
module FA_1007 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46709, net148762, net148733, net138080, n3, n4, n5;
  assign Co = net46709;

  NAND2_X1 U1 ( .A1(Ci), .A2(n5), .ZN(n4) );
  NAND2_X1 U2 ( .A1(n4), .A2(net138080), .ZN(net46709) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n5) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  CLKBUF_X1 U5 ( .A(A), .Z(net148733) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
  CLKBUF_X1 U7 ( .A(B), .Z(net148762) );
  NAND2_X1 U8 ( .A1(net148733), .A2(net148762), .ZN(net138080) );
endmodule


module FA_1006 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46706, n3, n4, n5, n6;
  assign Co = net46706;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46706) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_1005 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46703, n3, n4, n5, n6;
  assign Co = net46703;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46703) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_1004 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46700, n3, n4, n5, n6;
  assign Co = net46700;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46700) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_1003 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46697, n3, n4, n5, n6;
  assign Co = net46697;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46697) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_1002 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46694, n3, n4, n5, n6;
  assign Co = net46694;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46694) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_1001 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46691, n3, n4, n5, n6;
  assign Co = net46691;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46691) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_1000 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46688, n3, n4, n5, n6;
  assign Co = net46688;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46688) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_999 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46685, n3, n4, n5, n6;
  assign Co = net46685;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46685) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_998 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46682, n3, n4, n5, n6;
  assign Co = net46682;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46682) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_997 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46679, n3, n4, n5, n6;
  assign Co = net46679;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46679) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_996 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46676, n3, n4, n5, n6;
  assign Co = net46676;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46676) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_995 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46673, n3, n4, n5, n6;
  assign Co = net46673;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46673) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_994 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46670, n3, n4, n5, n6;
  assign Co = net46670;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46670) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_993 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46667, n3, n4, n5, n6;
  assign Co = net46667;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46667) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_992 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46664, n3, n4, n5, n6;
  assign Co = net46664;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46664) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_991 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46661, n3, n4, n5, n6;
  assign Co = net46661;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46661) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_990 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46658, n3, n4, n5, n6;
  assign Co = net46658;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46658) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_989 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46655, n3, n4, n5, n6;
  assign Co = net46655;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46655) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_988 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46652, n3, n4, n5, n6;
  assign Co = net46652;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46652) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_987 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46649, n3, n4, n5, n6;
  assign Co = net46649;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46649) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_986 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46646, n3, n4, n5, n6;
  assign Co = net46646;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46646) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_985 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46643, n3, n4, n5, n6;
  assign Co = net46643;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46643) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_984 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46640, net137989, net137988, n3, n4;
  assign Co = net46640;

  NAND2_X1 U1 ( .A1(Ci), .A2(n4), .ZN(net137989) );
  NAND2_X1 U2 ( .A1(net137989), .A2(net137988), .ZN(net46640) );
  INV_X1 U3 ( .A(n3), .ZN(n4) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(net137988) );
endmodule


module FA_983 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46637, n3, n4, n5, n6;
  assign Co = net46637;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46637) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_982 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46634, n3, n4, n5, n6;
  assign Co = net46634;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46634) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_981 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46631, n3, n4, n5, n6;
  assign Co = net46631;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46631) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_980 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46628, n3, n4, n5, n6;
  assign Co = net46628;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46628) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_979 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46625, n3, n4, n5, n6;
  assign Co = net46625;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46625) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_978 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46622, n3, n4, n5, n6;
  assign Co = net46622;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46622) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_977 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46619, n3, n4, n5, n6;
  assign Co = net46619;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46619) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_976 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46616, n3, n4, n5, n6;
  assign Co = net46616;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46616) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_975 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46613, n3, n4, n5, n6;
  assign Co = net46613;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46613) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_974 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46610, n3, n4, n5, n6;
  assign Co = net46610;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46610) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_973 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46607, n3, n4, n5, n6;
  assign Co = net46607;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46607) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_972 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46604, n3, n4, n5, n6;
  assign Co = net46604;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46604) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_971 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46601, n3, n4, n5, n6;
  assign Co = net46601;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46601) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_970 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46598, n3, n4, n5, n6;
  assign Co = net46598;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46598) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_969 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46595, n3, n4, n5, n6;
  assign Co = net46595;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46595) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_968 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46592, n3, n4, n5, n6;
  assign Co = net46592;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46592) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_967 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46589, n3, n4, n5, n6;
  assign Co = net46589;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46589) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_966 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46586, n3, n4, n5, n6;
  assign Co = net46586;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n4), .A2(n5), .ZN(net46586) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_965 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46583, net137913, net137912, n3, n4;
  assign Co = net46583;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(net137913) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n3) );
  INV_X1 U4 ( .A(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net137912) );
  NAND2_X1 U6 ( .A1(net137913), .A2(net137912), .ZN(net46583) );
endmodule


module FA_964 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46580, n3, n4, n5, n6;
  assign Co = net46580;

  NAND2_X1 U1 ( .A1(n4), .A2(n5), .ZN(net46580) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_963 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46577, n3, n4, n5, n6;
  assign Co = net46577;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net46577) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_962 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46574, n3, n4, n5, n6;
  assign Co = net46574;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net46574) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U4 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_961 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46571, n3, n4, n5, n6;
  assign Co = net46571;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net46571) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U4 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_960 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46568, n3, n4, n5, n6;
  assign Co = net46568;

  NAND2_X1 U1 ( .A1(n4), .A2(n5), .ZN(net46568) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_959 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46565, n3, n4, n5, n6;
  assign Co = net46565;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net46565) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U4 ( .A(n3), .ZN(n6) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_958 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46562, n3, n4, n5, n6;
  assign Co = net46562;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net46562) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_957 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46559, n3, n4, n5, n6;
  assign Co = net46559;

  NAND2_X1 U1 ( .A1(n4), .A2(n5), .ZN(net46559) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_956 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46556, n3, n4, n5, n6;
  assign Co = net46556;

  NAND2_X1 U1 ( .A1(n4), .A2(n5), .ZN(net46556) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_955 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46553, n3, n4, n5, n6;
  assign Co = net46553;

  NAND2_X1 U1 ( .A1(n4), .A2(n5), .ZN(net46553) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_954 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46550, n3, n4, n5, n6;
  assign Co = net46550;

  NAND2_X1 U1 ( .A1(n4), .A2(n5), .ZN(net46550) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_953 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46547, n3, n4, n5, n6;
  assign Co = net46547;

  NAND2_X1 U1 ( .A1(n4), .A2(n5), .ZN(net46547) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_952 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46544, n3, n4, n5, n6;
  assign Co = net46544;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net46544) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  INV_X1 U3 ( .A(n3), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_951 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net137856, net137857, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(net137857) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n3) );
  INV_X1 U4 ( .A(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net137856) );
  NAND2_X1 U6 ( .A1(net137856), .A2(net137857), .ZN(Co) );
endmodule


module FA_950 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_949 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_948 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_947 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_946 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_945 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_944 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  OAI21_X1 U1 ( .B1(n5), .B2(n6), .A(n4), .ZN(Co) );
  XNOR2_X1 U2 ( .A(n5), .B(Ci), .ZN(S) );
  CLKBUF_X1 U3 ( .A(B), .Z(n3) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n5) );
  INV_X1 U5 ( .A(Ci), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n3), .A2(A), .ZN(n4) );
endmodule


module FA_943 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_942 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_941 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_940 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n4), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_939 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_938 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_937 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_936 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_935 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_934 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_933 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_932 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_931 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_930 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_929 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_928 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_927 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_926 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_925 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_924 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_923 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_922 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_921 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_920 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46448, net137734, net137732, n3, n4, n5;
  assign Co = net46448;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(net137734) );
  XNOR2_X1 U3 ( .A(Ci), .B(n3), .ZN(S) );
  CLKBUF_X1 U4 ( .A(B), .Z(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(n4), .ZN(net137732) );
  NAND2_X1 U6 ( .A1(n5), .A2(net137732), .ZN(net46448) );
  NAND2_X1 U7 ( .A1(net137734), .A2(Ci), .ZN(n5) );
endmodule


module FA_919 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46445, n3, n4, n5, n6;
  assign Co = net46445;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net46445) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n3) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_918 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net137724, net137725, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(net137725) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(net137724) );
  XOR2_X1 U5 ( .A(A), .B(B), .Z(n4) );
  NAND2_X1 U6 ( .A1(net137725), .A2(net137724), .ZN(Co) );
endmodule


module FA_917 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_916 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_915 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_914 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_913 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_912 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  BUF_X1 U2 ( .A(n8), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n5) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_911 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_910 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_909 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_908 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_907 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_906 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_905 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_904 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_903 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_902 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_901 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net137656, net137657, net137658, n3, n4;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n4) );
  INV_X1 U3 ( .A(n4), .ZN(net137658) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(net137656) );
  XNOR2_X1 U5 ( .A(Ci), .B(n4), .ZN(S) );
  NAND2_X1 U6 ( .A1(Ci), .A2(net137658), .ZN(net137657) );
  NAND2_X1 U7 ( .A1(net137656), .A2(net137657), .ZN(Co) );
endmodule


module FA_900 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_899 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_898 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_897 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_896 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_895 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_894 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_893 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_892 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_891 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_890 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_889 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_888 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(Ci), .B(n6), .ZN(S) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U6 ( .A1(n5), .A2(n4), .ZN(Co) );
endmodule


module FA_887 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46349, net137600, n3, n4, n5;
  assign Co = net46349;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  NAND2_X1 U2 ( .A1(net137600), .A2(n5), .ZN(net46349) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(net137600) );
  XNOR2_X1 U5 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n4) );
endmodule


module FA_886 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net137596, net137597, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(net137597) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n3) );
  INV_X1 U4 ( .A(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net137596) );
  NAND2_X1 U6 ( .A1(net137596), .A2(net137597), .ZN(Co) );
endmodule


module FA_885 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_884 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_883 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_882 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_881 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_880 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XNOR2_X1 U1 ( .A(n4), .B(Ci), .ZN(S) );
  OAI21_X1 U2 ( .B1(n5), .B2(n4), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_879 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_878 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_877 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_876 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_875 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_874 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_873 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  XNOR2_X1 U3 ( .A(B), .B(n4), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_872 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_871 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_870 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_869 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_868 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_867 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_866 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_865 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_864 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(n3), .B(B), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_863 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_862 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_861 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_860 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_859 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_858 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_857 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_856 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_855 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_854 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46250, net137468, n3, n4, n5;
  assign Co = net46250;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U3 ( .A(Ci), .B(n4), .ZN(S) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(net137468) );
  NAND2_X1 U5 ( .A1(n5), .A2(net137468), .ZN(net46250) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n3), .ZN(n5) );
endmodule


module FA_853 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net137464, net137465, n3, n4, n5;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n5), .ZN(net137465) );
  NAND2_X1 U5 ( .A1(A), .A2(n3), .ZN(net137464) );
  XOR2_X1 U6 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U7 ( .A1(net137465), .A2(net137464), .ZN(Co) );
endmodule


module FA_852 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_851 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_850 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_849 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_848 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(n4), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_847 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_846 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_845 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_844 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_843 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_842 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_841 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_840 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_839 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_838 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_837 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46199, net137401, net137400, net137399, n3;
  assign Co = net46199;

  NAND2_X1 U1 ( .A1(Ci), .A2(n3), .ZN(net137401) );
  NAND2_X1 U2 ( .A1(net137401), .A2(net137400), .ZN(net46199) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U4 ( .A(Ci), .B(net137399), .ZN(S) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(net137399) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(net137400) );
endmodule


module FA_836 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46196, n3, n4, n5, n6;
  assign Co = net46196;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net46196) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_835 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46193, n3, n4, n5, n6;
  assign Co = net46193;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n4), .A2(n5), .ZN(net46193) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_834 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net137388, net137389, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(net137389) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net137388) );
  NAND2_X1 U6 ( .A1(net137389), .A2(net137388), .ZN(Co) );
endmodule


module FA_833 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_832 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_831 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_830 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(n3), .B(B), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_829 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_828 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_827 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_826 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_825 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_824 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_823 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_822 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46154, net137340, n3, n4, n5, n6;
  assign Co = net46154;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(net137340), .A2(n6), .ZN(net46154) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net137340) );
  XNOR2_X1 U6 ( .A(Ci), .B(n5), .ZN(S) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n5) );
endmodule


module FA_821 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net137336, net137337, n3, n4;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n3), .ZN(net137337) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net137336) );
  NAND2_X1 U6 ( .A1(net137336), .A2(net137337), .ZN(Co) );
endmodule


module FA_820 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_819 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_818 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_817 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_816 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XNOR2_X1 U1 ( .A(n4), .B(Ci), .ZN(S) );
  OAI21_X1 U2 ( .B1(n5), .B2(n4), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_815 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_814 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_813 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_812 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_811 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_810 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_809 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_808 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_807 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_806 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_805 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_804 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_803 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n3), .A2(A), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_802 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XOR2_X1 U3 ( .A(Ci), .B(n4), .Z(S) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
endmodule


module FA_801 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_800 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_799 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_798 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_797 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_796 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_795 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_794 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_793 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_792 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_791 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_790 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_789 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46055, net137210, net137208, n3, n4, n5;
  assign Co = net46055;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(net137210) );
  XNOR2_X1 U3 ( .A(n3), .B(Ci), .ZN(S) );
  CLKBUF_X1 U4 ( .A(B), .Z(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(n4), .ZN(net137208) );
  NAND2_X1 U6 ( .A1(n5), .A2(net137208), .ZN(net46055) );
  NAND2_X1 U7 ( .A1(Ci), .A2(net137210), .ZN(n5) );
endmodule


module FA_788 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46052, n3, n4, n5, n6;
  assign Co = net46052;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net46052) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_787 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net137200, net137201, n3, n4, n5;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n5), .ZN(net137201) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(net137200) );
  XOR2_X1 U6 ( .A(B), .B(A), .Z(n5) );
  NAND2_X1 U7 ( .A1(net137201), .A2(net137200), .ZN(Co) );
endmodule


module FA_786 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_785 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_784 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_783 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_782 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_781 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_780 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_779 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_778 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_777 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_776 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_775 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_774 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_773 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_772 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_771 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_770 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45998, net137133, net137132, net137131, n3;
  assign Co = net45998;

  NAND2_X1 U1 ( .A1(Ci), .A2(n3), .ZN(net137133) );
  NAND2_X1 U2 ( .A1(net137133), .A2(net137132), .ZN(net45998) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U4 ( .A(Ci), .B(net137131), .ZN(S) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(net137131) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(net137132) );
endmodule


module FA_769 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45995, n3, n4, n5, n6;
  assign Co = net45995;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n4), .A2(n5), .ZN(net45995) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_768 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45992, n3, n4, n5, n6;
  assign Co = net45992;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n4), .A2(n5), .ZN(net45992) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_767 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45989, n3, n4, n5, n6;
  assign Co = net45989;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net45989) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n4) );
endmodule


module FA_766 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45986, n3, n4, n5, n6, n7;
  assign Co = net45986;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n3), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(net45986) );
  XNOR2_X1 U4 ( .A(n4), .B(Ci), .ZN(S) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n4) );
  CLKBUF_X1 U6 ( .A(B), .Z(n7) );
  NAND2_X1 U7 ( .A1(A), .A2(n7), .ZN(n5) );
endmodule


module FA_765 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45983, n3, n4, n5, n6;
  assign Co = net45983;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n4), .A2(n5), .ZN(net45983) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_764 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45980, n3, n4, n5, n6;
  assign Co = net45980;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net45980) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_763 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45977, n3, n4, n5, n6;
  assign Co = net45977;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n4), .A2(n5), .ZN(net45977) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
endmodule


module FA_762 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45974, n3, n4, n5, n6, n7;
  assign Co = net45974;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n7), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(net45974) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n7) );
  XNOR2_X1 U5 ( .A(Ci), .B(n4), .ZN(S) );
  NAND2_X1 U6 ( .A1(A), .A2(n3), .ZN(n5) );
  XNOR2_X1 U7 ( .A(A), .B(B), .ZN(n4) );
endmodule


module FA_761 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45971, n3, n4, n5, n6;
  assign Co = net45971;

  NAND2_X1 U1 ( .A1(n6), .A2(Ci), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n4), .A2(n5), .ZN(net45971) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_760 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net137092, net137093, n3, n4;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n3), .ZN(net137093) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n4) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(net137092) );
  NAND2_X1 U6 ( .A1(net137093), .A2(net137092), .ZN(Co) );
endmodule


module FA_759 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_758 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_757 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45959, net137080, n3, n4, n5, n6;
  assign Co = net45959;

  XNOR2_X1 U1 ( .A(n3), .B(B), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(net137080), .A2(n6), .ZN(net45959) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net137080) );
  XNOR2_X1 U6 ( .A(Ci), .B(n5), .ZN(S) );
  XNOR2_X1 U7 ( .A(A), .B(B), .ZN(n5) );
endmodule


module FA_756 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net137076, net137077, n3, n4;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(n4), .B(Ci), .ZN(S) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n3), .ZN(net137077) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net137076) );
  NAND2_X1 U6 ( .A1(net137076), .A2(net137077), .ZN(Co) );
endmodule


module FA_755 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_754 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_753 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_752 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(n5), .B(Ci), .ZN(S) );
  OAI21_X1 U3 ( .B1(n6), .B2(n5), .A(n4), .ZN(Co) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n5) );
  INV_X1 U5 ( .A(Ci), .ZN(n6) );
  NAND2_X1 U6 ( .A1(A), .A2(n3), .ZN(n4) );
endmodule


module FA_751 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_750 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(n4), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n8), .B(Ci), .ZN(S) );
endmodule


module FA_749 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(n4), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_748 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_747 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_746 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_745 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_744 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_743 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_742 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_741 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_740 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_739 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_738 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  XNOR2_X1 U3 ( .A(B), .B(n4), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(n3), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n8), .B(Ci), .ZN(S) );
endmodule


module FA_737 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_736 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_735 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_734 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_733 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_732 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_731 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_730 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(n3), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_729 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_728 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_727 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_726 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n3), .A2(A), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_725 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_724 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_723 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45857, net136945, net136944, net148804, net136943, n3;
  assign Co = net45857;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(net136943), .ZN(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(net136943) );
  NAND2_X1 U4 ( .A1(Ci), .A2(net148804), .ZN(net136945) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net136944) );
  XNOR2_X1 U6 ( .A(B), .B(n3), .ZN(net148804) );
  NAND2_X1 U7 ( .A1(net136945), .A2(net136944), .ZN(net45857) );
endmodule


module FA_722 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45854, n3, n4, n5, n6, n7;
  assign Co = net45854;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(net45854) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U7 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_721 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45851, n3, n4, n5, n6, n7;
  assign Co = net45851;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n7) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(net45851) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U7 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_720 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45848, n3, n4, n5, n6, n7;
  assign Co = net45848;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  NAND2_X1 U2 ( .A1(n6), .A2(n5), .ZN(net45848) );
  NAND2_X1 U3 ( .A1(n3), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n7), .ZN(n6) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n7) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U7 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_719 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45845, n3, n4, n5, n6;
  assign Co = net45845;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net45845) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_718 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45842, n3, n4, n5, n6;
  assign Co = net45842;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net45842) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_717 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136920, net136921, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(net136921) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net136920) );
  NAND2_X1 U6 ( .A1(net136921), .A2(net136920), .ZN(Co) );
endmodule


module FA_716 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_715 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_714 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_713 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_712 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_711 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_710 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_709 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_708 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_707 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_706 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_705 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(n3), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_704 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_703 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_702 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_701 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_700 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_699 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_698 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_697 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_696 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45776, net136837, net136836, net136835, n3;
  assign Co = net45776;

  NAND2_X1 U1 ( .A1(Ci), .A2(n3), .ZN(net136837) );
  NAND2_X1 U2 ( .A1(net136836), .A2(net136837), .ZN(net45776) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U4 ( .A(Ci), .B(net136835), .ZN(S) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(net136835) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(net136836) );
endmodule


module FA_695 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45773, n3, n4, n5, n6, n7;
  assign Co = net45773;

  NAND2_X1 U1 ( .A1(Ci), .A2(n6), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n4), .A2(n5), .ZN(net45773) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n6) );
  XNOR2_X1 U4 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U5 ( .A1(A), .A2(n7), .ZN(n4) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
  CLKBUF_X1 U7 ( .A(B), .Z(n7) );
endmodule


module FA_694 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136828, net136829, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(net136829) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net136828) );
  NAND2_X1 U6 ( .A1(net136829), .A2(net136828), .ZN(Co) );
endmodule


module FA_693 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_692 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136820, net136821, net152734, n3;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(net136820) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(net152734) );
  NAND2_X1 U5 ( .A1(Ci), .A2(net152734), .ZN(net136821) );
  NAND2_X1 U6 ( .A1(net136821), .A2(net136820), .ZN(Co) );
endmodule


module FA_691 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_690 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_689 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_688 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XNOR2_X1 U1 ( .A(n4), .B(Ci), .ZN(S) );
  OAI21_X1 U2 ( .B1(n4), .B2(n5), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_687 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n4), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_686 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_685 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_684 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_683 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_682 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_681 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_680 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_679 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_678 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_677 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_676 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_675 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_674 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_673 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_672 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_671 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_670 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_669 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_668 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_667 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_666 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_665 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_664 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_663 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_662 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_661 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_660 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_659 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136687, net136688, net136689, n3;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n3), .ZN(net136689) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(net136687) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(net136688) );
  NAND2_X1 U5 ( .A1(net136689), .A2(net136688), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(net136687), .ZN(S) );
endmodule


module FA_658 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136684, net136685, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(net136685) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net136684) );
  NAND2_X1 U6 ( .A1(net136685), .A2(net136684), .ZN(Co) );
endmodule


module FA_657 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_656 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_655 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_654 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_653 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45647, net136664, n3, n4, n5;
  assign Co = net45647;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  NAND2_X1 U2 ( .A1(n5), .A2(net136664), .ZN(net45647) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(net136664) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n5) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U6 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_652 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136660, net136661, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n5) );
  XNOR2_X1 U2 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n4), .ZN(net136661) );
  XNOR2_X1 U5 ( .A(n5), .B(B), .ZN(n4) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(net136660) );
  NAND2_X1 U7 ( .A1(net136661), .A2(net136660), .ZN(Co) );
endmodule


module FA_651 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_650 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_649 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_648 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_647 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_646 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_645 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_644 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_643 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_642 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  BUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U4 ( .A1(n4), .A2(A), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(Ci), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n3), .B(Ci), .ZN(S) );
endmodule


module FA_641 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_640 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_639 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_638 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_637 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_636 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_635 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_634 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_633 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_632 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_631 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_630 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136572, net136573, net149086, n3, n4;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U3 ( .A1(A), .A2(n4), .ZN(net136572) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(net149086) );
  CLKBUF_X1 U5 ( .A(B), .Z(n4) );
  NAND2_X1 U6 ( .A1(Ci), .A2(net149086), .ZN(net136573) );
  NAND2_X1 U7 ( .A1(net136573), .A2(net136572), .ZN(Co) );
endmodule


module FA_629 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_628 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45572, net136564, n3, n4, n5, n6;
  assign Co = net45572;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  NAND2_X1 U2 ( .A1(net136564), .A2(n5), .ZN(net45572) );
  NAND2_X1 U3 ( .A1(n3), .A2(Ci), .ZN(n5) );
  NAND2_X1 U4 ( .A1(A), .A2(n6), .ZN(net136564) );
  CLKBUF_X1 U5 ( .A(B), .Z(n6) );
  XNOR2_X1 U6 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n4) );
endmodule


module FA_627 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136560, net136561, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n4), .A2(Ci), .ZN(net136561) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net136560) );
  NAND2_X1 U6 ( .A1(net136560), .A2(net136561), .ZN(Co) );
endmodule


module FA_626 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_625 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_624 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XNOR2_X1 U1 ( .A(n4), .B(Ci), .ZN(S) );
  OAI21_X1 U2 ( .B1(n4), .B2(n5), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_623 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_622 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_621 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  XNOR2_X1 U3 ( .A(B), .B(n4), .ZN(n5) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(n3), .ZN(n7) );
  NAND2_X1 U6 ( .A1(n5), .A2(Ci), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n8), .B(Ci), .ZN(S) );
endmodule


module FA_620 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_619 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_618 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_617 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_616 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_615 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_614 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_613 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_612 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_611 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_610 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_609 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_608 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_607 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_606 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_605 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_604 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_603 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_602 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_601 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_600 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_599 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(n3), .B(B), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_598 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_597 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n4), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_596 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_595 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_594 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136427, net136428, net136429, n3;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n3), .ZN(net136429) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(net136427) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(net136428) );
  NAND2_X1 U5 ( .A1(net136429), .A2(net136428), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(net136427), .ZN(S) );
endmodule


module FA_593 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136424, net136425, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(net136425) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net136424) );
  NAND2_X1 U6 ( .A1(net136425), .A2(net136424), .ZN(Co) );
endmodule


module FA_592 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_591 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_590 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_589 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n4), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_588 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136404, net136405, net148805, n3, n4;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(net148805), .ZN(net136405) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net136404) );
  XNOR2_X1 U6 ( .A(B), .B(n4), .ZN(net148805) );
  NAND2_X1 U7 ( .A1(net136404), .A2(net136405), .ZN(Co) );
endmodule


module FA_587 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_586 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_585 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_584 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_583 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_582 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_581 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_580 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_579 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_578 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  INV_X1 U2 ( .A(A), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(n4), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_577 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_576 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_575 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  XNOR2_X1 U3 ( .A(B), .B(n4), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_574 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_573 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_572 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_571 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_570 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_569 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  CLKBUF_X1 U3 ( .A(B), .Z(n5) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(n5), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n4), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_568 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_567 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_566 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45386, net136317, net136316, net136315, n3, n4;
  assign Co = net45386;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n4), .ZN(net136317) );
  NAND2_X1 U3 ( .A1(net136316), .A2(net136317), .ZN(net45386) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(net136315), .ZN(S) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(net136315) );
  NAND2_X1 U7 ( .A1(A), .A2(n3), .ZN(net136316) );
endmodule


module FA_565 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136312, net136313, n3, n4, n5;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n5), .ZN(net136313) );
  XOR2_X1 U5 ( .A(A), .B(B), .Z(n5) );
  NAND2_X1 U6 ( .A1(A), .A2(n3), .ZN(net136312) );
  NAND2_X1 U7 ( .A1(net136312), .A2(net136313), .ZN(Co) );
endmodule


module FA_564 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_563 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136304, net136305, net149729, n3;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(Ci), .ZN(S) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(net136304) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(net149729) );
  NAND2_X1 U5 ( .A1(Ci), .A2(net149729), .ZN(net136305) );
  NAND2_X1 U6 ( .A1(net136304), .A2(net136305), .ZN(Co) );
endmodule


module FA_562 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_561 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_560 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XNOR2_X1 U1 ( .A(n4), .B(Ci), .ZN(S) );
  OAI21_X1 U2 ( .B1(n4), .B2(n5), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_559 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_558 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_557 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_556 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_555 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n3), .A2(A), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_554 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_553 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_552 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_551 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_550 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_549 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_548 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_547 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_546 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n4), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_545 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  XNOR2_X1 U3 ( .A(n4), .B(B), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_544 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_543 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_542 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_541 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_540 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_539 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_538 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_537 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_536 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_535 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_534 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_533 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_532 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_531 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_530 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_529 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136167, net136168, net136169, n3;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n3), .ZN(net136169) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(net136167) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(net136168) );
  NAND2_X1 U5 ( .A1(net136169), .A2(net136168), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(net136167), .ZN(S) );
endmodule


module FA_528 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136164, net136165, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(net136165) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n4) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(net136164) );
  NAND2_X1 U6 ( .A1(net136165), .A2(net136164), .ZN(Co) );
endmodule


module FA_527 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_526 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_525 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_524 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45260, net136149, net136148, net136147, n3;
  assign Co = net45260;

  NAND2_X1 U1 ( .A1(net136149), .A2(net136148), .ZN(net45260) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n3), .ZN(net136149) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n3) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(net136148) );
  XNOR2_X1 U5 ( .A(Ci), .B(net136147), .ZN(S) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(net136147) );
endmodule


module FA_523 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45257, n3, n4, n5, n6;
  assign Co = net45257;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net45257) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_522 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45254, n3, n4, n5, n6;
  assign Co = net45254;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net45254) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_521 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45251, n3, n4, n5, n6;
  assign Co = net45251;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net45251) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n6) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_520 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45248, n3, n4, n5, n6, n7;
  assign Co = net45248;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net45248) );
  NAND2_X1 U2 ( .A1(A), .A2(n6), .ZN(n4) );
  CLKBUF_X1 U3 ( .A(B), .Z(n6) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n7), .ZN(n5) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n7) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_519 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45245, n3, n4, n5, n6, n7;
  assign Co = net45245;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net45245) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U4 ( .A(n7), .B(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_518 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45242, n3, n4, n5, n6, n7;
  assign Co = net45242;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(net45242) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U7 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_517 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45239, n3, n4, n5, n6;
  assign Co = net45239;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net45239) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U5 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_516 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45236, n3, n4, n5, n6, n7;
  assign Co = net45236;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net45236) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n7), .ZN(n5) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n6), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(B), .Z(n6) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_515 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45233, n3, n4, n5, n6, n7;
  assign Co = net45233;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(net45233) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U5 ( .A1(n7), .A2(Ci), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U7 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_514 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45230, n3, n4, n5, n6, n7;
  assign Co = net45230;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net45230) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U5 ( .A(B), .B(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_513 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45227, n3, n4, n5, n6, n7;
  assign Co = net45227;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(net45227) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U7 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_512 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45224, n3, n4, n5, n6, n7;
  assign Co = net45224;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net45224) );
  NAND2_X1 U2 ( .A1(A), .A2(n6), .ZN(n4) );
  CLKBUF_X1 U3 ( .A(B), .Z(n6) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n7), .ZN(n5) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n7) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_511 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45221, n3, n4, n5, n6, n7;
  assign Co = net45221;

  NAND2_X1 U1 ( .A1(n4), .A2(n5), .ZN(net45221) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n7), .ZN(n5) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n6), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(B), .Z(n6) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_510 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45218, n3, n4, n5, n6, n7;
  assign Co = net45218;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n4), .A2(n5), .ZN(net45218) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(n7), .ZN(n6) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n4) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_509 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136088, net136089, n3, n4, n5;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n5), .ZN(net136089) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n5) );
  NAND2_X1 U6 ( .A1(A), .A2(n3), .ZN(net136088) );
  NAND2_X1 U7 ( .A1(net136088), .A2(net136089), .ZN(Co) );
endmodule


module FA_508 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_507 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_506 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_505 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_504 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_503 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_502 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_501 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45191, net136057, net136056, net136055, n3, n4;
  assign Co = net45191;

  NAND2_X1 U1 ( .A1(Ci), .A2(n3), .ZN(net136057) );
  NAND2_X1 U2 ( .A1(net136056), .A2(net136057), .ZN(net45191) );
  XOR2_X1 U3 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U4 ( .A(Ci), .B(net136055), .ZN(S) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(net136055) );
  NAND2_X1 U6 ( .A1(A), .A2(n4), .ZN(net136056) );
  CLKBUF_X1 U7 ( .A(B), .Z(n4) );
endmodule


module FA_500 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136052, net136053, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(net136053) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(net136052) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n4) );
  NAND2_X1 U6 ( .A1(net136052), .A2(net136053), .ZN(Co) );
endmodule


module FA_499 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net136048, net136049, net149575, n3, n4;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U3 ( .A(Ci), .B(n4), .ZN(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(net149575) );
  NAND2_X1 U5 ( .A1(A), .A2(n3), .ZN(net136048) );
  NAND2_X1 U6 ( .A1(Ci), .A2(net149575), .ZN(net136049) );
  NAND2_X1 U7 ( .A1(net136048), .A2(net136049), .ZN(Co) );
endmodule


module FA_498 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_497 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(n7), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_496 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U1 ( .A(n4), .B(n5), .Z(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n4) );
  OAI21_X1 U3 ( .B1(n4), .B2(n5), .A(n3), .ZN(Co) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_495 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_494 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_493 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_492 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_491 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_490 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_489 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_488 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(n3), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_487 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_486 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_485 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_484 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_483 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_482 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_481 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_480 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_479 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_478 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_477 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_476 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_475 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_474 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_473 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_472 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_471 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_470 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_469 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_468 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_467 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_466 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_465 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_464 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135907, net135908, net135909, n3;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n3), .ZN(net135909) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(net135907) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(net135908) );
  NAND2_X1 U5 ( .A1(net135909), .A2(net135908), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(net135907), .ZN(S) );
endmodule


module FA_463 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135904, net135905, n3, n4;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(net135905) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n4) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net135904) );
  NAND2_X1 U6 ( .A1(net135904), .A2(net135905), .ZN(Co) );
endmodule


module FA_462 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_461 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_460 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(n3), .B(B), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_459 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_458 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_457 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_456 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_455 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_454 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_453 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_452 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_451 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_450 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_449 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_448 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_447 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_446 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_445 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45023, net135833, net135832, net135831, n3;
  assign Co = net45023;

  NAND2_X1 U1 ( .A1(net135833), .A2(net135832), .ZN(net45023) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(net135832) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n3), .ZN(net135833) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(net135831) );
  XNOR2_X1 U6 ( .A(Ci), .B(net135831), .ZN(S) );
endmodule


module FA_444 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45020, n3, n4, n5, n6, n7;
  assign Co = net45020;

  NAND2_X1 U1 ( .A1(n4), .A2(n5), .ZN(net45020) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(n7), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(B), .Z(n7) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_443 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45017, n3, n4, n5, n6, n7;
  assign Co = net45017;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  NAND2_X1 U2 ( .A1(n6), .A2(n5), .ZN(net45017) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n7), .ZN(n6) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n7) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(n5) );
  XNOR2_X1 U6 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n4) );
endmodule


module FA_442 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45014, n3, n4, n5, n6, n7, n8;
  assign Co = net45014;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n8) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(net45014) );
  NAND2_X1 U4 ( .A1(A), .A2(n7), .ZN(n5) );
  CLKBUF_X1 U5 ( .A(B), .Z(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n8), .ZN(n6) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U8 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_441 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45011, n3, n4, n5, n6, n7, n8;
  assign Co = net45011;

  INV_X1 U1 ( .A(A), .ZN(n8) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  NAND2_X1 U3 ( .A1(n5), .A2(n6), .ZN(net45011) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n7), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n8), .ZN(n7) );
  NAND2_X1 U6 ( .A1(n3), .A2(A), .ZN(n5) );
  XNOR2_X1 U7 ( .A(n4), .B(Ci), .ZN(S) );
  XNOR2_X1 U8 ( .A(B), .B(A), .ZN(n4) );
endmodule


module FA_440 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45008, n3, n4, n5, n6, n7, n8;
  assign Co = net45008;

  INV_X1 U1 ( .A(A), .ZN(n8) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  NAND2_X1 U3 ( .A1(n6), .A2(n5), .ZN(net45008) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n7), .ZN(n6) );
  XNOR2_X1 U5 ( .A(B), .B(n8), .ZN(n7) );
  NAND2_X1 U6 ( .A1(n3), .A2(A), .ZN(n5) );
  XNOR2_X1 U7 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U8 ( .A(B), .B(A), .ZN(n4) );
endmodule


module FA_439 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net45005, n3, n4, n5, n6, n7;
  assign Co = net45005;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  NAND2_X1 U2 ( .A1(n6), .A2(n5), .ZN(net45005) );
  NAND2_X1 U3 ( .A1(n3), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n7), .ZN(n6) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(n7) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U7 ( .A(Ci), .B(n4), .ZN(S) );
endmodule


module FA_438 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135804, net135805, n3, n4, n5;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n5), .ZN(net135805) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(net135804) );
  XOR2_X1 U6 ( .A(B), .B(A), .Z(n5) );
  NAND2_X1 U7 ( .A1(net135805), .A2(net135804), .ZN(Co) );
endmodule


module FA_437 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_436 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135796, net135797, net148884, n3;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n3), .ZN(S) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(net148884) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(net135796) );
  NAND2_X1 U5 ( .A1(net148884), .A2(Ci), .ZN(net135797) );
  NAND2_X1 U6 ( .A1(net135797), .A2(net135796), .ZN(Co) );
endmodule


module FA_435 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135792, net135793, net149073, n3, n4, n5;

  XNOR2_X1 U1 ( .A(n3), .B(B), .ZN(net149073) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n5) );
  XNOR2_X1 U5 ( .A(n5), .B(Ci), .ZN(S) );
  NAND2_X1 U6 ( .A1(A), .A2(n4), .ZN(net135792) );
  NAND2_X1 U7 ( .A1(Ci), .A2(net149073), .ZN(net135793) );
  NAND2_X1 U8 ( .A1(net135792), .A2(net135793), .ZN(Co) );
endmodule


module FA_434 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_433 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_432 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U1 ( .A(n4), .B(n5), .Z(S) );
  OAI21_X1 U2 ( .B1(n4), .B2(n5), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_431 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_430 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_429 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_428 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_427 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_426 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_425 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_424 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_423 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n3), .A2(A), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_422 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n3), .A2(A), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_421 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_420 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(n3), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_419 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_418 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_417 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_416 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_415 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_414 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_413 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_412 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_411 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_410 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_409 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_408 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_407 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_406 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_405 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_404 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_403 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_402 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_401 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_400 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_399 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135647, net135648, net135649, n3;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n3), .ZN(net135649) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(net135647) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(net135648) );
  NAND2_X1 U5 ( .A1(net135649), .A2(net135648), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(net135647), .ZN(S) );
endmodule


module FA_398 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44882, n3, n4, n5, n6, n7;
  assign Co = net44882;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net44882) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U5 ( .A(B), .B(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_397 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44879, n3, n4, n5, n6, n7;
  assign Co = net44879;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net44879) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U5 ( .A(n7), .B(B), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_396 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44876, n3, n4, n5, n6, n7;
  assign Co = net44876;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net44876) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U5 ( .A(B), .B(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_395 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135632, net135633, n3, n4, n5;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n5) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n5), .ZN(net135633) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(net135632) );
  NAND2_X1 U7 ( .A1(net135633), .A2(net135632), .ZN(Co) );
endmodule


module FA_394 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_393 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_392 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_391 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_390 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_389 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_388 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_387 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_386 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_385 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_384 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_383 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_382 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_381 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_380 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_379 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_378 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_377 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_376 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n4), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_375 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_374 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135548, net135549, net148779, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n5) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U4 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U5 ( .A(B), .B(n5), .ZN(net148779) );
  NAND2_X1 U6 ( .A1(A), .A2(n3), .ZN(net135548) );
  NAND2_X1 U7 ( .A1(Ci), .A2(net148779), .ZN(net135549) );
  NAND2_X1 U8 ( .A1(net135549), .A2(net135548), .ZN(Co) );
endmodule


module FA_373 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  XNOR2_X1 U3 ( .A(B), .B(n4), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_372 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44804, net135541, net135540, net135539, n3, n4;
  assign Co = net44804;

  NAND2_X1 U1 ( .A1(n3), .A2(Ci), .ZN(net135541) );
  NAND2_X1 U2 ( .A1(net135541), .A2(net135540), .ZN(net44804) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U4 ( .A(Ci), .B(net135539), .ZN(S) );
  CLKBUF_X1 U5 ( .A(B), .Z(n4) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(net135539) );
  NAND2_X1 U7 ( .A1(n4), .A2(A), .ZN(net135540) );
endmodule


module FA_371 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135536, net135537, net149082, n3;

  XNOR2_X1 U1 ( .A(n3), .B(Ci), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(net149082), .ZN(net135537) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(net135536) );
  XOR2_X1 U5 ( .A(B), .B(A), .Z(net149082) );
  NAND2_X1 U6 ( .A1(net135537), .A2(net135536), .ZN(Co) );
endmodule


module FA_370 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_369 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(n7), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_368 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U1 ( .A(n4), .B(n5), .Z(S) );
  OAI21_X1 U2 ( .B1(n4), .B2(n5), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_367 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_366 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_365 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_364 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_363 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_362 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_361 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_360 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_359 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_358 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_357 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n3), .A2(A), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_356 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_355 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_354 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_353 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_352 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_351 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_350 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n3), .A2(A), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_349 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_348 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_347 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_346 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_345 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_344 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_343 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n3), .A2(A), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_342 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_341 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_340 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_339 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_338 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_337 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_336 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_335 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_334 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_333 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_332 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_331 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135376, net135377, net148753, n3;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n3), .ZN(S) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(net135376) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(net148753) );
  NAND2_X1 U5 ( .A1(Ci), .A2(net148753), .ZN(net135377) );
  NAND2_X1 U6 ( .A1(net135377), .A2(net135376), .ZN(Co) );
endmodule


module FA_330 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(n3), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_329 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_328 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_327 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_326 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_325 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_324 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_323 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_322 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_321 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_320 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_319 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_318 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_317 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_316 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_315 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_314 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  XNOR2_X1 U3 ( .A(B), .B(n4), .ZN(n5) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_313 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_312 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_311 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_310 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44618, net135293, net135292, net135291, n3;
  assign Co = net44618;

  NAND2_X1 U1 ( .A1(net135293), .A2(net135292), .ZN(net44618) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(net135292) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n3), .ZN(net135293) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(net135291) );
  XNOR2_X1 U6 ( .A(Ci), .B(net135291), .ZN(S) );
endmodule


module FA_309 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44615, n3, n4, n5, n6, n7;
  assign Co = net44615;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net44615) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n6) );
  NAND2_X1 U4 ( .A1(A), .A2(n7), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(B), .Z(n7) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n3) );
endmodule


module FA_308 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44612, n3, n4, n5, n6;
  assign Co = net44612;

  NAND2_X1 U1 ( .A1(n5), .A2(n4), .ZN(net44612) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n6) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U6 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_307 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44609, net135281, net135280, net135279, n3, n4;
  assign Co = net44609;

  NAND2_X1 U1 ( .A1(Ci), .A2(n3), .ZN(net135281) );
  NAND2_X1 U2 ( .A1(net135281), .A2(net135280), .ZN(net44609) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U4 ( .A(Ci), .B(net135279), .ZN(S) );
  XNOR2_X1 U5 ( .A(B), .B(A), .ZN(net135279) );
  CLKBUF_X1 U6 ( .A(B), .Z(n4) );
  NAND2_X1 U7 ( .A1(A), .A2(n4), .ZN(net135280) );
endmodule


module FA_306 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135276, net135277, n3, n4, n5;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n4), .ZN(net135277) );
  CLKBUF_X1 U5 ( .A(B), .Z(n5) );
  NAND2_X1 U6 ( .A1(A), .A2(n5), .ZN(net135276) );
  NAND2_X1 U7 ( .A1(net135276), .A2(net135277), .ZN(Co) );
endmodule


module FA_305 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n7) );
  INV_X1 U5 ( .A(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_304 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U1 ( .A(n4), .B(n5), .Z(S) );
  OAI21_X1 U2 ( .B1(n4), .B2(n5), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_303 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_302 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_301 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_300 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_299 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_298 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_297 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_296 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_295 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_294 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_293 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_292 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_291 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_290 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_289 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_288 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_287 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_286 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_285 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_284 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_283 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_282 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_281 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_280 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_279 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_278 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(n4), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_277 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_276 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_275 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_274 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_273 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(n3), .B(B), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_272 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_271 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_270 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_269 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_268 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_267 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135120, net135121, net147396, n3, n4;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U4 ( .A(B), .B(n4), .ZN(net147396) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(net135120) );
  NAND2_X1 U6 ( .A1(Ci), .A2(net147396), .ZN(net135121) );
  NAND2_X1 U7 ( .A1(net135121), .A2(net135120), .ZN(Co) );
endmodule


module FA_266 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_265 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(n4), .A2(Ci), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_264 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_263 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n4), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_262 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_261 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_260 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_259 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_258 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_257 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_256 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_255 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_254 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_253 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_252 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_251 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_250 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_249 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_248 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_247 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_246 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(n4), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_245 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_244 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_243 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135024, net135025, net148778, n3, n4, n5;

  INV_X1 U1 ( .A(A), .ZN(n5) );
  CLKBUF_X1 U2 ( .A(B), .Z(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U4 ( .A(Ci), .B(n4), .ZN(S) );
  XNOR2_X1 U5 ( .A(B), .B(n5), .ZN(net148778) );
  NAND2_X1 U6 ( .A1(n3), .A2(A), .ZN(net135024) );
  NAND2_X1 U7 ( .A1(Ci), .A2(net148778), .ZN(net135025) );
  NAND2_X1 U8 ( .A1(net135024), .A2(net135025), .ZN(Co) );
endmodule


module FA_242 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net135020, net135021, net148887, n3, n4;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n3), .ZN(S) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(net148887) );
  NAND2_X1 U5 ( .A1(n4), .A2(A), .ZN(net135020) );
  NAND2_X1 U6 ( .A1(Ci), .A2(net148887), .ZN(net135021) );
  NAND2_X1 U7 ( .A1(net135020), .A2(net135021), .ZN(Co) );
endmodule


module FA_241 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8, n9;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  CLKBUF_X1 U2 ( .A(n9), .Z(n4) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n5) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n9) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(n8) );
  INV_X1 U6 ( .A(n4), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n5), .A2(n6), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n8), .A2(n7), .ZN(Co) );
  XNOR2_X1 U9 ( .A(n9), .B(Ci), .ZN(S) );
endmodule


module FA_240 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U1 ( .A(n4), .B(n5), .Z(S) );
  OAI21_X1 U2 ( .B1(n4), .B2(n5), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_239 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_238 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_237 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_236 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_235 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_234 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_233 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_232 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_231 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(n6), .B(Ci), .ZN(S) );
endmodule


module FA_230 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_229 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_228 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_227 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_226 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_225 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_224 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  BUF_X1 U1 ( .A(n7), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_223 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_222 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_221 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_220 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_219 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(n7), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_218 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_217 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_216 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_215 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_214 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_213 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_212 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_211 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_210 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(B), .ZN(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_209 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_208 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_207 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_206 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_205 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_204 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_203 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net134863, net134864, net134865, n3;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n3), .ZN(net134865) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(net134864) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(net134863) );
  NAND2_X1 U5 ( .A1(net134865), .A2(net134864), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(net134863), .ZN(S) );
endmodule


module FA_202 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_201 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_200 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_199 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(n3), .B(B), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_198 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_197 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44279, n3, n4, n5, n6, n7;
  assign Co = net44279;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net44279) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U5 ( .A(B), .B(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_196 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44276, n3, n4, n5, n6, n7;
  assign Co = net44276;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net44276) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U5 ( .A(B), .B(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_195 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_194 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_193 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44267, n3, n4, n5, n6, n7;
  assign Co = net44267;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net44267) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U5 ( .A(B), .B(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_192 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_191 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_190 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44258, n3, n4, n5, n6, n7;
  assign Co = net44258;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net44258) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U5 ( .A(n7), .B(B), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_189 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_188 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44252, n3, n4, n5, n6, n7;
  assign Co = net44252;

  INV_X1 U1 ( .A(A), .ZN(n7) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net44252) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n4) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U5 ( .A(B), .B(n7), .ZN(n6) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_187 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_186 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_185 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_184 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_183 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_182 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44234, n3, n4, n5, n6, n7, n8;
  assign Co = net44234;

  INV_X1 U1 ( .A(A), .ZN(n8) );
  NAND2_X1 U2 ( .A1(n5), .A2(n4), .ZN(net44234) );
  NAND2_X1 U3 ( .A1(n7), .A2(A), .ZN(n4) );
  CLKBUF_X1 U4 ( .A(B), .Z(n7) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n6), .ZN(n5) );
  XNOR2_X1 U6 ( .A(B), .B(n8), .ZN(n6) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U8 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_181 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net134776, net134777, n3, n4, n5;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  NAND2_X1 U3 ( .A1(Ci), .A2(n4), .ZN(net134777) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(n4) );
  CLKBUF_X1 U5 ( .A(B), .Z(n5) );
  NAND2_X1 U6 ( .A1(A), .A2(n5), .ZN(net134776) );
  NAND2_X1 U7 ( .A1(net134777), .A2(net134776), .ZN(Co) );
endmodule


module FA_180 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  CLKBUF_X1 U2 ( .A(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n4), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_179 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net134768, net134769, net148793, n3, n4;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(Ci), .B(n3), .ZN(S) );
  XNOR2_X1 U4 ( .A(B), .B(n4), .ZN(net148793) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(net134768) );
  NAND2_X1 U6 ( .A1(Ci), .A2(net148793), .ZN(net134769) );
  NAND2_X1 U7 ( .A1(net134769), .A2(net134768), .ZN(Co) );
endmodule


module FA_178 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net134764, net134765, net148581, n3, n4;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(Ci), .B(n3), .ZN(S) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(net148581) );
  NAND2_X1 U5 ( .A1(n4), .A2(A), .ZN(net134764) );
  NAND2_X1 U6 ( .A1(Ci), .A2(net148581), .ZN(net134765) );
  NAND2_X1 U7 ( .A1(net134765), .A2(net134764), .ZN(Co) );
endmodule


module FA_177 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n7) );
  INV_X1 U5 ( .A(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_176 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U1 ( .A(n4), .B(n5), .Z(S) );
  OAI21_X1 U2 ( .B1(n4), .B2(n5), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_175 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_174 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_173 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_172 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_171 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_170 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_169 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_168 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_167 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_166 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_165 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_164 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_163 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_162 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_161 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_160 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_159 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_158 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_157 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_156 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_155 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_154 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_153 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_152 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  BUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_151 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_150 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_149 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_148 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_147 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_146 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n3), .ZN(n4) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n5) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n5), .B(n4), .ZN(S) );
endmodule


module FA_145 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_144 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_143 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n5) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n3), .B(n4), .ZN(S) );
endmodule


module FA_142 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_141 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_140 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_139 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XOR2_X1 U2 ( .A(A), .B(B), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_138 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(n7), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(Ci), .ZN(S) );
endmodule


module FA_137 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(n7), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(Ci), .ZN(S) );
endmodule


module FA_136 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_135 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  BUF_X1 U1 ( .A(n7), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n3), .ZN(S) );
endmodule


module FA_134 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_133 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  BUF_X1 U1 ( .A(Ci), .Z(n3) );
  INV_X1 U2 ( .A(A), .ZN(n4) );
  XNOR2_X1 U3 ( .A(n4), .B(B), .ZN(n5) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n3), .B(n8), .ZN(S) );
endmodule


module FA_132 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_131 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_130 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_129 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_128 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_127 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_126 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_125 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n6) );
  NAND2_X1 U3 ( .A1(B), .A2(A), .ZN(n5) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_124 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n6) );
  XNOR2_X1 U3 ( .A(n4), .B(B), .ZN(n3) );
  INV_X1 U4 ( .A(n3), .ZN(n5) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n8) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n3), .ZN(n7) );
  NAND2_X1 U7 ( .A1(n7), .A2(n8), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n6), .B(n5), .ZN(S) );
endmodule


module FA_123 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_122 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  BUF_X1 U1 ( .A(B), .Z(n3) );
  CLKBUF_X1 U2 ( .A(n3), .Z(n4) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n5) );
  XNOR2_X1 U4 ( .A(n3), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n4), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_121 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(n7) );
  XNOR2_X1 U3 ( .A(B), .B(n4), .ZN(n3) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n7), .B(Ci), .ZN(S) );
endmodule


module FA_120 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(n3), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_119 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XNOR2_X1 U1 ( .A(B), .B(n3), .ZN(n4) );
  INV_X32 U2 ( .A(A), .ZN(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_118 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_117 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net134520, net134521, net147405, n3, n4;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n4) );
  XNOR2_X1 U3 ( .A(Ci), .B(n4), .ZN(S) );
  XOR2_X1 U4 ( .A(B), .B(A), .Z(net147405) );
  NAND2_X1 U5 ( .A1(n3), .A2(A), .ZN(net134520) );
  NAND2_X1 U6 ( .A1(Ci), .A2(net147405), .ZN(net134521) );
  NAND2_X1 U7 ( .A1(net134521), .A2(net134520), .ZN(Co) );
endmodule


module FA_116 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(B), .Z(n3) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U4 ( .A1(n3), .A2(A), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_115 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44033, net134513, net134512, net134511, n3, n4, n5;
  assign Co = net44033;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  NAND2_X1 U3 ( .A1(net134513), .A2(net134512), .ZN(net44033) );
  NAND2_X1 U4 ( .A1(n4), .A2(A), .ZN(net134512) );
  CLKBUF_X1 U5 ( .A(B), .Z(n4) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(net134513) );
  XNOR2_X1 U7 ( .A(B), .B(A), .ZN(net134511) );
  XNOR2_X1 U8 ( .A(Ci), .B(net134511), .ZN(S) );
endmodule


module FA_114 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net44030, net134509, net134508, net134507, n3, n4;
  assign Co = net44030;

  NAND2_X1 U1 ( .A1(n3), .A2(Ci), .ZN(net134509) );
  NAND2_X1 U2 ( .A1(net134509), .A2(net134508), .ZN(net44030) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U4 ( .A(Ci), .B(net134507), .ZN(S) );
  CLKBUF_X1 U5 ( .A(B), .Z(n4) );
  XNOR2_X1 U6 ( .A(B), .B(A), .ZN(net134507) );
  NAND2_X1 U7 ( .A1(A), .A2(n4), .ZN(net134508) );
endmodule


module FA_113 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net134504, net134506, net149730, net149817, n3, n4, n5;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(net149817) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n3) );
  CLKBUF_X1 U4 ( .A(n3), .Z(net149730) );
  CLKBUF_X1 U5 ( .A(B), .Z(n4) );
  NAND2_X1 U6 ( .A1(n4), .A2(A), .ZN(net134504) );
  INV_X1 U7 ( .A(net149730), .ZN(net134506) );
  NAND2_X1 U8 ( .A1(net149817), .A2(net134506), .ZN(n5) );
  NAND2_X1 U9 ( .A1(net134504), .A2(n5), .ZN(Co) );
endmodule


module FA_112 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5;

  XOR2_X1 U1 ( .A(n4), .B(n5), .Z(S) );
  OAI21_X1 U2 ( .B1(n4), .B2(n5), .A(n3), .ZN(Co) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n4) );
  INV_X1 U4 ( .A(Ci), .ZN(n5) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n3) );
endmodule


module FA_111 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_110 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_109 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_108 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_107 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_106 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_105 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_104 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_103 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_102 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_101 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_100 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_99 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(n3), .A2(Ci), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_98 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_97 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_96 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  INV_X1 U1 ( .A(A), .ZN(n4) );
  INV_X1 U2 ( .A(n3), .ZN(n7) );
  XNOR2_X1 U3 ( .A(n4), .B(B), .ZN(n3) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(Ci), .B(n7), .ZN(S) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(n7), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U5 ( .A(n7), .ZN(n4) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U7 ( .A1(n6), .A2(n5), .ZN(Co) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n5) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n4), .B(n3), .ZN(S) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n5) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n4), .B(n3), .ZN(S) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(n7), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U5 ( .A(n7), .ZN(n4) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U7 ( .A1(n6), .A2(n5), .ZN(Co) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n6), .A2(n5), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(n7), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U5 ( .A(n7), .ZN(n4) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U7 ( .A1(n6), .A2(n5), .ZN(Co) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n5) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n4), .B(n3), .ZN(S) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(n3), .B(n7), .ZN(S) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U5 ( .A(n7), .ZN(n4) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U7 ( .A1(n6), .A2(n5), .ZN(Co) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(n4), .B(n3), .ZN(S) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U6 ( .A(n8), .ZN(n5) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U8 ( .A1(n6), .A2(n7), .ZN(Co) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(Ci), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n4), .B(n3), .ZN(S) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(Ci), .B(n6), .ZN(S) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U4 ( .A(n6), .ZN(n3) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U6 ( .A1(n4), .A2(n5), .ZN(Co) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n4), .A2(n5), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(n4), .B(n3), .ZN(S) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U6 ( .A(n8), .ZN(n5) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U8 ( .A1(n6), .A2(n7), .ZN(Co) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  CLKBUF_X1 U1 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n7) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n6) );
  INV_X1 U4 ( .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n4), .ZN(n5) );
  NAND2_X1 U6 ( .A1(n5), .A2(n6), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n3), .B(n7), .ZN(S) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(n4), .B(n3), .ZN(S) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U6 ( .A(n8), .ZN(n5) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U8 ( .A1(n6), .A2(n7), .ZN(Co) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(n4), .B(n3), .ZN(S) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U6 ( .A(n8), .ZN(n5) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U8 ( .A1(n6), .A2(n7), .ZN(Co) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  BUF_X1 U1 ( .A(Ci), .Z(n4) );
  CLKBUF_X1 U2 ( .A(n8), .Z(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n5) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n7), .A2(n6), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n4), .B(n3), .ZN(S) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n6) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n5) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n3), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n5), .A2(n4), .ZN(Co) );
  XNOR2_X1 U6 ( .A(Ci), .B(n6), .ZN(S) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n5) );
  XOR2_X1 U2 ( .A(n6), .B(n3), .Z(S) );
  CLKBUF_X1 U3 ( .A(n4), .Z(n3) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(Ci), .Z(n6) );
  NAND2_X1 U6 ( .A1(B), .A2(A), .ZN(n8) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n7), .A2(n8), .ZN(Co) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n5) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n4), .B(n3), .ZN(S) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(n4), .B(n3), .ZN(S) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(B), .A2(A), .ZN(n7) );
  INV_X1 U6 ( .A(n8), .ZN(n5) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U8 ( .A1(n6), .A2(n7), .ZN(Co) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n4), .B(n8), .ZN(S) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n7) );
  INV_X1 U5 ( .A(n8), .ZN(n5) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n4), .B(n3), .ZN(S) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7;

  XOR2_X1 U1 ( .A(A), .B(B), .Z(n3) );
  INV_X1 U2 ( .A(n3), .ZN(n4) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n5) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n7) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n5), .B(n4), .ZN(S) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  CLKBUF_X1 U1 ( .A(n8), .Z(n3) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(n4) );
  XNOR2_X1 U3 ( .A(n4), .B(n3), .ZN(S) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(A), .A2(B), .ZN(n7) );
  INV_X1 U6 ( .A(n8), .ZN(n5) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U8 ( .A1(n6), .A2(n7), .ZN(Co) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net134264, n3, n4, n5, n6;

  BUF_X1 U1 ( .A(Ci), .Z(n5) );
  XOR2_X1 U2 ( .A(B), .B(A), .Z(n3) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n4) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(net134264) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n3), .ZN(n6) );
  NAND2_X1 U6 ( .A1(n6), .A2(net134264), .ZN(Co) );
  XNOR2_X1 U7 ( .A(n5), .B(n4), .ZN(S) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8, n9;

  INV_X1 U1 ( .A(A), .ZN(n5) );
  INV_X1 U2 ( .A(n4), .ZN(n9) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n3) );
  XNOR2_X1 U4 ( .A(B), .B(n5), .ZN(n4) );
  CLKBUF_X1 U5 ( .A(B), .Z(n6) );
  NAND2_X1 U6 ( .A1(A), .A2(n6), .ZN(n8) );
  NAND2_X1 U7 ( .A1(Ci), .A2(n4), .ZN(n7) );
  NAND2_X1 U8 ( .A1(n7), .A2(n8), .ZN(Co) );
  XNOR2_X1 U9 ( .A(n3), .B(n9), .ZN(S) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  BUF_X1 U1 ( .A(Ci), .Z(n3) );
  BUF_X1 U2 ( .A(B), .Z(n4) );
  XOR2_X1 U3 ( .A(B), .B(A), .Z(n5) );
  XNOR2_X1 U4 ( .A(n4), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n4), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(n3), .B(n8), .ZN(S) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n4, n5, n6, n7, n8;

  INV_X1 U1 ( .A(A), .ZN(n3) );
  XNOR2_X1 U2 ( .A(B), .B(n3), .ZN(n5) );
  CLKBUF_X1 U3 ( .A(B), .Z(n4) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n8) );
  NAND2_X1 U5 ( .A1(n4), .A2(A), .ZN(n7) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n5), .ZN(n6) );
  NAND2_X1 U7 ( .A1(n6), .A2(n7), .ZN(Co) );
  XNOR2_X1 U8 ( .A(Ci), .B(n8), .ZN(S) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net134248, net134250, net148436, net148468, n3, n4, n5;

  XNOR2_X1 U1 ( .A(Ci), .B(n3), .ZN(S) );
  CLKBUF_X1 U2 ( .A(Ci), .Z(net148436) );
  XNOR2_X1 U3 ( .A(B), .B(A), .ZN(n3) );
  CLKBUF_X1 U4 ( .A(n3), .Z(net148468) );
  CLKBUF_X1 U5 ( .A(B), .Z(n4) );
  NAND2_X1 U6 ( .A1(n4), .A2(A), .ZN(net134248) );
  INV_X1 U7 ( .A(net148468), .ZN(net134250) );
  NAND2_X1 U8 ( .A1(net148436), .A2(net134250), .ZN(n5) );
  NAND2_X1 U9 ( .A1(net134248), .A2(n5), .ZN(Co) );
endmodule


module RCA_generic_N64_14 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_944 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_943 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_942 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_941 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_940 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_939 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_938 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_937 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_936 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_935 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_934 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_933 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_932 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_931 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_930 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_929 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_928 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_927 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_926 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_925 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_924 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_923 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_922 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_921 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_920 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_919 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_918 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_917 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_916 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_915 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_914 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_913 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_912 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_911 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_910 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_909 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_908 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_907 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_906 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_905 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_904 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_903 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_902 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_901 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_900 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_899 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_898 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_897 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_896 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_895 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_894 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_893 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_892 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_891 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_890 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_889 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_888 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_887 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_886 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_885 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_884 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_883 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_882 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_881 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_13 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_880 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_879 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_878 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_877 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_876 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_875 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_874 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_873 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_872 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_871 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_870 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_869 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_868 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_867 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_866 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_865 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_864 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_863 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_862 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_861 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_860 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_859 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_858 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_857 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_856 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_855 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_854 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_853 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_852 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_851 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_850 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_849 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_848 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_847 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_846 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_845 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_844 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_843 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_842 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_841 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_840 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_839 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_838 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_837 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_836 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_835 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_834 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_833 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_832 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_831 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_830 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_829 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_828 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_827 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_826 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_825 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_824 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_823 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_822 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_821 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_820 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_819 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_818 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_817 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_12 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_816 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_815 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_814 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_813 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_812 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_811 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_810 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_809 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_808 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_807 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_806 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_805 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_804 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_803 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_802 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_801 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_800 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_799 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_798 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_797 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_796 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_795 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_794 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_793 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_792 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_791 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_790 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_789 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_788 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_787 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_786 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_785 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_784 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_783 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_782 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_781 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_780 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_779 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_778 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_777 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_776 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_775 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_774 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_773 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_772 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_771 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_770 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_769 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_768 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_767 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_766 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_765 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_764 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_763 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_762 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_761 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_760 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_759 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_758 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_757 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_756 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_755 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_754 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_753 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_11 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_752 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_751 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_750 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_749 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_748 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_747 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_746 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_745 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_744 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_743 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_742 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_741 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_740 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_739 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_738 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_737 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_736 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_735 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_734 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_733 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_732 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_731 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_730 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_729 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_728 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_727 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_726 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_725 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_724 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_723 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_722 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_721 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_720 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_719 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_718 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_717 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_716 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_715 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_714 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_713 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_712 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_711 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_710 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_709 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_708 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_707 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_706 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_705 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_704 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_703 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_702 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_701 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_700 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_699 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_698 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_697 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_696 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_695 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_694 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_693 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_692 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_691 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_690 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_689 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_10 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_688 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_687 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_686 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_685 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_684 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_683 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_682 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_681 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_680 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_679 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_678 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_677 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_676 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_675 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_674 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_673 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_672 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_671 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_670 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_669 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_668 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_667 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_666 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_665 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_664 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_663 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_662 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_661 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_660 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_659 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_658 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_657 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_656 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_655 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_654 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_653 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_652 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_651 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_650 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_649 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_648 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_647 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_646 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_645 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_644 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_643 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_642 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_641 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_640 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_639 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_638 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_637 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_636 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_635 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_634 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_633 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_632 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_631 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_630 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_629 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_628 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_627 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_626 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_625 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_9 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_624 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_623 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_622 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_621 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_620 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_619 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_618 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_617 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_616 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_615 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_614 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_613 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_612 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_611 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_610 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_609 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_608 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_607 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_606 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_605 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_604 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_603 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_602 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_601 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_600 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_599 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_598 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_597 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_596 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_595 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_594 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_593 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_592 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_591 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_590 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_589 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_588 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_587 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_586 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_585 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_584 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_583 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_582 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_581 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_580 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_579 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_578 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_577 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_576 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_575 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_574 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_573 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_572 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_571 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_570 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_569 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_568 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_567 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_566 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_565 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_564 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_563 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_562 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_561 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_8 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_560 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_559 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_558 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_557 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_556 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_555 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_554 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_553 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_552 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_551 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_550 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_549 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_548 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_547 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_546 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_545 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_544 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_543 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_542 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_541 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_540 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_539 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_538 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_537 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_536 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_535 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_534 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_533 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_532 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_531 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_530 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_529 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_528 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_527 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_526 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_525 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_524 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_523 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_522 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_521 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_520 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_519 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_518 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_517 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_516 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_515 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_514 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_513 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_512 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_511 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_510 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_509 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_508 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_507 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_506 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_505 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_504 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_503 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_502 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_501 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_500 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_499 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_498 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_497 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_7 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_496 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_495 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_494 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_493 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_492 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_491 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_490 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_489 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_488 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_487 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_486 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_485 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_484 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_483 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_482 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_481 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_480 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_479 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_478 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_477 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_476 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_475 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_474 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_473 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_472 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_471 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_470 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_469 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_468 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_467 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_466 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_465 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_464 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_463 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_462 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_461 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_460 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_459 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_458 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_457 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_456 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_455 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_454 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_453 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_452 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_451 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_450 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_449 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_448 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_447 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_446 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_445 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_444 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_443 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_442 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_441 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_440 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_439 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_438 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_437 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_436 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_435 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_434 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_433 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_6 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_432 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_431 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_430 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_429 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_428 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_427 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_426 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_425 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_424 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_423 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_422 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_421 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_420 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_419 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_418 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_417 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_416 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_415 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_414 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_413 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_412 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_411 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_410 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_409 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_408 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_407 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_406 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_405 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_404 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_403 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_402 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_401 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_400 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_399 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_398 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_397 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_396 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_395 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_394 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_393 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_392 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_391 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_390 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_389 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_388 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_387 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_386 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_385 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_384 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_383 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_382 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_381 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_380 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_379 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_378 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_377 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_376 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_375 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_374 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_373 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_372 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_371 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_370 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_369 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_5 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_368 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_367 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_366 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_365 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_364 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_363 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_362 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_361 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_360 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_359 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_358 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_357 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_356 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_355 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_354 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_353 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_352 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_351 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_350 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_349 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_348 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_347 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_346 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_345 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_344 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_343 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_342 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_341 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_340 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_339 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_338 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_337 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_336 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_335 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_334 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_333 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_332 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_331 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_330 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_329 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_328 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_327 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_326 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_325 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_324 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_323 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_322 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_321 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_320 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_319 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_318 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_317 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_316 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_315 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_314 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_313 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_312 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_311 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_310 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_309 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_308 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_307 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_306 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_305 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_4 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_304 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_303 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_302 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_301 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_300 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_299 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_298 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_297 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_296 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_295 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_294 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_293 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_292 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_291 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_290 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_289 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_288 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_287 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_286 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_285 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_284 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_283 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_282 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_281 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_280 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_279 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_278 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_277 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_276 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_275 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_274 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_273 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_272 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_271 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_270 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_269 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_268 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_267 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_266 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_265 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_264 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_263 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_262 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_261 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_260 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_259 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_258 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_257 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_256 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_255 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_254 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_253 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_252 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_251 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_250 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_249 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_248 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_247 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_246 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_245 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_244 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_243 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_242 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_241 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_3 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_240 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_239 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_238 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_237 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_236 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_235 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_234 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_233 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_232 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_231 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_230 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_229 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_228 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_227 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_226 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_225 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_224 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_223 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_222 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_221 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_220 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_219 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_218 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_217 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_216 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_215 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_214 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_213 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_212 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_211 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_210 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_209 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_208 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_207 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_206 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_205 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_204 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_203 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_202 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_201 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_200 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_199 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_198 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_197 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_196 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_195 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_194 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_193 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_192 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_191 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_190 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_189 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_188 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_187 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_186 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_185 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_184 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_183 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_182 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_181 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_180 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_179 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_178 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_177 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_2 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_176 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_175 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_174 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_173 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_172 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_171 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_170 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_169 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_168 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_167 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_166 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_165 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_164 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_163 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_162 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_161 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_160 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_159 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_158 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_157 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_156 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_155 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_154 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_153 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_152 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_151 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_150 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_149 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_148 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_147 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_146 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_145 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_144 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_143 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_142 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_141 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_140 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_139 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_138 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_137 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_136 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_135 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_134 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_133 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_132 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_131 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_130 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_129 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_128 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_127 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_126 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_125 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_124 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_123 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_122 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_121 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_120 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_119 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_118 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_117 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_116 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_115 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_114 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_113 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module RCA_generic_N64_1 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_112 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_111 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_110 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_109 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_108 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_107 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_106 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_105 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_104 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_103 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_102 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_101 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_100 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_99 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14])
         );
  FA_98 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15])
         );
  FA_97 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16])
         );
  FA_96 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17])
         );
  FA_95 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18])
         );
  FA_94 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19])
         );
  FA_93 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20])
         );
  FA_92 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21])
         );
  FA_91 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22])
         );
  FA_90 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23])
         );
  FA_89 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24])
         );
  FA_88 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25])
         );
  FA_87 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26])
         );
  FA_86 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27])
         );
  FA_85 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28])
         );
  FA_84 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29])
         );
  FA_83 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30])
         );
  FA_82 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31])
         );
  FA_81 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32])
         );
  FA_80 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33])
         );
  FA_79 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34])
         );
  FA_78 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35])
         );
  FA_77 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36])
         );
  FA_76 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37])
         );
  FA_75 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38])
         );
  FA_74 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39])
         );
  FA_73 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40])
         );
  FA_72 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41])
         );
  FA_71 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42])
         );
  FA_70 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43])
         );
  FA_69 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44])
         );
  FA_68 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45])
         );
  FA_67 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46])
         );
  FA_66 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47])
         );
  FA_65 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48])
         );
  FA_64 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49])
         );
  FA_63 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50])
         );
  FA_62 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51])
         );
  FA_61 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52])
         );
  FA_60 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53])
         );
  FA_59 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54])
         );
  FA_58 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55])
         );
  FA_57 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56])
         );
  FA_56 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57])
         );
  FA_55 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58])
         );
  FA_54 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59])
         );
  FA_53 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60])
         );
  FA_52 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61])
         );
  FA_51 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62])
         );
  FA_50 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63])
         );
  FA_49 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module MUX51_GENERIC_N64_15 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   net141885, net141886, net141888, net142145, net146767, net146765,
         net146761, net146759, net146781, net146779, net146777, net146775,
         net146793, net146791, net146789, net146787, net146785, net146805,
         net146803, net146801, net146799, net146797, net146817, net146815,
         net146813, net146811, net146809, net148625, net142137, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408;

  AND2_X2 U1 ( .A1(n153), .A2(n149), .ZN(n139) );
  INV_X1 U2 ( .A(E[1]), .ZN(n140) );
  BUF_X1 U3 ( .A(net141885), .Z(net146781) );
  OR2_X1 U4 ( .A1(net142145), .A2(n140), .ZN(n160) );
  BUF_X4 U5 ( .A(n145), .Z(net146767) );
  NOR2_X1 U6 ( .A1(n151), .A2(SEL[2]), .ZN(n153) );
  AND2_X1 U7 ( .A1(SEL[1]), .A2(n152), .ZN(n141) );
  BUF_X2 U8 ( .A(net141886), .Z(net146787) );
  NOR2_X1 U9 ( .A1(n143), .A2(n144), .ZN(n142) );
  AND2_X1 U10 ( .A1(net141886), .A2(D[1]), .ZN(n143) );
  AND2_X1 U11 ( .A1(B[1]), .A2(n139), .ZN(n144) );
  CLKBUF_X1 U12 ( .A(n139), .Z(net146797) );
  AND2_X1 U13 ( .A1(n152), .A2(SEL[1]), .ZN(n145) );
  AND2_X1 U14 ( .A1(n148), .A2(n149), .ZN(n146) );
  AND2_X2 U15 ( .A1(n154), .A2(SEL[1]), .ZN(net141886) );
  INV_X1 U16 ( .A(n151), .ZN(n147) );
  NOR2_X1 U17 ( .A1(n147), .A2(SEL[1]), .ZN(n150) );
  INV_X1 U18 ( .A(SEL[1]), .ZN(n149) );
  INV_X1 U19 ( .A(SEL[0]), .ZN(n151) );
  NOR2_X1 U20 ( .A1(n151), .A2(SEL[2]), .ZN(n154) );
  NOR2_X1 U21 ( .A1(n155), .A2(SEL[2]), .ZN(n148) );
  NOR2_X1 U22 ( .A1(SEL[2]), .A2(n155), .ZN(n152) );
  NAND2_X1 U23 ( .A1(SEL[2]), .A2(E[0]), .ZN(net142137) );
  OAI21_X1 U24 ( .B1(SEL[2]), .B2(n150), .A(net148625), .ZN(net142145) );
  BUF_X1 U25 ( .A(SEL[0]), .Z(n155) );
  NAND2_X1 U26 ( .A1(n148), .A2(n149), .ZN(net148625) );
  NAND4_X1 U27 ( .A1(n158), .A2(net142137), .A3(n156), .A4(n157), .ZN(Y[0]) );
  NAND2_X1 U28 ( .A1(D[0]), .A2(net141886), .ZN(n157) );
  NAND2_X1 U29 ( .A1(B[0]), .A2(n139), .ZN(n156) );
  AOI22_X1 U30 ( .A1(C[0]), .A2(n141), .B1(n146), .B2(A[0]), .ZN(n158) );
  NAND3_X1 U31 ( .A1(n160), .A2(n159), .A3(n142), .ZN(Y[1]) );
  BUF_X4 U32 ( .A(net141888), .Z(net146809) );
  CLKBUF_X1 U33 ( .A(net141888), .Z(net146815) );
  BUF_X4 U34 ( .A(net141885), .Z(net146779) );
  CLKBUF_X1 U35 ( .A(net141886), .Z(net146791) );
  CLKBUF_X1 U36 ( .A(net141886), .Z(net146789) );
  CLKBUF_X1 U37 ( .A(net141886), .Z(net146785) );
  CLKBUF_X1 U38 ( .A(net141888), .Z(net146811) );
  CLKBUF_X1 U39 ( .A(net141888), .Z(net146813) );
  CLKBUF_X1 U40 ( .A(n139), .Z(net146803) );
  CLKBUF_X1 U41 ( .A(n139), .Z(net146801) );
  CLKBUF_X1 U42 ( .A(n139), .Z(net146799) );
  CLKBUF_X1 U43 ( .A(n145), .Z(net146759) );
  CLKBUF_X1 U44 ( .A(n145), .Z(net146761) );
  CLKBUF_X1 U45 ( .A(n145), .Z(net146765) );
  CLKBUF_X1 U46 ( .A(net141885), .Z(net146775) );
  CLKBUF_X1 U47 ( .A(net141885), .Z(net146777) );
  CLKBUF_X1 U48 ( .A(net141888), .Z(net146817) );
  CLKBUF_X1 U49 ( .A(n139), .Z(net146805) );
  CLKBUF_X1 U50 ( .A(net141886), .Z(net146793) );
  INV_X1 U51 ( .A(net142145), .ZN(net141888) );
  INV_X1 U52 ( .A(net148625), .ZN(net141885) );
  AOI22_X1 U53 ( .A1(C[1]), .A2(n145), .B1(A[1]), .B2(net141885), .ZN(n159) );
  NAND2_X1 U54 ( .A1(E[2]), .A2(net141888), .ZN(n164) );
  NAND2_X1 U55 ( .A1(B[2]), .A2(net146805), .ZN(n163) );
  NAND2_X1 U56 ( .A1(D[2]), .A2(net146787), .ZN(n162) );
  AOI22_X1 U57 ( .A1(C[2]), .A2(net146759), .B1(A[2]), .B2(net146775), .ZN(
        n161) );
  NAND4_X1 U58 ( .A1(n164), .A2(n163), .A3(n162), .A4(n161), .ZN(Y[2]) );
  NAND2_X1 U59 ( .A1(E[3]), .A2(net146815), .ZN(n168) );
  NAND2_X1 U60 ( .A1(B[3]), .A2(net146797), .ZN(n167) );
  NAND2_X1 U61 ( .A1(D[3]), .A2(net146785), .ZN(n166) );
  AOI22_X1 U62 ( .A1(C[3]), .A2(net146759), .B1(A[3]), .B2(net146781), .ZN(
        n165) );
  NAND4_X1 U63 ( .A1(n168), .A2(n167), .A3(n166), .A4(n165), .ZN(Y[3]) );
  NAND2_X1 U64 ( .A1(E[4]), .A2(net146811), .ZN(n172) );
  NAND2_X1 U65 ( .A1(B[4]), .A2(net146799), .ZN(n171) );
  NAND2_X1 U66 ( .A1(D[4]), .A2(net146793), .ZN(n170) );
  AOI22_X1 U67 ( .A1(C[4]), .A2(net146761), .B1(A[4]), .B2(net146781), .ZN(
        n169) );
  NAND4_X1 U68 ( .A1(n172), .A2(n171), .A3(n170), .A4(n169), .ZN(Y[4]) );
  NAND2_X1 U69 ( .A1(E[5]), .A2(net146813), .ZN(n176) );
  NAND2_X1 U70 ( .A1(B[5]), .A2(net146801), .ZN(n175) );
  NAND2_X1 U71 ( .A1(D[5]), .A2(net146791), .ZN(n174) );
  AOI22_X1 U72 ( .A1(C[5]), .A2(net146761), .B1(A[5]), .B2(net146781), .ZN(
        n173) );
  NAND4_X1 U73 ( .A1(n176), .A2(n175), .A3(n174), .A4(n173), .ZN(Y[5]) );
  NAND2_X1 U74 ( .A1(E[6]), .A2(net146817), .ZN(n180) );
  NAND2_X1 U75 ( .A1(B[6]), .A2(net146803), .ZN(n179) );
  NAND2_X1 U76 ( .A1(D[6]), .A2(net146789), .ZN(n178) );
  AOI22_X1 U77 ( .A1(C[6]), .A2(net146765), .B1(A[6]), .B2(net146777), .ZN(
        n177) );
  NAND4_X1 U78 ( .A1(n180), .A2(n179), .A3(n178), .A4(n177), .ZN(Y[6]) );
  NAND2_X1 U79 ( .A1(E[7]), .A2(net146809), .ZN(n184) );
  NAND2_X1 U80 ( .A1(B[7]), .A2(net146803), .ZN(n183) );
  NAND2_X1 U81 ( .A1(D[7]), .A2(net146787), .ZN(n182) );
  AOI22_X1 U82 ( .A1(C[7]), .A2(net146767), .B1(A[7]), .B2(net146779), .ZN(
        n181) );
  NAND4_X1 U83 ( .A1(n184), .A2(n183), .A3(n182), .A4(n181), .ZN(Y[7]) );
  NAND2_X1 U84 ( .A1(E[8]), .A2(net146809), .ZN(n188) );
  NAND2_X1 U85 ( .A1(B[8]), .A2(net146803), .ZN(n187) );
  NAND2_X1 U86 ( .A1(D[8]), .A2(net146785), .ZN(n186) );
  AOI22_X1 U87 ( .A1(C[8]), .A2(net146767), .B1(A[8]), .B2(net146779), .ZN(
        n185) );
  NAND4_X1 U88 ( .A1(n188), .A2(n187), .A3(n186), .A4(n185), .ZN(Y[8]) );
  NAND2_X1 U89 ( .A1(E[9]), .A2(net146809), .ZN(n192) );
  NAND2_X1 U90 ( .A1(B[9]), .A2(net146803), .ZN(n191) );
  NAND2_X1 U91 ( .A1(D[9]), .A2(net146793), .ZN(n190) );
  AOI22_X1 U92 ( .A1(C[9]), .A2(net146767), .B1(A[9]), .B2(net146779), .ZN(
        n189) );
  NAND4_X1 U93 ( .A1(n192), .A2(n191), .A3(n190), .A4(n189), .ZN(Y[9]) );
  NAND2_X1 U94 ( .A1(E[10]), .A2(net146809), .ZN(n196) );
  NAND2_X1 U95 ( .A1(B[10]), .A2(net146803), .ZN(n195) );
  NAND2_X1 U96 ( .A1(D[10]), .A2(net146791), .ZN(n194) );
  AOI22_X1 U97 ( .A1(C[10]), .A2(net146767), .B1(A[10]), .B2(net146779), .ZN(
        n193) );
  NAND4_X1 U98 ( .A1(n196), .A2(n195), .A3(n194), .A4(n193), .ZN(Y[10]) );
  NAND2_X1 U99 ( .A1(E[11]), .A2(net146809), .ZN(n200) );
  NAND2_X1 U100 ( .A1(B[11]), .A2(net146803), .ZN(n199) );
  NAND2_X1 U101 ( .A1(D[11]), .A2(net146789), .ZN(n198) );
  AOI22_X1 U102 ( .A1(C[11]), .A2(net146767), .B1(A[11]), .B2(net146779), .ZN(
        n197) );
  NAND4_X1 U103 ( .A1(n200), .A2(n199), .A3(n198), .A4(n197), .ZN(Y[11]) );
  NAND2_X1 U104 ( .A1(E[12]), .A2(net146809), .ZN(n204) );
  NAND2_X1 U105 ( .A1(B[12]), .A2(net146797), .ZN(n203) );
  NAND2_X1 U106 ( .A1(D[12]), .A2(net146787), .ZN(n202) );
  AOI22_X1 U107 ( .A1(C[12]), .A2(net146767), .B1(A[12]), .B2(net146779), .ZN(
        n201) );
  NAND4_X1 U108 ( .A1(n204), .A2(n203), .A3(n202), .A4(n201), .ZN(Y[12]) );
  NAND2_X1 U109 ( .A1(E[13]), .A2(net146809), .ZN(n208) );
  NAND2_X1 U110 ( .A1(B[13]), .A2(net146797), .ZN(n207) );
  NAND2_X1 U111 ( .A1(D[13]), .A2(net146785), .ZN(n206) );
  AOI22_X1 U112 ( .A1(C[13]), .A2(net146767), .B1(A[13]), .B2(net146779), .ZN(
        n205) );
  NAND4_X1 U113 ( .A1(n208), .A2(n207), .A3(n206), .A4(n205), .ZN(Y[13]) );
  NAND2_X1 U114 ( .A1(E[14]), .A2(net146809), .ZN(n212) );
  NAND2_X1 U115 ( .A1(B[14]), .A2(net146797), .ZN(n211) );
  NAND2_X1 U116 ( .A1(D[14]), .A2(net146793), .ZN(n210) );
  AOI22_X1 U117 ( .A1(C[14]), .A2(net146767), .B1(A[14]), .B2(net146779), .ZN(
        n209) );
  NAND4_X1 U118 ( .A1(n212), .A2(n211), .A3(n210), .A4(n209), .ZN(Y[14]) );
  NAND2_X1 U119 ( .A1(E[15]), .A2(net146809), .ZN(n216) );
  NAND2_X1 U120 ( .A1(B[15]), .A2(net146797), .ZN(n215) );
  NAND2_X1 U121 ( .A1(D[15]), .A2(net146791), .ZN(n214) );
  AOI22_X1 U122 ( .A1(C[15]), .A2(net146767), .B1(A[15]), .B2(net146779), .ZN(
        n213) );
  NAND4_X1 U123 ( .A1(n216), .A2(n215), .A3(n214), .A4(n213), .ZN(Y[15]) );
  NAND2_X1 U124 ( .A1(E[16]), .A2(net146809), .ZN(n220) );
  NAND2_X1 U125 ( .A1(B[16]), .A2(net146797), .ZN(n219) );
  NAND2_X1 U126 ( .A1(D[16]), .A2(net146789), .ZN(n218) );
  AOI22_X1 U127 ( .A1(C[16]), .A2(net146767), .B1(A[16]), .B2(net146779), .ZN(
        n217) );
  NAND4_X1 U128 ( .A1(n220), .A2(n219), .A3(n218), .A4(n217), .ZN(Y[16]) );
  NAND2_X1 U129 ( .A1(E[17]), .A2(net146809), .ZN(n224) );
  NAND2_X1 U130 ( .A1(B[17]), .A2(net146797), .ZN(n223) );
  NAND2_X1 U131 ( .A1(D[17]), .A2(net146787), .ZN(n222) );
  AOI22_X1 U132 ( .A1(C[17]), .A2(net146767), .B1(A[17]), .B2(net146779), .ZN(
        n221) );
  NAND4_X1 U133 ( .A1(n224), .A2(n223), .A3(n222), .A4(n221), .ZN(Y[17]) );
  NAND2_X1 U134 ( .A1(E[18]), .A2(net146817), .ZN(n228) );
  NAND2_X1 U135 ( .A1(B[18]), .A2(net146797), .ZN(n227) );
  NAND2_X1 U136 ( .A1(D[18]), .A2(net146785), .ZN(n226) );
  AOI22_X1 U137 ( .A1(C[18]), .A2(net146767), .B1(A[18]), .B2(net146779), .ZN(
        n225) );
  NAND4_X1 U138 ( .A1(n228), .A2(n227), .A3(n226), .A4(n225), .ZN(Y[18]) );
  NAND2_X1 U139 ( .A1(E[19]), .A2(net146809), .ZN(n232) );
  NAND2_X1 U140 ( .A1(B[19]), .A2(net146797), .ZN(n231) );
  NAND2_X1 U141 ( .A1(D[19]), .A2(net146793), .ZN(n230) );
  AOI22_X1 U142 ( .A1(C[19]), .A2(net146767), .B1(A[19]), .B2(net146779), .ZN(
        n229) );
  NAND4_X1 U143 ( .A1(n232), .A2(n231), .A3(n230), .A4(n229), .ZN(Y[19]) );
  NAND2_X1 U144 ( .A1(E[20]), .A2(net146817), .ZN(n236) );
  NAND2_X1 U145 ( .A1(B[20]), .A2(net146797), .ZN(n235) );
  NAND2_X1 U146 ( .A1(D[20]), .A2(net146791), .ZN(n234) );
  AOI22_X1 U147 ( .A1(C[20]), .A2(net146767), .B1(A[20]), .B2(net146779), .ZN(
        n233) );
  NAND4_X1 U148 ( .A1(n236), .A2(n235), .A3(n234), .A4(n233), .ZN(Y[20]) );
  NAND2_X1 U149 ( .A1(E[21]), .A2(net146809), .ZN(n240) );
  NAND2_X1 U150 ( .A1(B[21]), .A2(net146797), .ZN(n239) );
  NAND2_X1 U151 ( .A1(D[21]), .A2(net146789), .ZN(n238) );
  AOI22_X1 U152 ( .A1(C[21]), .A2(net146767), .B1(A[21]), .B2(net146779), .ZN(
        n237) );
  NAND4_X1 U153 ( .A1(n240), .A2(n239), .A3(n238), .A4(n237), .ZN(Y[21]) );
  NAND2_X1 U154 ( .A1(E[22]), .A2(net146817), .ZN(n244) );
  NAND2_X1 U155 ( .A1(B[22]), .A2(net146797), .ZN(n243) );
  NAND2_X1 U156 ( .A1(D[22]), .A2(net146787), .ZN(n242) );
  AOI22_X1 U157 ( .A1(C[22]), .A2(net146767), .B1(A[22]), .B2(net146779), .ZN(
        n241) );
  NAND4_X1 U158 ( .A1(n244), .A2(n243), .A3(n242), .A4(n241), .ZN(Y[22]) );
  NAND2_X1 U159 ( .A1(E[23]), .A2(net146809), .ZN(n248) );
  NAND2_X1 U160 ( .A1(B[23]), .A2(net146797), .ZN(n247) );
  NAND2_X1 U161 ( .A1(D[23]), .A2(net146785), .ZN(n246) );
  AOI22_X1 U162 ( .A1(C[23]), .A2(net146767), .B1(A[23]), .B2(net146779), .ZN(
        n245) );
  NAND4_X1 U163 ( .A1(n248), .A2(n247), .A3(n246), .A4(n245), .ZN(Y[23]) );
  NAND2_X1 U164 ( .A1(E[24]), .A2(net146817), .ZN(n252) );
  NAND2_X1 U165 ( .A1(B[24]), .A2(net146799), .ZN(n251) );
  NAND2_X1 U166 ( .A1(D[24]), .A2(net146793), .ZN(n250) );
  AOI22_X1 U167 ( .A1(C[24]), .A2(net146767), .B1(A[24]), .B2(net146779), .ZN(
        n249) );
  NAND4_X1 U168 ( .A1(n252), .A2(n251), .A3(n250), .A4(n249), .ZN(Y[24]) );
  NAND2_X1 U169 ( .A1(E[25]), .A2(net146809), .ZN(n256) );
  NAND2_X1 U170 ( .A1(B[25]), .A2(net146799), .ZN(n255) );
  NAND2_X1 U171 ( .A1(D[25]), .A2(net146791), .ZN(n254) );
  AOI22_X1 U172 ( .A1(C[25]), .A2(net146767), .B1(A[25]), .B2(net146779), .ZN(
        n253) );
  NAND4_X1 U173 ( .A1(n256), .A2(n255), .A3(n254), .A4(n253), .ZN(Y[25]) );
  NAND2_X1 U174 ( .A1(E[26]), .A2(net146817), .ZN(n260) );
  NAND2_X1 U175 ( .A1(B[26]), .A2(net146799), .ZN(n259) );
  NAND2_X1 U176 ( .A1(D[26]), .A2(net146789), .ZN(n258) );
  AOI22_X1 U177 ( .A1(C[26]), .A2(net146767), .B1(A[26]), .B2(net146779), .ZN(
        n257) );
  NAND4_X1 U178 ( .A1(n260), .A2(n259), .A3(n258), .A4(n257), .ZN(Y[26]) );
  NAND2_X1 U179 ( .A1(E[27]), .A2(net146809), .ZN(n264) );
  NAND2_X1 U180 ( .A1(B[27]), .A2(net146799), .ZN(n263) );
  NAND2_X1 U181 ( .A1(D[27]), .A2(net146787), .ZN(n262) );
  AOI22_X1 U182 ( .A1(C[27]), .A2(net146767), .B1(A[27]), .B2(net146779), .ZN(
        n261) );
  NAND4_X1 U183 ( .A1(n264), .A2(n263), .A3(n262), .A4(n261), .ZN(Y[27]) );
  NAND2_X1 U184 ( .A1(E[28]), .A2(net146817), .ZN(n268) );
  NAND2_X1 U185 ( .A1(B[28]), .A2(net146799), .ZN(n267) );
  NAND2_X1 U186 ( .A1(D[28]), .A2(net146785), .ZN(n266) );
  AOI22_X1 U187 ( .A1(C[28]), .A2(net146767), .B1(A[28]), .B2(net146779), .ZN(
        n265) );
  NAND4_X1 U188 ( .A1(n268), .A2(n267), .A3(n266), .A4(n265), .ZN(Y[28]) );
  NAND2_X1 U189 ( .A1(E[29]), .A2(net146809), .ZN(n272) );
  NAND2_X1 U190 ( .A1(B[29]), .A2(net146799), .ZN(n271) );
  NAND2_X1 U191 ( .A1(D[29]), .A2(net146793), .ZN(n270) );
  AOI22_X1 U192 ( .A1(C[29]), .A2(net146767), .B1(A[29]), .B2(net146779), .ZN(
        n269) );
  NAND4_X1 U193 ( .A1(n272), .A2(n271), .A3(n270), .A4(n269), .ZN(Y[29]) );
  NAND2_X1 U194 ( .A1(E[30]), .A2(net146817), .ZN(n276) );
  NAND2_X1 U195 ( .A1(B[30]), .A2(net146799), .ZN(n275) );
  NAND2_X1 U196 ( .A1(D[30]), .A2(net146791), .ZN(n274) );
  AOI22_X1 U197 ( .A1(C[30]), .A2(net146767), .B1(A[30]), .B2(net146777), .ZN(
        n273) );
  NAND4_X1 U198 ( .A1(n276), .A2(n275), .A3(n274), .A4(n273), .ZN(Y[30]) );
  NAND2_X1 U199 ( .A1(E[31]), .A2(net146809), .ZN(n280) );
  NAND2_X1 U200 ( .A1(B[31]), .A2(net146799), .ZN(n279) );
  NAND2_X1 U201 ( .A1(D[31]), .A2(net146789), .ZN(n278) );
  AOI22_X1 U202 ( .A1(C[31]), .A2(net146765), .B1(A[31]), .B2(net146779), .ZN(
        n277) );
  NAND4_X1 U203 ( .A1(n280), .A2(n279), .A3(n278), .A4(n277), .ZN(Y[31]) );
  NAND2_X1 U204 ( .A1(E[32]), .A2(net146817), .ZN(n284) );
  NAND2_X1 U205 ( .A1(B[32]), .A2(net146799), .ZN(n283) );
  NAND2_X1 U206 ( .A1(D[32]), .A2(net146787), .ZN(n282) );
  AOI22_X1 U207 ( .A1(C[32]), .A2(net146767), .B1(A[32]), .B2(net146779), .ZN(
        n281) );
  NAND4_X1 U208 ( .A1(n284), .A2(n283), .A3(n282), .A4(n281), .ZN(Y[32]) );
  NAND2_X1 U209 ( .A1(E[33]), .A2(net146817), .ZN(n288) );
  NAND2_X1 U210 ( .A1(B[33]), .A2(net146799), .ZN(n287) );
  NAND2_X1 U211 ( .A1(D[33]), .A2(net146785), .ZN(n286) );
  AOI22_X1 U212 ( .A1(C[33]), .A2(net146767), .B1(A[33]), .B2(net146779), .ZN(
        n285) );
  NAND4_X1 U213 ( .A1(n288), .A2(n287), .A3(n286), .A4(n285), .ZN(Y[33]) );
  NAND2_X1 U214 ( .A1(E[34]), .A2(net146817), .ZN(n292) );
  NAND2_X1 U215 ( .A1(B[34]), .A2(net146799), .ZN(n291) );
  NAND2_X1 U216 ( .A1(D[34]), .A2(net146793), .ZN(n290) );
  AOI22_X1 U217 ( .A1(C[34]), .A2(net146765), .B1(A[34]), .B2(net146777), .ZN(
        n289) );
  NAND4_X1 U218 ( .A1(n292), .A2(n291), .A3(n290), .A4(n289), .ZN(Y[34]) );
  NAND2_X1 U219 ( .A1(E[35]), .A2(net146809), .ZN(n296) );
  NAND2_X1 U220 ( .A1(B[35]), .A2(net146799), .ZN(n295) );
  NAND2_X1 U221 ( .A1(D[35]), .A2(net146791), .ZN(n294) );
  AOI22_X1 U222 ( .A1(C[35]), .A2(net146767), .B1(A[35]), .B2(net146779), .ZN(
        n293) );
  NAND4_X1 U223 ( .A1(n296), .A2(n295), .A3(n294), .A4(n293), .ZN(Y[35]) );
  NAND2_X1 U224 ( .A1(E[36]), .A2(net146813), .ZN(n300) );
  NAND2_X1 U225 ( .A1(B[36]), .A2(net146801), .ZN(n299) );
  NAND2_X1 U226 ( .A1(D[36]), .A2(net146789), .ZN(n298) );
  AOI22_X1 U227 ( .A1(C[36]), .A2(net146765), .B1(A[36]), .B2(net146779), .ZN(
        n297) );
  NAND4_X1 U228 ( .A1(n300), .A2(n299), .A3(n298), .A4(n297), .ZN(Y[36]) );
  NAND2_X1 U229 ( .A1(E[37]), .A2(net146809), .ZN(n304) );
  NAND2_X1 U230 ( .A1(B[37]), .A2(net146801), .ZN(n303) );
  NAND2_X1 U231 ( .A1(D[37]), .A2(net146787), .ZN(n302) );
  AOI22_X1 U232 ( .A1(C[37]), .A2(net146767), .B1(A[37]), .B2(net146779), .ZN(
        n301) );
  NAND4_X1 U233 ( .A1(n304), .A2(n303), .A3(n302), .A4(n301), .ZN(Y[37]) );
  NAND2_X1 U234 ( .A1(E[38]), .A2(net146817), .ZN(n308) );
  NAND2_X1 U235 ( .A1(B[38]), .A2(net146801), .ZN(n307) );
  NAND2_X1 U236 ( .A1(D[38]), .A2(net146785), .ZN(n306) );
  AOI22_X1 U237 ( .A1(C[38]), .A2(net146767), .B1(A[38]), .B2(net146777), .ZN(
        n305) );
  NAND4_X1 U238 ( .A1(n308), .A2(n307), .A3(n306), .A4(n305), .ZN(Y[38]) );
  NAND2_X1 U239 ( .A1(E[39]), .A2(net146813), .ZN(n312) );
  NAND2_X1 U240 ( .A1(B[39]), .A2(net146801), .ZN(n311) );
  NAND2_X1 U241 ( .A1(D[39]), .A2(net146793), .ZN(n310) );
  AOI22_X1 U242 ( .A1(C[39]), .A2(net146765), .B1(A[39]), .B2(net146779), .ZN(
        n309) );
  NAND4_X1 U243 ( .A1(n312), .A2(n311), .A3(n310), .A4(n309), .ZN(Y[39]) );
  NAND2_X1 U244 ( .A1(E[40]), .A2(net146809), .ZN(n316) );
  NAND2_X1 U245 ( .A1(B[40]), .A2(net146801), .ZN(n315) );
  NAND2_X1 U246 ( .A1(D[40]), .A2(net146791), .ZN(n314) );
  AOI22_X1 U247 ( .A1(C[40]), .A2(net146767), .B1(A[40]), .B2(net146779), .ZN(
        n313) );
  NAND4_X1 U248 ( .A1(n316), .A2(n315), .A3(n314), .A4(n313), .ZN(Y[40]) );
  NAND2_X1 U249 ( .A1(E[41]), .A2(net146817), .ZN(n320) );
  NAND2_X1 U250 ( .A1(B[41]), .A2(net146801), .ZN(n319) );
  NAND2_X1 U251 ( .A1(D[41]), .A2(net146789), .ZN(n318) );
  AOI22_X1 U252 ( .A1(C[41]), .A2(net146765), .B1(A[41]), .B2(net146777), .ZN(
        n317) );
  NAND4_X1 U253 ( .A1(n320), .A2(n319), .A3(n318), .A4(n317), .ZN(Y[41]) );
  NAND2_X1 U254 ( .A1(E[42]), .A2(net146813), .ZN(n324) );
  NAND2_X1 U255 ( .A1(B[42]), .A2(net146801), .ZN(n323) );
  NAND2_X1 U256 ( .A1(D[42]), .A2(net146787), .ZN(n322) );
  AOI22_X1 U257 ( .A1(C[42]), .A2(net146767), .B1(A[42]), .B2(net146779), .ZN(
        n321) );
  NAND4_X1 U258 ( .A1(n324), .A2(n323), .A3(n322), .A4(n321), .ZN(Y[42]) );
  NAND2_X1 U259 ( .A1(E[43]), .A2(net146809), .ZN(n328) );
  NAND2_X1 U260 ( .A1(B[43]), .A2(net146801), .ZN(n327) );
  NAND2_X1 U261 ( .A1(D[43]), .A2(net146785), .ZN(n326) );
  AOI22_X1 U262 ( .A1(C[43]), .A2(net146765), .B1(A[43]), .B2(net146779), .ZN(
        n325) );
  NAND4_X1 U263 ( .A1(n328), .A2(n327), .A3(n326), .A4(n325), .ZN(Y[43]) );
  NAND2_X1 U264 ( .A1(E[44]), .A2(net146813), .ZN(n332) );
  NAND2_X1 U265 ( .A1(B[44]), .A2(net146801), .ZN(n331) );
  NAND2_X1 U266 ( .A1(D[44]), .A2(net146793), .ZN(n330) );
  AOI22_X1 U267 ( .A1(C[44]), .A2(net146767), .B1(A[44]), .B2(net146779), .ZN(
        n329) );
  NAND4_X1 U268 ( .A1(n332), .A2(n331), .A3(n330), .A4(n329), .ZN(Y[44]) );
  NAND2_X1 U269 ( .A1(E[45]), .A2(net146817), .ZN(n336) );
  NAND2_X1 U270 ( .A1(B[45]), .A2(net146801), .ZN(n335) );
  NAND2_X1 U271 ( .A1(D[45]), .A2(net146791), .ZN(n334) );
  AOI22_X1 U272 ( .A1(C[45]), .A2(net146767), .B1(A[45]), .B2(net146777), .ZN(
        n333) );
  NAND4_X1 U273 ( .A1(n336), .A2(n335), .A3(n334), .A4(n333), .ZN(Y[45]) );
  NAND2_X1 U274 ( .A1(E[46]), .A2(net146809), .ZN(n340) );
  NAND2_X1 U275 ( .A1(B[46]), .A2(net146801), .ZN(n339) );
  NAND2_X1 U276 ( .A1(D[46]), .A2(net146789), .ZN(n338) );
  AOI22_X1 U277 ( .A1(C[46]), .A2(net146765), .B1(A[46]), .B2(net146779), .ZN(
        n337) );
  NAND4_X1 U278 ( .A1(n340), .A2(n339), .A3(n338), .A4(n337), .ZN(Y[46]) );
  NAND2_X1 U279 ( .A1(E[47]), .A2(net146813), .ZN(n344) );
  NAND2_X1 U280 ( .A1(B[47]), .A2(net146801), .ZN(n343) );
  NAND2_X1 U281 ( .A1(D[47]), .A2(net146787), .ZN(n342) );
  AOI22_X1 U282 ( .A1(C[47]), .A2(net146767), .B1(A[47]), .B2(net146779), .ZN(
        n341) );
  NAND4_X1 U283 ( .A1(n344), .A2(n343), .A3(n342), .A4(n341), .ZN(Y[47]) );
  NAND2_X1 U284 ( .A1(E[48]), .A2(net146817), .ZN(n348) );
  NAND2_X1 U285 ( .A1(B[48]), .A2(net146803), .ZN(n347) );
  NAND2_X1 U286 ( .A1(D[48]), .A2(net146785), .ZN(n346) );
  AOI22_X1 U287 ( .A1(C[48]), .A2(net146765), .B1(A[48]), .B2(net146779), .ZN(
        n345) );
  NAND4_X1 U288 ( .A1(n348), .A2(n347), .A3(n346), .A4(n345), .ZN(Y[48]) );
  NAND2_X1 U289 ( .A1(E[49]), .A2(net146809), .ZN(n352) );
  NAND2_X1 U290 ( .A1(B[49]), .A2(net146803), .ZN(n351) );
  NAND2_X1 U291 ( .A1(D[49]), .A2(net146793), .ZN(n350) );
  AOI22_X1 U292 ( .A1(C[49]), .A2(net146765), .B1(A[49]), .B2(net146781), .ZN(
        n349) );
  NAND4_X1 U293 ( .A1(n352), .A2(n351), .A3(n350), .A4(n349), .ZN(Y[49]) );
  NAND2_X1 U294 ( .A1(E[50]), .A2(net146811), .ZN(n356) );
  NAND2_X1 U295 ( .A1(B[50]), .A2(net146803), .ZN(n355) );
  NAND2_X1 U296 ( .A1(D[50]), .A2(net146791), .ZN(n354) );
  AOI22_X1 U297 ( .A1(C[50]), .A2(net146765), .B1(A[50]), .B2(net146777), .ZN(
        n353) );
  NAND4_X1 U298 ( .A1(n356), .A2(n355), .A3(n354), .A4(n353), .ZN(Y[50]) );
  NAND2_X1 U299 ( .A1(E[51]), .A2(net146813), .ZN(n360) );
  NAND2_X1 U300 ( .A1(B[51]), .A2(net146803), .ZN(n359) );
  NAND2_X1 U301 ( .A1(D[51]), .A2(net146789), .ZN(n358) );
  AOI22_X1 U302 ( .A1(C[51]), .A2(net146767), .B1(A[51]), .B2(net146779), .ZN(
        n357) );
  NAND4_X1 U303 ( .A1(n360), .A2(n359), .A3(n358), .A4(n357), .ZN(Y[51]) );
  NAND2_X1 U304 ( .A1(E[52]), .A2(net146817), .ZN(n364) );
  NAND2_X1 U305 ( .A1(B[52]), .A2(net146803), .ZN(n363) );
  NAND2_X1 U306 ( .A1(D[52]), .A2(net146787), .ZN(n362) );
  AOI22_X1 U307 ( .A1(C[52]), .A2(net146765), .B1(A[52]), .B2(net146779), .ZN(
        n361) );
  NAND4_X1 U308 ( .A1(n364), .A2(n363), .A3(n362), .A4(n361), .ZN(Y[52]) );
  NAND2_X1 U309 ( .A1(E[53]), .A2(net146809), .ZN(n368) );
  NAND2_X1 U310 ( .A1(B[53]), .A2(net146803), .ZN(n367) );
  NAND2_X1 U311 ( .A1(D[53]), .A2(net146785), .ZN(n366) );
  AOI22_X1 U312 ( .A1(C[53]), .A2(net146767), .B1(A[53]), .B2(net146779), .ZN(
        n365) );
  NAND4_X1 U313 ( .A1(n368), .A2(n367), .A3(n366), .A4(n365), .ZN(Y[53]) );
  NAND2_X1 U314 ( .A1(E[54]), .A2(net146811), .ZN(n372) );
  NAND2_X1 U315 ( .A1(B[54]), .A2(net146803), .ZN(n371) );
  NAND2_X1 U316 ( .A1(D[54]), .A2(net146793), .ZN(n370) );
  AOI22_X1 U317 ( .A1(C[54]), .A2(net146767), .B1(A[54]), .B2(net146781), .ZN(
        n369) );
  NAND4_X1 U318 ( .A1(n372), .A2(n371), .A3(n370), .A4(n369), .ZN(Y[54]) );
  NAND2_X1 U319 ( .A1(E[55]), .A2(net146813), .ZN(n376) );
  NAND2_X1 U320 ( .A1(B[55]), .A2(net146803), .ZN(n375) );
  NAND2_X1 U321 ( .A1(D[55]), .A2(net146791), .ZN(n374) );
  AOI22_X1 U322 ( .A1(C[55]), .A2(net146765), .B1(A[55]), .B2(net146777), .ZN(
        n373) );
  NAND4_X1 U323 ( .A1(n376), .A2(n375), .A3(n374), .A4(n373), .ZN(Y[55]) );
  NAND2_X1 U324 ( .A1(E[56]), .A2(net146817), .ZN(n380) );
  NAND2_X1 U325 ( .A1(B[56]), .A2(net146803), .ZN(n379) );
  NAND2_X1 U326 ( .A1(D[56]), .A2(net146789), .ZN(n378) );
  AOI22_X1 U327 ( .A1(C[56]), .A2(net146767), .B1(A[56]), .B2(net146779), .ZN(
        n377) );
  NAND4_X1 U328 ( .A1(n380), .A2(n379), .A3(n378), .A4(n377), .ZN(Y[56]) );
  NAND2_X1 U329 ( .A1(E[57]), .A2(net146809), .ZN(n384) );
  NAND2_X1 U330 ( .A1(B[57]), .A2(net146803), .ZN(n383) );
  NAND2_X1 U331 ( .A1(D[57]), .A2(net146787), .ZN(n382) );
  AOI22_X1 U332 ( .A1(C[57]), .A2(net146765), .B1(A[57]), .B2(net146779), .ZN(
        n381) );
  NAND4_X1 U333 ( .A1(n384), .A2(n383), .A3(n382), .A4(n381), .ZN(Y[57]) );
  NAND2_X1 U334 ( .A1(E[58]), .A2(net146811), .ZN(n388) );
  NAND2_X1 U335 ( .A1(B[58]), .A2(net146803), .ZN(n387) );
  NAND2_X1 U336 ( .A1(D[58]), .A2(net146785), .ZN(n386) );
  AOI22_X1 U337 ( .A1(C[58]), .A2(net146767), .B1(A[58]), .B2(net146779), .ZN(
        n385) );
  NAND4_X1 U338 ( .A1(n388), .A2(n387), .A3(n386), .A4(n385), .ZN(Y[58]) );
  NAND2_X1 U339 ( .A1(E[59]), .A2(net146813), .ZN(n392) );
  NAND2_X1 U340 ( .A1(B[59]), .A2(net146803), .ZN(n391) );
  NAND2_X1 U341 ( .A1(D[59]), .A2(net146793), .ZN(n390) );
  AOI22_X1 U342 ( .A1(C[59]), .A2(net146767), .B1(A[59]), .B2(net146777), .ZN(
        n389) );
  NAND4_X1 U343 ( .A1(n392), .A2(n391), .A3(n390), .A4(n389), .ZN(Y[59]) );
  NAND2_X1 U344 ( .A1(E[60]), .A2(net146813), .ZN(n396) );
  NAND2_X1 U345 ( .A1(B[60]), .A2(net146805), .ZN(n395) );
  NAND2_X1 U346 ( .A1(D[60]), .A2(net146791), .ZN(n394) );
  AOI22_X1 U347 ( .A1(C[60]), .A2(net146765), .B1(A[60]), .B2(net146781), .ZN(
        n393) );
  NAND4_X1 U348 ( .A1(n396), .A2(n395), .A3(n394), .A4(n393), .ZN(Y[60]) );
  NAND2_X1 U349 ( .A1(E[61]), .A2(net146817), .ZN(n400) );
  NAND2_X1 U350 ( .A1(B[61]), .A2(net146805), .ZN(n399) );
  NAND2_X1 U351 ( .A1(D[61]), .A2(net146789), .ZN(n398) );
  AOI22_X1 U352 ( .A1(C[61]), .A2(net146767), .B1(A[61]), .B2(net146779), .ZN(
        n397) );
  NAND4_X1 U353 ( .A1(n400), .A2(n399), .A3(n398), .A4(n397), .ZN(Y[61]) );
  NAND2_X1 U354 ( .A1(E[62]), .A2(net146809), .ZN(n404) );
  NAND2_X1 U355 ( .A1(B[62]), .A2(net146805), .ZN(n403) );
  NAND2_X1 U356 ( .A1(D[62]), .A2(net146787), .ZN(n402) );
  AOI22_X1 U357 ( .A1(C[62]), .A2(net146765), .B1(A[62]), .B2(net146777), .ZN(
        n401) );
  NAND4_X1 U358 ( .A1(n404), .A2(n403), .A3(n402), .A4(n401), .ZN(Y[62]) );
  NAND2_X1 U359 ( .A1(E[63]), .A2(net146813), .ZN(n408) );
  NAND2_X1 U360 ( .A1(B[63]), .A2(net146805), .ZN(n407) );
  NAND2_X1 U361 ( .A1(D[63]), .A2(net146785), .ZN(n406) );
  AOI22_X1 U362 ( .A1(C[63]), .A2(net146767), .B1(A[63]), .B2(net146779), .ZN(
        n405) );
  NAND4_X1 U363 ( .A1(n408), .A2(n407), .A3(n406), .A4(n405), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_14 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441;

  BUF_X2 U1 ( .A(n434), .Z(n150) );
  BUF_X2 U2 ( .A(n437), .Z(n140) );
  BUF_X2 U3 ( .A(n437), .Z(n139) );
  OR2_X2 U4 ( .A1(n176), .A2(n142), .ZN(n180) );
  NAND4_X1 U5 ( .A1(n209), .A2(n208), .A3(n207), .A4(n206), .ZN(Y[6]) );
  NAND4_X1 U6 ( .A1(n201), .A2(n200), .A3(n199), .A4(n198), .ZN(Y[4]) );
  NAND4_X1 U7 ( .A1(n213), .A2(n212), .A3(n211), .A4(n210), .ZN(Y[7]) );
  CLKBUF_X1 U8 ( .A(n436), .Z(n162) );
  BUF_X1 U9 ( .A(n436), .Z(n163) );
  BUF_X2 U10 ( .A(n436), .Z(n164) );
  INV_X1 U11 ( .A(n181), .ZN(n141) );
  CLKBUF_X1 U12 ( .A(n143), .Z(n144) );
  BUF_X2 U13 ( .A(n143), .Z(n146) );
  BUF_X2 U14 ( .A(n437), .Z(n168) );
  AND4_X2 U15 ( .A1(n178), .A2(n179), .A3(n181), .A4(n180), .ZN(n143) );
  NAND2_X1 U16 ( .A1(n177), .A2(n174), .ZN(n142) );
  CLKBUF_X1 U17 ( .A(n437), .Z(n169) );
  BUF_X1 U18 ( .A(n435), .Z(n156) );
  CLKBUF_X1 U19 ( .A(n435), .Z(n157) );
  CLKBUF_X1 U20 ( .A(n434), .Z(n151) );
  CLKBUF_X1 U21 ( .A(n143), .Z(n145) );
  CLKBUF_X1 U22 ( .A(n437), .Z(n170) );
  CLKBUF_X1 U23 ( .A(n435), .Z(n158) );
  CLKBUF_X1 U24 ( .A(n434), .Z(n152) );
  CLKBUF_X1 U25 ( .A(n437), .Z(n171) );
  CLKBUF_X1 U26 ( .A(n435), .Z(n159) );
  CLKBUF_X1 U27 ( .A(n434), .Z(n153) );
  CLKBUF_X1 U28 ( .A(n143), .Z(n147) );
  CLKBUF_X1 U29 ( .A(n141), .Z(n165) );
  CLKBUF_X1 U30 ( .A(n437), .Z(n172) );
  CLKBUF_X1 U31 ( .A(n435), .Z(n160) );
  CLKBUF_X1 U32 ( .A(n434), .Z(n154) );
  CLKBUF_X1 U33 ( .A(n143), .Z(n148) );
  CLKBUF_X1 U34 ( .A(n141), .Z(n166) );
  NAND2_X1 U35 ( .A1(n177), .A2(n175), .ZN(n181) );
  CLKBUF_X1 U36 ( .A(n143), .Z(n149) );
  CLKBUF_X1 U37 ( .A(n434), .Z(n155) );
  CLKBUF_X1 U38 ( .A(n435), .Z(n161) );
  CLKBUF_X1 U39 ( .A(n141), .Z(n167) );
  CLKBUF_X1 U40 ( .A(n437), .Z(n173) );
  INV_X1 U41 ( .A(SEL[1]), .ZN(n176) );
  INV_X1 U42 ( .A(SEL[2]), .ZN(n174) );
  NAND3_X1 U43 ( .A1(SEL[0]), .A2(n176), .A3(n174), .ZN(n178) );
  NAND3_X1 U44 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n174), .ZN(n179) );
  INV_X1 U45 ( .A(SEL[0]), .ZN(n177) );
  NOR2_X1 U46 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n175) );
  NAND2_X1 U47 ( .A1(E[0]), .A2(n144), .ZN(n185) );
  INV_X1 U48 ( .A(n178), .ZN(n434) );
  NAND2_X1 U49 ( .A1(B[0]), .A2(n150), .ZN(n184) );
  INV_X1 U50 ( .A(n179), .ZN(n435) );
  NAND2_X1 U51 ( .A1(D[0]), .A2(n156), .ZN(n183) );
  INV_X1 U52 ( .A(n180), .ZN(n437) );
  INV_X1 U53 ( .A(n181), .ZN(n436) );
  AOI22_X1 U54 ( .A1(C[0]), .A2(n168), .B1(A[0]), .B2(n162), .ZN(n182) );
  NAND4_X1 U55 ( .A1(n185), .A2(n184), .A3(n183), .A4(n182), .ZN(Y[0]) );
  NAND2_X1 U56 ( .A1(E[1]), .A2(n144), .ZN(n189) );
  NAND2_X1 U57 ( .A1(B[1]), .A2(n150), .ZN(n188) );
  NAND2_X1 U58 ( .A1(D[1]), .A2(n156), .ZN(n187) );
  AOI22_X1 U59 ( .A1(C[1]), .A2(n140), .B1(A[1]), .B2(n162), .ZN(n186) );
  NAND4_X1 U60 ( .A1(n189), .A2(n188), .A3(n187), .A4(n186), .ZN(Y[1]) );
  NAND2_X1 U61 ( .A1(E[2]), .A2(n146), .ZN(n193) );
  NAND2_X1 U62 ( .A1(B[2]), .A2(n150), .ZN(n192) );
  NAND2_X1 U63 ( .A1(D[2]), .A2(n156), .ZN(n191) );
  AOI22_X1 U64 ( .A1(C[2]), .A2(n139), .B1(A[2]), .B2(n164), .ZN(n190) );
  NAND4_X1 U65 ( .A1(n193), .A2(n192), .A3(n191), .A4(n190), .ZN(Y[2]) );
  NAND2_X1 U66 ( .A1(E[3]), .A2(n145), .ZN(n197) );
  NAND2_X1 U67 ( .A1(B[3]), .A2(n150), .ZN(n196) );
  NAND2_X1 U68 ( .A1(D[3]), .A2(n156), .ZN(n195) );
  AOI22_X1 U69 ( .A1(C[3]), .A2(n173), .B1(A[3]), .B2(n163), .ZN(n194) );
  NAND4_X1 U70 ( .A1(n197), .A2(n196), .A3(n195), .A4(n194), .ZN(Y[3]) );
  NAND2_X1 U71 ( .A1(E[4]), .A2(n149), .ZN(n201) );
  NAND2_X1 U72 ( .A1(B[4]), .A2(n150), .ZN(n200) );
  NAND2_X1 U73 ( .A1(D[4]), .A2(n156), .ZN(n199) );
  AOI22_X1 U74 ( .A1(C[4]), .A2(n172), .B1(A[4]), .B2(n164), .ZN(n198) );
  NAND2_X1 U75 ( .A1(E[5]), .A2(n148), .ZN(n205) );
  NAND2_X1 U76 ( .A1(B[5]), .A2(n150), .ZN(n204) );
  NAND2_X1 U77 ( .A1(D[5]), .A2(n156), .ZN(n203) );
  AOI22_X1 U78 ( .A1(C[5]), .A2(n171), .B1(A[5]), .B2(n163), .ZN(n202) );
  NAND4_X1 U79 ( .A1(n205), .A2(n204), .A3(n203), .A4(n202), .ZN(Y[5]) );
  NAND2_X1 U80 ( .A1(E[6]), .A2(n147), .ZN(n209) );
  NAND2_X1 U81 ( .A1(B[6]), .A2(n150), .ZN(n208) );
  NAND2_X1 U82 ( .A1(D[6]), .A2(n156), .ZN(n207) );
  AOI22_X1 U83 ( .A1(C[6]), .A2(n170), .B1(A[6]), .B2(n164), .ZN(n206) );
  NAND2_X1 U84 ( .A1(E[7]), .A2(n146), .ZN(n213) );
  NAND2_X1 U85 ( .A1(B[7]), .A2(n150), .ZN(n212) );
  NAND2_X1 U86 ( .A1(D[7]), .A2(n156), .ZN(n211) );
  AOI22_X1 U87 ( .A1(C[7]), .A2(n169), .B1(A[7]), .B2(n163), .ZN(n210) );
  NAND2_X1 U88 ( .A1(E[8]), .A2(n145), .ZN(n217) );
  NAND2_X1 U89 ( .A1(B[8]), .A2(n150), .ZN(n216) );
  NAND2_X1 U90 ( .A1(D[8]), .A2(n156), .ZN(n215) );
  AOI22_X1 U91 ( .A1(C[8]), .A2(n173), .B1(A[8]), .B2(n164), .ZN(n214) );
  NAND4_X1 U92 ( .A1(n217), .A2(n216), .A3(n215), .A4(n214), .ZN(Y[8]) );
  NAND2_X1 U93 ( .A1(E[9]), .A2(n149), .ZN(n221) );
  NAND2_X1 U94 ( .A1(B[9]), .A2(n150), .ZN(n220) );
  NAND2_X1 U95 ( .A1(D[9]), .A2(n156), .ZN(n219) );
  AOI22_X1 U96 ( .A1(C[9]), .A2(n172), .B1(A[9]), .B2(n163), .ZN(n218) );
  NAND4_X1 U97 ( .A1(n221), .A2(n220), .A3(n219), .A4(n218), .ZN(Y[9]) );
  NAND2_X1 U98 ( .A1(E[10]), .A2(n148), .ZN(n225) );
  NAND2_X1 U99 ( .A1(B[10]), .A2(n150), .ZN(n224) );
  NAND2_X1 U100 ( .A1(D[10]), .A2(n156), .ZN(n223) );
  AOI22_X1 U101 ( .A1(C[10]), .A2(n171), .B1(A[10]), .B2(n164), .ZN(n222) );
  NAND4_X1 U102 ( .A1(n225), .A2(n224), .A3(n223), .A4(n222), .ZN(Y[10]) );
  NAND2_X1 U103 ( .A1(E[11]), .A2(n147), .ZN(n229) );
  NAND2_X1 U104 ( .A1(B[11]), .A2(n150), .ZN(n228) );
  NAND2_X1 U105 ( .A1(D[11]), .A2(n156), .ZN(n227) );
  AOI22_X1 U106 ( .A1(C[11]), .A2(n170), .B1(A[11]), .B2(n163), .ZN(n226) );
  NAND4_X1 U107 ( .A1(n229), .A2(n228), .A3(n227), .A4(n226), .ZN(Y[11]) );
  NAND2_X1 U108 ( .A1(E[12]), .A2(n146), .ZN(n233) );
  NAND2_X1 U109 ( .A1(B[12]), .A2(n151), .ZN(n232) );
  NAND2_X1 U110 ( .A1(D[12]), .A2(n157), .ZN(n231) );
  AOI22_X1 U111 ( .A1(C[12]), .A2(n169), .B1(A[12]), .B2(n164), .ZN(n230) );
  NAND4_X1 U112 ( .A1(n233), .A2(n232), .A3(n231), .A4(n230), .ZN(Y[12]) );
  NAND2_X1 U113 ( .A1(E[13]), .A2(n145), .ZN(n237) );
  NAND2_X1 U114 ( .A1(B[13]), .A2(n151), .ZN(n236) );
  NAND2_X1 U115 ( .A1(D[13]), .A2(n157), .ZN(n235) );
  AOI22_X1 U116 ( .A1(C[13]), .A2(n140), .B1(A[13]), .B2(n163), .ZN(n234) );
  NAND4_X1 U117 ( .A1(n237), .A2(n236), .A3(n235), .A4(n234), .ZN(Y[13]) );
  NAND2_X1 U118 ( .A1(E[14]), .A2(n149), .ZN(n241) );
  NAND2_X1 U119 ( .A1(B[14]), .A2(n151), .ZN(n240) );
  NAND2_X1 U120 ( .A1(D[14]), .A2(n157), .ZN(n239) );
  AOI22_X1 U121 ( .A1(C[14]), .A2(n139), .B1(A[14]), .B2(n164), .ZN(n238) );
  NAND4_X1 U122 ( .A1(n241), .A2(n240), .A3(n239), .A4(n238), .ZN(Y[14]) );
  NAND2_X1 U123 ( .A1(E[15]), .A2(n148), .ZN(n245) );
  NAND2_X1 U124 ( .A1(B[15]), .A2(n151), .ZN(n244) );
  NAND2_X1 U125 ( .A1(D[15]), .A2(n157), .ZN(n243) );
  AOI22_X1 U126 ( .A1(C[15]), .A2(n140), .B1(A[15]), .B2(n163), .ZN(n242) );
  NAND4_X1 U127 ( .A1(n245), .A2(n244), .A3(n243), .A4(n242), .ZN(Y[15]) );
  NAND2_X1 U128 ( .A1(E[16]), .A2(n147), .ZN(n249) );
  NAND2_X1 U129 ( .A1(B[16]), .A2(n151), .ZN(n248) );
  NAND2_X1 U130 ( .A1(D[16]), .A2(n157), .ZN(n247) );
  AOI22_X1 U131 ( .A1(C[16]), .A2(n139), .B1(A[16]), .B2(n164), .ZN(n246) );
  NAND4_X1 U132 ( .A1(n249), .A2(n248), .A3(n247), .A4(n246), .ZN(Y[16]) );
  NAND2_X1 U133 ( .A1(E[17]), .A2(n146), .ZN(n253) );
  NAND2_X1 U134 ( .A1(B[17]), .A2(n151), .ZN(n252) );
  NAND2_X1 U135 ( .A1(D[17]), .A2(n157), .ZN(n251) );
  AOI22_X1 U136 ( .A1(C[17]), .A2(n173), .B1(A[17]), .B2(n163), .ZN(n250) );
  NAND4_X1 U137 ( .A1(n253), .A2(n252), .A3(n251), .A4(n250), .ZN(Y[17]) );
  NAND2_X1 U138 ( .A1(E[18]), .A2(n145), .ZN(n257) );
  NAND2_X1 U139 ( .A1(B[18]), .A2(n151), .ZN(n256) );
  NAND2_X1 U140 ( .A1(D[18]), .A2(n157), .ZN(n255) );
  AOI22_X1 U141 ( .A1(C[18]), .A2(n172), .B1(A[18]), .B2(n164), .ZN(n254) );
  NAND4_X1 U142 ( .A1(n257), .A2(n256), .A3(n255), .A4(n254), .ZN(Y[18]) );
  NAND2_X1 U143 ( .A1(E[19]), .A2(n149), .ZN(n261) );
  NAND2_X1 U144 ( .A1(B[19]), .A2(n151), .ZN(n260) );
  NAND2_X1 U145 ( .A1(D[19]), .A2(n157), .ZN(n259) );
  AOI22_X1 U146 ( .A1(C[19]), .A2(n171), .B1(A[19]), .B2(n163), .ZN(n258) );
  NAND4_X1 U147 ( .A1(n261), .A2(n260), .A3(n259), .A4(n258), .ZN(Y[19]) );
  NAND2_X1 U148 ( .A1(E[20]), .A2(n148), .ZN(n265) );
  NAND2_X1 U149 ( .A1(B[20]), .A2(n151), .ZN(n264) );
  NAND2_X1 U150 ( .A1(D[20]), .A2(n157), .ZN(n263) );
  AOI22_X1 U151 ( .A1(C[20]), .A2(n170), .B1(A[20]), .B2(n164), .ZN(n262) );
  NAND4_X1 U152 ( .A1(n265), .A2(n264), .A3(n263), .A4(n262), .ZN(Y[20]) );
  NAND2_X1 U153 ( .A1(E[21]), .A2(n147), .ZN(n269) );
  NAND2_X1 U154 ( .A1(B[21]), .A2(n151), .ZN(n268) );
  NAND2_X1 U155 ( .A1(D[21]), .A2(n157), .ZN(n267) );
  AOI22_X1 U156 ( .A1(C[21]), .A2(n169), .B1(A[21]), .B2(n163), .ZN(n266) );
  NAND4_X1 U157 ( .A1(n269), .A2(n268), .A3(n267), .A4(n266), .ZN(Y[21]) );
  NAND2_X1 U158 ( .A1(E[22]), .A2(n146), .ZN(n273) );
  NAND2_X1 U159 ( .A1(B[22]), .A2(n151), .ZN(n272) );
  NAND2_X1 U160 ( .A1(D[22]), .A2(n157), .ZN(n271) );
  AOI22_X1 U161 ( .A1(C[22]), .A2(n140), .B1(A[22]), .B2(n164), .ZN(n270) );
  NAND4_X1 U162 ( .A1(n273), .A2(n272), .A3(n271), .A4(n270), .ZN(Y[22]) );
  NAND2_X1 U163 ( .A1(E[23]), .A2(n145), .ZN(n277) );
  NAND2_X1 U164 ( .A1(B[23]), .A2(n151), .ZN(n276) );
  NAND2_X1 U165 ( .A1(D[23]), .A2(n157), .ZN(n275) );
  AOI22_X1 U166 ( .A1(C[23]), .A2(n140), .B1(A[23]), .B2(n163), .ZN(n274) );
  NAND4_X1 U167 ( .A1(n277), .A2(n276), .A3(n275), .A4(n274), .ZN(Y[23]) );
  NAND2_X1 U168 ( .A1(E[24]), .A2(n149), .ZN(n281) );
  NAND2_X1 U169 ( .A1(B[24]), .A2(n152), .ZN(n280) );
  NAND2_X1 U170 ( .A1(D[24]), .A2(n158), .ZN(n279) );
  AOI22_X1 U171 ( .A1(C[24]), .A2(n140), .B1(A[24]), .B2(n164), .ZN(n278) );
  NAND4_X1 U172 ( .A1(n281), .A2(n280), .A3(n279), .A4(n278), .ZN(Y[24]) );
  NAND2_X1 U173 ( .A1(E[25]), .A2(n148), .ZN(n285) );
  NAND2_X1 U174 ( .A1(B[25]), .A2(n152), .ZN(n284) );
  NAND2_X1 U175 ( .A1(D[25]), .A2(n158), .ZN(n283) );
  AOI22_X1 U176 ( .A1(C[25]), .A2(n139), .B1(A[25]), .B2(n163), .ZN(n282) );
  NAND4_X1 U177 ( .A1(n285), .A2(n284), .A3(n283), .A4(n282), .ZN(Y[25]) );
  NAND2_X1 U178 ( .A1(E[26]), .A2(n147), .ZN(n289) );
  NAND2_X1 U179 ( .A1(B[26]), .A2(n152), .ZN(n288) );
  NAND2_X1 U180 ( .A1(D[26]), .A2(n158), .ZN(n287) );
  AOI22_X1 U181 ( .A1(C[26]), .A2(n139), .B1(A[26]), .B2(n164), .ZN(n286) );
  NAND4_X1 U182 ( .A1(n289), .A2(n288), .A3(n287), .A4(n286), .ZN(Y[26]) );
  NAND2_X1 U183 ( .A1(E[27]), .A2(n146), .ZN(n293) );
  NAND2_X1 U184 ( .A1(B[27]), .A2(n152), .ZN(n292) );
  NAND2_X1 U185 ( .A1(D[27]), .A2(n158), .ZN(n291) );
  AOI22_X1 U186 ( .A1(C[27]), .A2(n139), .B1(A[27]), .B2(n163), .ZN(n290) );
  NAND4_X1 U187 ( .A1(n293), .A2(n292), .A3(n291), .A4(n290), .ZN(Y[27]) );
  NAND2_X1 U188 ( .A1(E[28]), .A2(n145), .ZN(n297) );
  NAND2_X1 U189 ( .A1(B[28]), .A2(n152), .ZN(n296) );
  NAND2_X1 U190 ( .A1(D[28]), .A2(n158), .ZN(n295) );
  AOI22_X1 U191 ( .A1(C[28]), .A2(n140), .B1(A[28]), .B2(n164), .ZN(n294) );
  NAND4_X1 U192 ( .A1(n297), .A2(n296), .A3(n295), .A4(n294), .ZN(Y[28]) );
  NAND2_X1 U193 ( .A1(E[29]), .A2(n149), .ZN(n301) );
  NAND2_X1 U194 ( .A1(B[29]), .A2(n152), .ZN(n300) );
  NAND2_X1 U195 ( .A1(D[29]), .A2(n158), .ZN(n299) );
  AOI22_X1 U196 ( .A1(C[29]), .A2(n139), .B1(A[29]), .B2(n163), .ZN(n298) );
  NAND4_X1 U197 ( .A1(n301), .A2(n300), .A3(n299), .A4(n298), .ZN(Y[29]) );
  NAND2_X1 U198 ( .A1(E[30]), .A2(n148), .ZN(n305) );
  NAND2_X1 U199 ( .A1(B[30]), .A2(n152), .ZN(n304) );
  NAND2_X1 U200 ( .A1(D[30]), .A2(n158), .ZN(n303) );
  AOI22_X1 U201 ( .A1(C[30]), .A2(n140), .B1(A[30]), .B2(n164), .ZN(n302) );
  NAND4_X1 U202 ( .A1(n305), .A2(n304), .A3(n303), .A4(n302), .ZN(Y[30]) );
  NAND2_X1 U203 ( .A1(E[31]), .A2(n147), .ZN(n309) );
  NAND2_X1 U204 ( .A1(B[31]), .A2(n152), .ZN(n308) );
  NAND2_X1 U205 ( .A1(D[31]), .A2(n158), .ZN(n307) );
  AOI22_X1 U206 ( .A1(C[31]), .A2(n139), .B1(A[31]), .B2(n163), .ZN(n306) );
  NAND4_X1 U207 ( .A1(n309), .A2(n308), .A3(n307), .A4(n306), .ZN(Y[31]) );
  NAND2_X1 U208 ( .A1(E[32]), .A2(n146), .ZN(n313) );
  NAND2_X1 U209 ( .A1(B[32]), .A2(n152), .ZN(n312) );
  NAND2_X1 U210 ( .A1(D[32]), .A2(n158), .ZN(n311) );
  AOI22_X1 U211 ( .A1(C[32]), .A2(n173), .B1(A[32]), .B2(n164), .ZN(n310) );
  NAND4_X1 U212 ( .A1(n313), .A2(n312), .A3(n311), .A4(n310), .ZN(Y[32]) );
  NAND2_X1 U213 ( .A1(E[33]), .A2(n145), .ZN(n317) );
  NAND2_X1 U214 ( .A1(B[33]), .A2(n152), .ZN(n316) );
  NAND2_X1 U215 ( .A1(D[33]), .A2(n158), .ZN(n315) );
  AOI22_X1 U216 ( .A1(C[33]), .A2(n172), .B1(A[33]), .B2(n163), .ZN(n314) );
  NAND4_X1 U217 ( .A1(n317), .A2(n316), .A3(n315), .A4(n314), .ZN(Y[33]) );
  NAND2_X1 U218 ( .A1(E[34]), .A2(n149), .ZN(n321) );
  NAND2_X1 U219 ( .A1(B[34]), .A2(n152), .ZN(n320) );
  NAND2_X1 U220 ( .A1(D[34]), .A2(n158), .ZN(n319) );
  AOI22_X1 U221 ( .A1(C[34]), .A2(n171), .B1(A[34]), .B2(n164), .ZN(n318) );
  NAND4_X1 U222 ( .A1(n321), .A2(n320), .A3(n319), .A4(n318), .ZN(Y[34]) );
  NAND2_X1 U223 ( .A1(E[35]), .A2(n148), .ZN(n325) );
  NAND2_X1 U224 ( .A1(B[35]), .A2(n152), .ZN(n324) );
  NAND2_X1 U225 ( .A1(D[35]), .A2(n158), .ZN(n323) );
  AOI22_X1 U226 ( .A1(C[35]), .A2(n170), .B1(A[35]), .B2(n163), .ZN(n322) );
  NAND4_X1 U227 ( .A1(n325), .A2(n324), .A3(n323), .A4(n322), .ZN(Y[35]) );
  NAND2_X1 U228 ( .A1(E[36]), .A2(n147), .ZN(n329) );
  NAND2_X1 U229 ( .A1(B[36]), .A2(n153), .ZN(n328) );
  NAND2_X1 U230 ( .A1(D[36]), .A2(n159), .ZN(n327) );
  AOI22_X1 U231 ( .A1(C[36]), .A2(n169), .B1(A[36]), .B2(n165), .ZN(n326) );
  NAND4_X1 U232 ( .A1(n329), .A2(n328), .A3(n327), .A4(n326), .ZN(Y[36]) );
  NAND2_X1 U233 ( .A1(E[37]), .A2(n146), .ZN(n333) );
  NAND2_X1 U234 ( .A1(B[37]), .A2(n153), .ZN(n332) );
  NAND2_X1 U235 ( .A1(D[37]), .A2(n159), .ZN(n331) );
  AOI22_X1 U236 ( .A1(C[37]), .A2(n140), .B1(A[37]), .B2(n165), .ZN(n330) );
  NAND4_X1 U237 ( .A1(n333), .A2(n332), .A3(n331), .A4(n330), .ZN(Y[37]) );
  NAND2_X1 U238 ( .A1(E[38]), .A2(n145), .ZN(n337) );
  NAND2_X1 U239 ( .A1(B[38]), .A2(n153), .ZN(n336) );
  NAND2_X1 U240 ( .A1(D[38]), .A2(n159), .ZN(n335) );
  AOI22_X1 U241 ( .A1(C[38]), .A2(n139), .B1(A[38]), .B2(n165), .ZN(n334) );
  NAND4_X1 U242 ( .A1(n337), .A2(n336), .A3(n335), .A4(n334), .ZN(Y[38]) );
  NAND2_X1 U243 ( .A1(E[39]), .A2(n149), .ZN(n341) );
  NAND2_X1 U244 ( .A1(B[39]), .A2(n153), .ZN(n340) );
  NAND2_X1 U245 ( .A1(D[39]), .A2(n159), .ZN(n339) );
  AOI22_X1 U246 ( .A1(C[39]), .A2(n140), .B1(A[39]), .B2(n165), .ZN(n338) );
  NAND4_X1 U247 ( .A1(n341), .A2(n340), .A3(n339), .A4(n338), .ZN(Y[39]) );
  NAND2_X1 U248 ( .A1(E[40]), .A2(n148), .ZN(n345) );
  NAND2_X1 U249 ( .A1(B[40]), .A2(n153), .ZN(n344) );
  NAND2_X1 U250 ( .A1(D[40]), .A2(n159), .ZN(n343) );
  AOI22_X1 U251 ( .A1(C[40]), .A2(n139), .B1(A[40]), .B2(n165), .ZN(n342) );
  NAND4_X1 U252 ( .A1(n345), .A2(n344), .A3(n343), .A4(n342), .ZN(Y[40]) );
  NAND2_X1 U253 ( .A1(E[41]), .A2(n147), .ZN(n349) );
  NAND2_X1 U254 ( .A1(B[41]), .A2(n153), .ZN(n348) );
  NAND2_X1 U255 ( .A1(D[41]), .A2(n159), .ZN(n347) );
  AOI22_X1 U256 ( .A1(C[41]), .A2(n173), .B1(A[41]), .B2(n165), .ZN(n346) );
  NAND4_X1 U257 ( .A1(n349), .A2(n348), .A3(n347), .A4(n346), .ZN(Y[41]) );
  NAND2_X1 U258 ( .A1(E[42]), .A2(n146), .ZN(n353) );
  NAND2_X1 U259 ( .A1(B[42]), .A2(n153), .ZN(n352) );
  NAND2_X1 U260 ( .A1(D[42]), .A2(n159), .ZN(n351) );
  AOI22_X1 U261 ( .A1(C[42]), .A2(n172), .B1(A[42]), .B2(n165), .ZN(n350) );
  NAND4_X1 U262 ( .A1(n353), .A2(n352), .A3(n351), .A4(n350), .ZN(Y[42]) );
  NAND2_X1 U263 ( .A1(E[43]), .A2(n145), .ZN(n357) );
  NAND2_X1 U264 ( .A1(B[43]), .A2(n153), .ZN(n356) );
  NAND2_X1 U265 ( .A1(D[43]), .A2(n159), .ZN(n355) );
  AOI22_X1 U266 ( .A1(C[43]), .A2(n171), .B1(A[43]), .B2(n165), .ZN(n354) );
  NAND4_X1 U267 ( .A1(n357), .A2(n356), .A3(n355), .A4(n354), .ZN(Y[43]) );
  NAND2_X1 U268 ( .A1(E[44]), .A2(n149), .ZN(n361) );
  NAND2_X1 U269 ( .A1(B[44]), .A2(n153), .ZN(n360) );
  NAND2_X1 U270 ( .A1(D[44]), .A2(n159), .ZN(n359) );
  AOI22_X1 U271 ( .A1(C[44]), .A2(n170), .B1(A[44]), .B2(n165), .ZN(n358) );
  NAND4_X1 U272 ( .A1(n361), .A2(n360), .A3(n359), .A4(n358), .ZN(Y[44]) );
  NAND2_X1 U273 ( .A1(E[45]), .A2(n148), .ZN(n365) );
  NAND2_X1 U274 ( .A1(B[45]), .A2(n153), .ZN(n364) );
  NAND2_X1 U275 ( .A1(D[45]), .A2(n159), .ZN(n363) );
  AOI22_X1 U276 ( .A1(C[45]), .A2(n169), .B1(A[45]), .B2(n165), .ZN(n362) );
  NAND4_X1 U277 ( .A1(n365), .A2(n364), .A3(n363), .A4(n362), .ZN(Y[45]) );
  NAND2_X1 U278 ( .A1(E[46]), .A2(n147), .ZN(n369) );
  NAND2_X1 U279 ( .A1(B[46]), .A2(n153), .ZN(n368) );
  NAND2_X1 U280 ( .A1(D[46]), .A2(n159), .ZN(n367) );
  AOI22_X1 U281 ( .A1(C[46]), .A2(n140), .B1(A[46]), .B2(n165), .ZN(n366) );
  NAND4_X1 U282 ( .A1(n369), .A2(n368), .A3(n367), .A4(n366), .ZN(Y[46]) );
  NAND2_X1 U283 ( .A1(E[47]), .A2(n146), .ZN(n373) );
  NAND2_X1 U284 ( .A1(B[47]), .A2(n153), .ZN(n372) );
  NAND2_X1 U285 ( .A1(D[47]), .A2(n159), .ZN(n371) );
  AOI22_X1 U286 ( .A1(C[47]), .A2(n139), .B1(A[47]), .B2(n165), .ZN(n370) );
  NAND4_X1 U287 ( .A1(n373), .A2(n372), .A3(n371), .A4(n370), .ZN(Y[47]) );
  NAND2_X1 U288 ( .A1(E[48]), .A2(n145), .ZN(n377) );
  NAND2_X1 U289 ( .A1(B[48]), .A2(n154), .ZN(n376) );
  NAND2_X1 U290 ( .A1(D[48]), .A2(n160), .ZN(n375) );
  AOI22_X1 U291 ( .A1(C[48]), .A2(n140), .B1(A[48]), .B2(n166), .ZN(n374) );
  NAND4_X1 U292 ( .A1(n377), .A2(n376), .A3(n375), .A4(n374), .ZN(Y[48]) );
  NAND2_X1 U293 ( .A1(E[49]), .A2(n149), .ZN(n381) );
  NAND2_X1 U294 ( .A1(B[49]), .A2(n154), .ZN(n380) );
  NAND2_X1 U295 ( .A1(D[49]), .A2(n160), .ZN(n379) );
  AOI22_X1 U296 ( .A1(C[49]), .A2(n139), .B1(A[49]), .B2(n166), .ZN(n378) );
  NAND4_X1 U297 ( .A1(n381), .A2(n380), .A3(n379), .A4(n378), .ZN(Y[49]) );
  NAND2_X1 U298 ( .A1(E[50]), .A2(n148), .ZN(n385) );
  NAND2_X1 U299 ( .A1(B[50]), .A2(n154), .ZN(n384) );
  NAND2_X1 U300 ( .A1(D[50]), .A2(n160), .ZN(n383) );
  AOI22_X1 U301 ( .A1(C[50]), .A2(n140), .B1(A[50]), .B2(n166), .ZN(n382) );
  NAND4_X1 U302 ( .A1(n385), .A2(n384), .A3(n383), .A4(n382), .ZN(Y[50]) );
  NAND2_X1 U303 ( .A1(E[51]), .A2(n147), .ZN(n389) );
  NAND2_X1 U304 ( .A1(B[51]), .A2(n154), .ZN(n388) );
  NAND2_X1 U305 ( .A1(D[51]), .A2(n160), .ZN(n387) );
  AOI22_X1 U306 ( .A1(C[51]), .A2(n139), .B1(A[51]), .B2(n166), .ZN(n386) );
  NAND4_X1 U307 ( .A1(n389), .A2(n388), .A3(n387), .A4(n386), .ZN(Y[51]) );
  NAND2_X1 U308 ( .A1(E[52]), .A2(n146), .ZN(n393) );
  NAND2_X1 U309 ( .A1(B[52]), .A2(n154), .ZN(n392) );
  NAND2_X1 U310 ( .A1(D[52]), .A2(n160), .ZN(n391) );
  AOI22_X1 U311 ( .A1(C[52]), .A2(n173), .B1(A[52]), .B2(n166), .ZN(n390) );
  NAND4_X1 U312 ( .A1(n393), .A2(n392), .A3(n391), .A4(n390), .ZN(Y[52]) );
  NAND2_X1 U313 ( .A1(E[53]), .A2(n145), .ZN(n397) );
  NAND2_X1 U314 ( .A1(B[53]), .A2(n154), .ZN(n396) );
  NAND2_X1 U315 ( .A1(D[53]), .A2(n160), .ZN(n395) );
  AOI22_X1 U316 ( .A1(C[53]), .A2(n172), .B1(A[53]), .B2(n166), .ZN(n394) );
  NAND4_X1 U317 ( .A1(n397), .A2(n396), .A3(n395), .A4(n394), .ZN(Y[53]) );
  NAND2_X1 U318 ( .A1(E[54]), .A2(n149), .ZN(n401) );
  NAND2_X1 U319 ( .A1(B[54]), .A2(n154), .ZN(n400) );
  NAND2_X1 U320 ( .A1(D[54]), .A2(n160), .ZN(n399) );
  AOI22_X1 U321 ( .A1(C[54]), .A2(n171), .B1(A[54]), .B2(n166), .ZN(n398) );
  NAND4_X1 U322 ( .A1(n401), .A2(n400), .A3(n399), .A4(n398), .ZN(Y[54]) );
  NAND2_X1 U323 ( .A1(E[55]), .A2(n148), .ZN(n405) );
  NAND2_X1 U324 ( .A1(B[55]), .A2(n154), .ZN(n404) );
  NAND2_X1 U325 ( .A1(D[55]), .A2(n160), .ZN(n403) );
  AOI22_X1 U326 ( .A1(C[55]), .A2(n170), .B1(A[55]), .B2(n166), .ZN(n402) );
  NAND4_X1 U327 ( .A1(n405), .A2(n404), .A3(n403), .A4(n402), .ZN(Y[55]) );
  NAND2_X1 U328 ( .A1(E[56]), .A2(n147), .ZN(n409) );
  NAND2_X1 U329 ( .A1(B[56]), .A2(n154), .ZN(n408) );
  NAND2_X1 U330 ( .A1(D[56]), .A2(n160), .ZN(n407) );
  AOI22_X1 U331 ( .A1(C[56]), .A2(n169), .B1(A[56]), .B2(n166), .ZN(n406) );
  NAND4_X1 U332 ( .A1(n409), .A2(n408), .A3(n407), .A4(n406), .ZN(Y[56]) );
  NAND2_X1 U333 ( .A1(E[57]), .A2(n146), .ZN(n413) );
  NAND2_X1 U334 ( .A1(B[57]), .A2(n154), .ZN(n412) );
  NAND2_X1 U335 ( .A1(D[57]), .A2(n160), .ZN(n411) );
  AOI22_X1 U336 ( .A1(C[57]), .A2(n173), .B1(A[57]), .B2(n166), .ZN(n410) );
  NAND4_X1 U337 ( .A1(n413), .A2(n412), .A3(n411), .A4(n410), .ZN(Y[57]) );
  NAND2_X1 U338 ( .A1(E[58]), .A2(n145), .ZN(n417) );
  NAND2_X1 U339 ( .A1(B[58]), .A2(n154), .ZN(n416) );
  NAND2_X1 U340 ( .A1(D[58]), .A2(n160), .ZN(n415) );
  AOI22_X1 U341 ( .A1(C[58]), .A2(n172), .B1(A[58]), .B2(n166), .ZN(n414) );
  NAND4_X1 U342 ( .A1(n417), .A2(n416), .A3(n415), .A4(n414), .ZN(Y[58]) );
  NAND2_X1 U343 ( .A1(E[59]), .A2(n149), .ZN(n421) );
  NAND2_X1 U344 ( .A1(B[59]), .A2(n154), .ZN(n420) );
  NAND2_X1 U345 ( .A1(D[59]), .A2(n160), .ZN(n419) );
  AOI22_X1 U346 ( .A1(C[59]), .A2(n171), .B1(A[59]), .B2(n166), .ZN(n418) );
  NAND4_X1 U347 ( .A1(n421), .A2(n420), .A3(n419), .A4(n418), .ZN(Y[59]) );
  NAND2_X1 U348 ( .A1(E[60]), .A2(n148), .ZN(n425) );
  NAND2_X1 U349 ( .A1(B[60]), .A2(n155), .ZN(n424) );
  NAND2_X1 U350 ( .A1(D[60]), .A2(n161), .ZN(n423) );
  AOI22_X1 U351 ( .A1(C[60]), .A2(n170), .B1(A[60]), .B2(n167), .ZN(n422) );
  NAND4_X1 U352 ( .A1(n425), .A2(n424), .A3(n423), .A4(n422), .ZN(Y[60]) );
  NAND2_X1 U353 ( .A1(E[61]), .A2(n147), .ZN(n429) );
  NAND2_X1 U354 ( .A1(B[61]), .A2(n155), .ZN(n428) );
  NAND2_X1 U355 ( .A1(D[61]), .A2(n161), .ZN(n427) );
  AOI22_X1 U356 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n167), .ZN(n426) );
  NAND4_X1 U357 ( .A1(n429), .A2(n428), .A3(n427), .A4(n426), .ZN(Y[61]) );
  NAND2_X1 U358 ( .A1(E[62]), .A2(n146), .ZN(n433) );
  NAND2_X1 U359 ( .A1(B[62]), .A2(n155), .ZN(n432) );
  NAND2_X1 U360 ( .A1(D[62]), .A2(n161), .ZN(n431) );
  AOI22_X1 U361 ( .A1(C[62]), .A2(n140), .B1(A[62]), .B2(n167), .ZN(n430) );
  NAND4_X1 U362 ( .A1(n433), .A2(n432), .A3(n431), .A4(n430), .ZN(Y[62]) );
  NAND2_X1 U363 ( .A1(E[63]), .A2(n145), .ZN(n441) );
  NAND2_X1 U364 ( .A1(B[63]), .A2(n155), .ZN(n440) );
  NAND2_X1 U365 ( .A1(D[63]), .A2(n161), .ZN(n439) );
  AOI22_X1 U366 ( .A1(C[63]), .A2(n139), .B1(A[63]), .B2(n167), .ZN(n438) );
  NAND4_X1 U367 ( .A1(n441), .A2(n440), .A3(n439), .A4(n438), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_13 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X1 U1 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND4_X2 U2 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND4_X2 U3 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND4_X2 U4 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND4_X2 U5 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  BUF_X2 U6 ( .A(n434), .Z(n164) );
  CLKBUF_X1 U7 ( .A(n434), .Z(n165) );
  BUF_X2 U8 ( .A(n432), .Z(n152) );
  BUF_X2 U9 ( .A(n431), .Z(n146) );
  BUF_X2 U10 ( .A(n139), .Z(n140) );
  CLKBUF_X1 U11 ( .A(n139), .Z(n141) );
  BUF_X2 U12 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U13 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U14 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U15 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U16 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U17 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U18 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U19 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U20 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U21 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U22 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U23 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U24 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U25 ( .A(n433), .Z(n161) );
  CLKBUF_X1 U26 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U27 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U28 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U29 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U30 ( .A(n433), .Z(n162) );
  AND4_X1 U31 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U32 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U33 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U34 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U35 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U36 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U37 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U38 ( .A(n434), .Z(n169) );
  INV_X1 U39 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U40 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U41 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U42 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U43 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U44 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U45 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U46 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U47 ( .A(n175), .ZN(n431) );
  NAND2_X1 U48 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U49 ( .A(n176), .ZN(n432) );
  NAND2_X1 U50 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U51 ( .A(n177), .ZN(n434) );
  INV_X1 U52 ( .A(n178), .ZN(n433) );
  AOI22_X1 U53 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U54 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U55 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U56 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U57 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U58 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U59 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U60 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U61 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U62 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U63 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U64 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U65 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U66 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U67 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U68 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U69 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U70 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U71 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U72 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U73 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U74 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U75 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U76 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U77 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U78 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND2_X1 U79 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U80 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U81 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U82 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND2_X1 U83 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U84 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U85 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U86 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND2_X1 U87 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U88 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U89 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U90 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U91 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U92 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U93 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U94 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U95 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND2_X1 U96 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U97 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U98 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U99 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U100 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U101 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U102 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U103 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U104 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND2_X1 U105 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U106 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U107 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U108 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U109 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U110 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U111 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U112 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U113 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U114 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U115 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U116 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U117 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U118 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U119 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U120 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U121 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U122 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U123 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U124 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U125 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U126 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U127 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U128 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U129 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U130 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U131 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U132 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U133 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U134 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U135 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U136 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U137 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U138 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U139 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U140 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U141 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U142 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U143 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U144 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U145 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U146 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U147 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U148 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U149 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U150 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U151 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U152 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U153 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U154 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U155 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U156 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U157 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U158 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U159 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U160 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U161 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U162 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U163 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U164 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U165 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U166 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U167 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U168 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U169 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U170 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U171 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U172 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U173 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U174 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U175 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U176 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U177 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U178 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U179 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U180 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U181 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U182 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U183 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U184 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U185 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U186 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U187 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U188 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U189 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U190 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U191 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U192 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U193 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U194 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U195 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U196 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U197 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U198 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U199 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U200 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U201 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U202 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U203 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U204 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U205 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U206 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U207 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U208 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U209 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U210 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U211 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U212 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U213 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U214 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U215 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U216 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U217 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U218 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U219 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U220 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U221 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U222 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U223 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U224 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U225 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U226 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U227 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U228 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U229 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U230 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U231 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U232 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U233 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U234 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U235 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U236 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U237 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U238 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U239 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U240 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U241 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U242 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U243 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U244 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U245 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U246 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U247 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U248 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U249 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U250 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U251 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U252 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U253 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U254 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U255 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U256 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U257 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U258 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U259 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U260 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U261 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U262 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U263 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U264 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U265 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U266 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U267 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U268 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U269 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U270 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U271 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U272 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U273 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U274 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U275 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U276 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U277 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U278 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U279 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U280 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U281 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U282 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U283 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U284 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U285 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U286 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U287 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U288 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U289 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U290 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U291 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U292 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U293 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U294 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U295 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U296 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U297 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U298 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U299 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U300 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U301 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U302 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U303 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U304 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U305 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U306 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U307 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U308 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U309 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U310 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U311 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U312 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U313 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U314 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U315 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U316 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U317 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U318 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U319 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U320 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U321 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U322 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U323 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U324 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U325 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U326 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U327 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U328 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U329 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U330 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U331 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U332 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U333 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U334 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U335 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U336 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U337 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U338 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U339 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U340 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U341 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U342 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U343 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U344 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U345 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U346 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U347 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U348 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U349 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U350 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U351 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U352 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U353 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND4_X1 U354 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND2_X1 U355 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U356 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U357 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U358 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND4_X1 U359 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_12 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X2 U1 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND4_X2 U2 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  BUF_X1 U3 ( .A(n434), .Z(n164) );
  BUF_X1 U4 ( .A(n432), .Z(n152) );
  BUF_X1 U5 ( .A(n431), .Z(n146) );
  BUF_X1 U6 ( .A(n139), .Z(n140) );
  BUF_X1 U7 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U8 ( .A(n434), .Z(n165) );
  CLKBUF_X1 U9 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U10 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U11 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U12 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U13 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U14 ( .A(n139), .Z(n141) );
  CLKBUF_X1 U15 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U16 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U17 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U18 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U19 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U20 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U21 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U22 ( .A(n433), .Z(n161) );
  CLKBUF_X1 U23 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U24 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U25 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U26 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U27 ( .A(n433), .Z(n162) );
  AND4_X1 U28 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U29 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U30 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U31 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U32 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U33 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U34 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U35 ( .A(n434), .Z(n169) );
  INV_X1 U36 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U37 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U38 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U39 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U40 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U41 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U42 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U43 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U44 ( .A(n175), .ZN(n431) );
  NAND2_X1 U45 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U46 ( .A(n176), .ZN(n432) );
  NAND2_X1 U47 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U48 ( .A(n177), .ZN(n434) );
  INV_X1 U49 ( .A(n178), .ZN(n433) );
  AOI22_X1 U50 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U51 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U52 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U53 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U54 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U55 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND2_X1 U56 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U57 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U58 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U59 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U60 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U61 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U62 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U63 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U64 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U65 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U66 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U67 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U68 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U69 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U70 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U71 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U72 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U73 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U74 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U75 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U76 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U77 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U78 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U79 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U80 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U81 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U82 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U83 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U84 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND4_X1 U85 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  NAND2_X1 U86 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U87 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U88 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U89 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND2_X1 U90 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U91 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U92 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U93 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U94 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U95 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U96 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U97 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U98 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U99 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U100 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U101 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U102 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U103 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND4_X1 U104 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND2_X1 U105 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U106 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U107 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U108 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U109 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U110 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U111 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U112 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U113 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U114 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U115 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U116 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U117 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U118 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U119 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U120 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U121 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U122 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U123 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U124 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U125 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U126 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U127 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U128 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U129 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U130 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U131 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U132 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U133 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U134 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U135 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U136 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U137 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U138 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U139 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U140 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U141 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U142 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U143 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U144 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U145 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U146 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U147 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U148 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U149 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U150 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U151 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U152 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U153 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U154 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U155 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U156 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U157 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U158 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U159 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U160 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U161 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U162 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U163 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U164 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U165 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U166 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U167 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U168 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U169 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U170 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U171 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U172 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U173 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U174 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U175 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U176 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U177 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U178 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U179 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U180 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U181 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U182 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U183 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U184 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U185 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U186 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U187 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U188 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U189 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U190 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U191 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U192 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U193 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U194 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U195 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U196 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U197 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U198 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U199 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U200 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U201 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U202 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U203 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U204 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U205 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U206 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U207 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U208 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U209 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U210 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U211 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U212 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U213 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U214 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U215 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U216 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U217 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U218 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U219 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U220 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U221 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U222 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U223 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U224 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U225 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U226 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U227 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U228 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U229 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U230 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U231 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U232 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U233 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U234 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U235 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U236 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U237 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U238 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U239 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U240 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U241 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U242 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U243 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U244 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U245 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U246 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U247 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U248 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U249 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U250 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U251 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U252 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U253 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U254 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U255 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U256 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U257 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U258 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U259 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U260 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U261 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U262 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U263 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U264 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U265 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U266 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U267 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U268 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U269 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U270 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U271 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U272 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U273 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U274 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U275 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U276 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U277 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U278 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U279 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U280 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U281 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U282 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U283 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U284 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U285 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U286 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U287 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U288 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U289 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U290 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U291 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U292 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U293 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U294 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U295 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U296 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U297 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U298 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U299 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U300 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U301 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U302 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U303 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U304 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U305 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U306 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U307 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U308 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U309 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U310 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U311 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U312 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U313 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U314 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U315 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U316 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U317 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U318 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U319 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U320 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U321 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U322 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U323 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U324 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U325 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U326 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U327 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U328 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U329 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U330 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U331 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U332 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U333 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U334 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U335 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U336 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U337 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U338 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U339 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U340 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U341 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U342 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U343 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U344 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U345 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U346 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U347 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U348 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U349 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U350 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U351 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U352 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U353 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND4_X1 U354 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND2_X1 U355 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U356 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U357 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U358 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND4_X1 U359 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_11 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X2 U1 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND4_X2 U2 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND4_X2 U3 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND4_X2 U4 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  BUF_X2 U5 ( .A(n434), .Z(n164) );
  BUF_X2 U6 ( .A(n432), .Z(n152) );
  BUF_X1 U7 ( .A(n431), .Z(n146) );
  BUF_X1 U8 ( .A(n139), .Z(n140) );
  BUF_X1 U9 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U10 ( .A(n434), .Z(n165) );
  CLKBUF_X1 U11 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U12 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U13 ( .A(n139), .Z(n141) );
  CLKBUF_X1 U14 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U15 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U16 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U17 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U18 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U19 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U20 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U21 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U22 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U23 ( .A(n433), .Z(n161) );
  CLKBUF_X1 U24 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U25 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U26 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U27 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U28 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U29 ( .A(n433), .Z(n162) );
  AND4_X1 U30 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U31 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U32 ( .A1(n174), .A2(n171), .ZN(n178) );
  NAND4_X1 U33 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  CLKBUF_X1 U34 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U35 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U36 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U37 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U38 ( .A(n434), .Z(n169) );
  INV_X1 U39 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U40 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U41 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U42 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U43 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U44 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U45 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U46 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U47 ( .A(n175), .ZN(n431) );
  NAND2_X1 U48 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U49 ( .A(n176), .ZN(n432) );
  NAND2_X1 U50 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U51 ( .A(n177), .ZN(n434) );
  INV_X1 U52 ( .A(n178), .ZN(n433) );
  AOI22_X1 U53 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U54 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U55 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U56 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U57 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U58 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U59 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U60 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U61 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U62 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U63 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND2_X1 U64 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U65 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U66 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U67 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND2_X1 U68 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U69 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U70 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U71 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U72 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U73 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U74 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U75 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U76 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U77 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U78 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U79 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U80 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U81 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND2_X1 U82 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U83 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U84 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U85 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND4_X1 U86 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  NAND2_X1 U87 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U88 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U89 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U90 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U91 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U92 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U93 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U94 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U95 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND2_X1 U96 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U97 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U98 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U99 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND2_X1 U100 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U101 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U102 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U103 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND4_X1 U104 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND2_X1 U105 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U106 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U107 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U108 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U109 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U110 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U111 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U112 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U113 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U114 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U115 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U116 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U117 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U118 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U119 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U120 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U121 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U122 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U123 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U124 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U125 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U126 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U127 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U128 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U129 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U130 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U131 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U132 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U133 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U134 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U135 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U136 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U137 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U138 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U139 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U140 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U141 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U142 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U143 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U144 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U145 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U146 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U147 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U148 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U149 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U150 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U151 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U152 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U153 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U154 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U155 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U156 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U157 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U158 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U159 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U160 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U161 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U162 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U163 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U164 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U165 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U166 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U167 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U168 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U169 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U170 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U171 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U172 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U173 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U174 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U175 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U176 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U177 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U178 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U179 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U180 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U181 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U182 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U183 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U184 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U185 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U186 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U187 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U188 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U189 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U190 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U191 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U192 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U193 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U194 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U195 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U196 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U197 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U198 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U199 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U200 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U201 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U202 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U203 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U204 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U205 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U206 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U207 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U208 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U209 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U210 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U211 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U212 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U213 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U214 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U215 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U216 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U217 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U218 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U219 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U220 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U221 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U222 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U223 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U224 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U225 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U226 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U227 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U228 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U229 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U230 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U231 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U232 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U233 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U234 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U235 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U236 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U237 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U238 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U239 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U240 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U241 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U242 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U243 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U244 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U245 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U246 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U247 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U248 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U249 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U250 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U251 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U252 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U253 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U254 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U255 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U256 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U257 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U258 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U259 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U260 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U261 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U262 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U263 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U264 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U265 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U266 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U267 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U268 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U269 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U270 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U271 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U272 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U273 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U274 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U275 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U276 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U277 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U278 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U279 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U280 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U281 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U282 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U283 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U284 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U285 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U286 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U287 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U288 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U289 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U290 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U291 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U292 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U293 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U294 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U295 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U296 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U297 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U298 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U299 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U300 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U301 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U302 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U303 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U304 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U305 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U306 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U307 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U308 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U309 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U310 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U311 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U312 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U313 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U314 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U315 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U316 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U317 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U318 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U319 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U320 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U321 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U322 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U323 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U324 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U325 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U326 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U327 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U328 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U329 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U330 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U331 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U332 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U333 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U334 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U335 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U336 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U337 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U338 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U339 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U340 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U341 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U342 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U343 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U344 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U345 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U346 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U347 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U348 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U349 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U350 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U351 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U352 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U353 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND4_X1 U354 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND2_X1 U355 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U356 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U357 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U358 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND4_X1 U359 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_10 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X2 U1 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND4_X2 U2 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  BUF_X2 U3 ( .A(n431), .Z(n146) );
  BUF_X2 U4 ( .A(n434), .Z(n164) );
  BUF_X2 U5 ( .A(n432), .Z(n152) );
  BUF_X1 U6 ( .A(n139), .Z(n140) );
  BUF_X1 U7 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U8 ( .A(n434), .Z(n165) );
  CLKBUF_X1 U9 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U10 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U11 ( .A(n139), .Z(n141) );
  CLKBUF_X1 U12 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U13 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U14 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U15 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U16 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U17 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U18 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U19 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U20 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U21 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U22 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U23 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U24 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U25 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U26 ( .A(n433), .Z(n162) );
  CLKBUF_X1 U27 ( .A(n433), .Z(n161) );
  AND4_X1 U28 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U29 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U30 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U31 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U32 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U33 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U34 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U35 ( .A(n434), .Z(n169) );
  INV_X1 U36 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U37 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U38 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U39 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U40 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U41 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U42 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U43 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U44 ( .A(n175), .ZN(n431) );
  NAND2_X1 U45 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U46 ( .A(n176), .ZN(n432) );
  NAND2_X1 U47 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U48 ( .A(n177), .ZN(n434) );
  INV_X1 U49 ( .A(n178), .ZN(n433) );
  AOI22_X1 U50 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U51 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U52 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U53 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U54 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U55 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND2_X1 U56 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U57 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U58 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U59 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U60 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U61 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U62 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U63 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U64 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U65 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U66 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U67 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U68 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U69 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U70 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U71 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U72 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U73 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U74 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U75 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U76 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U77 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U78 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U79 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U80 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U81 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U82 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U83 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U84 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND4_X1 U85 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  NAND2_X1 U86 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U87 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U88 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U89 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U90 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U91 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U92 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U93 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U94 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U95 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U96 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U97 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U98 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U99 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U100 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U101 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U102 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U103 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U104 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND4_X1 U105 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND2_X1 U106 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U107 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U108 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U109 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U110 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U111 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U112 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U113 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U114 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U115 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U116 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U117 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U118 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U119 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U120 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U121 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U122 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U123 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U124 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U125 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U126 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U127 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U128 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U129 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U130 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U131 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U132 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U133 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U134 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U135 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U136 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U137 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U138 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U139 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U140 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U141 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U142 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U143 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U144 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U145 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U146 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U147 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U148 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U149 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U150 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U151 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U152 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U153 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U154 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U155 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U156 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U157 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U158 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U159 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U160 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U161 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U162 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U163 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U164 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U165 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U166 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U167 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U168 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U169 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U170 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U171 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U172 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U173 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U174 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U175 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U176 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U177 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U178 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U179 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U180 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U181 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U182 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U183 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U184 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U185 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U186 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U187 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U188 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U189 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U190 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U191 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U192 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U193 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U194 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U195 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U196 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U197 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U198 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U199 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U200 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U201 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U202 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U203 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U204 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U205 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U206 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U207 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U208 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U209 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U210 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U211 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U212 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U213 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U214 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U215 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U216 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U217 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U218 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U219 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U220 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U221 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U222 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U223 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U224 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U225 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U226 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U227 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U228 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U229 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U230 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U231 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U232 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U233 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U234 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U235 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U236 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U237 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U238 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U239 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U240 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U241 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U242 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U243 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U244 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U245 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U246 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U247 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U248 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U249 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U250 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U251 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U252 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U253 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U254 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U255 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U256 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U257 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U258 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U259 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U260 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U261 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U262 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U263 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U264 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U265 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U266 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U267 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U268 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U269 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U270 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U271 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U272 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U273 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U274 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U275 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U276 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U277 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U278 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U279 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U280 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U281 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U282 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U283 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U284 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U285 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U286 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U287 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U288 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U289 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U290 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U291 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U292 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U293 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U294 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U295 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U296 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U297 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U298 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U299 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U300 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U301 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U302 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U303 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U304 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U305 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U306 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U307 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U308 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U309 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U310 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U311 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U312 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U313 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U314 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U315 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U316 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U317 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U318 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U319 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U320 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U321 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U322 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U323 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U324 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U325 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U326 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U327 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U328 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U329 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U330 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U331 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U332 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U333 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U334 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U335 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U336 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U337 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U338 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U339 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U340 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U341 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U342 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U343 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U344 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U345 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U346 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U347 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U348 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U349 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND2_X1 U350 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U351 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U352 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U353 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND4_X1 U354 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND2_X1 U355 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U356 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U357 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U358 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND4_X1 U359 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_9 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X2 U1 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND4_X2 U2 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND4_X2 U3 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND4_X2 U4 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND4_X2 U5 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  BUF_X2 U6 ( .A(n434), .Z(n164) );
  BUF_X2 U7 ( .A(n432), .Z(n152) );
  BUF_X2 U8 ( .A(n431), .Z(n146) );
  BUF_X2 U9 ( .A(n139), .Z(n140) );
  BUF_X2 U10 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U11 ( .A(n434), .Z(n165) );
  CLKBUF_X1 U12 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U13 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U14 ( .A(n139), .Z(n141) );
  CLKBUF_X1 U15 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U16 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U17 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U18 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U19 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U20 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U21 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U22 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U23 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U24 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U25 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U26 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U27 ( .A(n433), .Z(n162) );
  CLKBUF_X1 U28 ( .A(n433), .Z(n161) );
  CLKBUF_X1 U29 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U30 ( .A(n431), .Z(n150) );
  AND4_X1 U31 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U32 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U33 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U34 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U35 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U36 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U37 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U38 ( .A(n434), .Z(n169) );
  INV_X1 U39 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U40 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U41 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U42 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U43 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U44 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U45 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U46 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U47 ( .A(n175), .ZN(n431) );
  NAND2_X1 U48 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U49 ( .A(n176), .ZN(n432) );
  NAND2_X1 U50 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U51 ( .A(n177), .ZN(n434) );
  INV_X1 U52 ( .A(n178), .ZN(n433) );
  AOI22_X1 U53 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U54 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U55 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U56 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U57 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U58 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U59 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U60 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U61 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U62 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U63 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND2_X1 U64 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U65 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U66 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U67 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U68 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U69 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U70 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U71 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U72 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND2_X1 U73 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U74 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U75 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U76 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U77 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U78 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U79 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U80 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U81 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U82 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U83 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U84 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U85 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U86 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND2_X1 U87 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U88 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U89 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U90 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U91 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U92 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U93 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U94 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U95 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U96 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U97 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U98 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U99 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U100 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U101 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U102 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U103 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U104 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U105 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND2_X1 U106 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U107 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U108 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U109 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U110 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U111 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U112 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U113 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U114 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U115 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U116 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U117 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U118 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U119 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U120 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U121 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U122 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U123 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U124 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U125 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U126 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U127 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U128 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U129 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U130 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U131 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U132 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U133 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U134 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U135 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U136 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U137 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U138 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U139 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U140 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U141 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U142 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U143 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U144 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U145 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U146 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U147 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U148 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U149 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U150 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U151 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U152 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U153 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U154 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U155 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U156 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U157 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U158 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U159 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U160 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U161 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U162 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U163 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U164 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U165 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U166 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U167 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U168 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U169 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U170 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U171 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U172 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U173 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U174 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U175 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U176 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U177 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U178 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U179 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U180 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U181 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U182 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U183 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U184 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U185 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U186 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U187 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U188 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U189 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U190 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U191 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U192 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U193 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U194 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U195 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U196 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U197 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U198 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U199 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U200 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U201 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U202 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U203 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U204 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U205 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U206 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U207 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U208 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U209 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U210 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U211 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U212 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U213 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U214 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U215 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U216 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U217 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U218 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U219 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U220 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U221 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U222 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U223 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U224 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U225 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U226 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U227 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U228 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U229 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U230 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U231 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U232 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U233 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U234 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U235 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U236 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U237 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U238 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U239 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U240 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U241 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U242 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U243 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U244 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U245 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U246 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U247 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U248 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U249 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U250 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U251 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U252 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U253 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U254 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U255 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U256 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U257 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U258 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U259 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U260 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U261 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U262 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U263 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U264 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U265 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U266 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U267 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U268 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U269 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U270 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U271 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U272 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U273 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U274 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U275 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U276 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U277 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U278 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U279 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U280 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U281 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U282 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U283 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U284 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U285 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U286 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U287 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U288 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U289 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U290 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U291 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U292 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U293 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U294 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U295 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U296 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U297 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U298 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U299 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U300 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U301 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U302 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U303 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U304 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U305 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U306 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U307 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U308 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U309 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U310 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U311 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U312 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U313 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U314 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U315 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U316 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U317 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U318 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U319 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U320 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U321 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U322 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U323 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U324 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U325 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U326 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U327 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U328 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U329 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U330 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U331 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U332 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U333 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U334 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U335 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U336 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U337 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U338 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U339 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U340 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U341 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U342 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U343 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U344 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U345 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U346 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U347 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U348 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U349 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U350 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U351 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U352 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U353 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U354 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND4_X1 U355 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND2_X1 U356 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U357 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U358 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U359 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_8 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  AND4_X1 U1 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  BUF_X2 U2 ( .A(n139), .Z(n140) );
  BUF_X2 U3 ( .A(n434), .Z(n164) );
  CLKBUF_X1 U4 ( .A(n434), .Z(n165) );
  BUF_X2 U5 ( .A(n432), .Z(n152) );
  CLKBUF_X1 U6 ( .A(n432), .Z(n153) );
  BUF_X2 U7 ( .A(n431), .Z(n146) );
  CLKBUF_X1 U8 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U9 ( .A(n139), .Z(n141) );
  BUF_X2 U10 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U11 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U12 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U13 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U14 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U15 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U16 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U17 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U18 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U19 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U20 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U21 ( .A(n433), .Z(n161) );
  CLKBUF_X1 U22 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U23 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U24 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U25 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U26 ( .A(n433), .Z(n162) );
  NAND2_X1 U27 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U28 ( .A1(n174), .A2(n171), .ZN(n178) );
  NAND4_X1 U29 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  CLKBUF_X1 U30 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U31 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U32 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U33 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U34 ( .A(n434), .Z(n169) );
  INV_X1 U35 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U36 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U37 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U38 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U39 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U40 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U41 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U42 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U43 ( .A(n175), .ZN(n431) );
  NAND2_X1 U44 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U45 ( .A(n176), .ZN(n432) );
  NAND2_X1 U46 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U47 ( .A(n177), .ZN(n434) );
  INV_X1 U48 ( .A(n178), .ZN(n433) );
  AOI22_X1 U49 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U50 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U51 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U52 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U53 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U54 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U55 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U56 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U57 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U58 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U59 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U60 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U61 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U62 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U63 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U64 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U65 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U66 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U67 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U68 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U69 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U70 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U71 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U72 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U73 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U74 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U75 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U76 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U77 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U78 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U79 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U80 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U81 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U82 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U83 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U84 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND4_X1 U85 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  NAND2_X1 U86 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U87 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U88 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U89 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U90 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U91 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U92 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U93 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U94 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U95 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U96 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U97 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U98 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U99 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U100 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U101 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U102 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U103 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U104 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND4_X1 U105 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND2_X1 U106 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U107 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U108 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U109 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U110 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U111 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U112 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U113 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U114 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U115 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U116 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U117 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U118 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U119 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U120 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U121 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U122 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U123 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U124 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U125 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U126 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U127 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U128 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U129 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U130 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U131 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U132 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U133 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U134 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U135 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U136 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U137 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U138 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U139 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U140 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U141 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U142 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U143 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U144 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U145 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U146 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U147 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U148 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U149 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U150 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U151 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U152 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U153 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U154 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U155 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U156 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U157 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U158 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U159 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U160 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U161 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U162 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U163 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U164 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U165 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U166 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U167 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U168 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U169 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U170 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U171 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U172 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U173 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U174 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U175 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U176 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U177 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U178 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U179 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U180 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U181 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U182 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U183 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U184 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U185 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U186 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U187 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U188 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U189 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U190 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U191 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U192 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U193 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U194 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U195 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U196 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U197 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U198 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U199 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U200 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U201 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U202 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U203 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U204 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U205 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U206 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U207 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U208 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U209 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U210 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U211 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U212 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U213 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U214 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U215 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U216 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U217 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U218 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U219 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U220 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U221 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U222 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U223 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U224 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U225 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U226 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U227 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U228 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U229 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U230 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U231 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U232 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U233 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U234 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U235 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U236 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U237 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U238 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U239 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U240 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U241 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U242 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U243 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U244 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U245 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U246 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U247 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U248 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U249 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U250 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U251 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U252 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U253 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U254 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U255 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U256 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U257 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U258 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U259 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U260 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U261 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U262 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U263 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U264 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND2_X1 U265 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U266 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U267 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U268 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U269 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U270 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U271 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U272 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U273 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U274 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U275 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U276 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U277 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U278 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U279 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U280 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U281 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U282 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U283 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U284 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U285 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U286 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U287 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U288 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U289 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U290 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U291 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U292 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U293 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U294 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U295 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U296 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U297 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U298 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U299 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U300 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U301 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U302 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U303 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U304 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U305 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U306 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U307 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U308 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U309 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U310 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U311 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U312 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U313 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U314 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U315 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U316 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U317 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U318 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U319 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U320 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U321 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U322 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U323 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U324 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U325 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U326 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U327 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U328 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U329 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U330 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U331 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U332 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U333 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U334 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U335 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U336 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U337 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U338 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U339 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U340 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U341 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U342 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U343 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U344 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U345 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U346 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U347 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U348 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U349 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U350 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U351 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U352 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U353 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND4_X1 U354 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND2_X1 U355 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U356 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U357 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U358 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND4_X1 U359 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_7 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X2 U1 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND4_X2 U2 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  BUF_X2 U3 ( .A(n434), .Z(n164) );
  CLKBUF_X1 U4 ( .A(n434), .Z(n165) );
  BUF_X2 U5 ( .A(n432), .Z(n152) );
  BUF_X2 U6 ( .A(n431), .Z(n146) );
  BUF_X2 U7 ( .A(n139), .Z(n140) );
  CLKBUF_X1 U8 ( .A(n139), .Z(n141) );
  BUF_X2 U9 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U10 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U11 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U12 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U13 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U14 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U15 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U16 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U17 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U18 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U19 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U20 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U21 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U22 ( .A(n433), .Z(n161) );
  CLKBUF_X1 U23 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U24 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U25 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U26 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U27 ( .A(n433), .Z(n162) );
  AND4_X1 U28 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U29 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U30 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U31 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U32 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U33 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U34 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U35 ( .A(n434), .Z(n169) );
  INV_X1 U36 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U37 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U38 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U39 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U40 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U41 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U42 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U43 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U44 ( .A(n175), .ZN(n431) );
  NAND2_X1 U45 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U46 ( .A(n176), .ZN(n432) );
  NAND2_X1 U47 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U48 ( .A(n177), .ZN(n434) );
  INV_X1 U49 ( .A(n178), .ZN(n433) );
  AOI22_X1 U50 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U51 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U52 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U53 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U54 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U55 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U56 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U57 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U58 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U59 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U60 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U61 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U62 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U63 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U64 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U65 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U66 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U67 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U68 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U69 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U70 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND2_X1 U71 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U72 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U73 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U74 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U75 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U76 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U77 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U78 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U79 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U80 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U81 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U82 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U83 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U84 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND4_X1 U85 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  NAND2_X1 U86 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U87 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U88 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U89 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U90 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U91 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U92 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U93 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U94 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U95 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U96 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U97 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U98 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U99 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U100 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U101 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U102 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U103 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U104 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND4_X1 U105 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND2_X1 U106 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U107 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U108 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U109 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U110 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U111 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U112 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U113 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U114 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U115 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U116 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U117 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U118 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U119 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U120 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U121 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U122 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U123 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U124 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U125 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U126 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U127 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U128 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U129 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U130 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U131 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U132 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U133 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U134 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U135 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U136 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U137 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U138 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U139 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U140 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U141 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U142 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U143 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U144 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U145 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U146 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U147 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U148 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U149 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U150 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U151 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U152 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U153 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U154 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U155 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U156 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U157 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U158 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U159 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U160 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U161 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U162 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U163 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U164 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U165 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U166 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U167 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U168 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U169 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U170 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U171 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U172 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U173 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U174 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U175 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U176 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U177 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U178 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U179 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U180 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U181 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U182 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U183 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U184 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U185 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U186 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U187 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U188 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U189 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U190 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U191 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U192 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U193 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U194 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U195 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U196 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U197 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U198 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U199 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U200 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U201 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U202 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U203 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U204 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U205 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U206 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U207 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U208 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U209 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U210 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U211 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U212 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U213 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U214 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U215 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U216 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U217 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U218 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U219 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U220 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U221 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U222 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U223 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U224 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U225 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U226 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U227 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U228 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U229 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U230 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U231 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U232 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U233 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U234 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U235 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U236 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U237 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U238 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U239 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U240 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U241 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U242 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U243 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U244 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U245 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U246 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U247 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U248 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U249 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U250 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U251 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U252 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U253 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U254 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U255 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U256 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U257 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U258 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U259 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U260 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U261 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U262 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U263 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U264 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U265 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U266 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U267 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U268 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U269 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U270 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U271 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U272 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U273 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U274 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U275 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U276 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U277 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U278 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U279 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U280 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U281 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U282 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U283 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U284 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U285 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U286 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U287 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U288 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U289 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U290 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U291 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U292 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U293 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U294 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U295 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U296 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U297 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U298 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U299 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U300 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U301 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U302 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U303 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U304 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U305 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U306 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U307 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U308 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U309 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U310 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U311 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U312 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U313 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U314 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U315 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U316 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U317 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U318 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U319 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U320 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U321 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U322 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U323 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U324 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U325 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U326 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U327 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U328 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U329 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U330 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U331 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U332 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U333 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U334 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U335 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U336 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U337 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U338 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U339 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U340 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U341 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U342 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U343 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U344 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U345 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U346 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U347 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U348 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U349 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U350 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U351 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U352 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U353 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U354 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND4_X1 U355 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND2_X1 U356 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U357 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U358 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U359 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_6 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X2 U1 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND4_X2 U2 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND4_X2 U3 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  BUF_X2 U4 ( .A(n434), .Z(n164) );
  BUF_X2 U5 ( .A(n432), .Z(n152) );
  BUF_X2 U6 ( .A(n431), .Z(n146) );
  BUF_X2 U7 ( .A(n139), .Z(n140) );
  BUF_X2 U8 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U9 ( .A(n434), .Z(n165) );
  CLKBUF_X1 U10 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U11 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U12 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U13 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U14 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U15 ( .A(n139), .Z(n141) );
  CLKBUF_X1 U16 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U17 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U18 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U19 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U20 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U21 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U22 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U23 ( .A(n433), .Z(n161) );
  CLKBUF_X1 U24 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U25 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U26 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U27 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U28 ( .A(n433), .Z(n162) );
  AND4_X1 U29 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U30 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U31 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U32 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U33 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U34 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U35 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U36 ( .A(n434), .Z(n169) );
  INV_X1 U37 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U38 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U39 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U40 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U41 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U43 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U44 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U45 ( .A(n175), .ZN(n431) );
  NAND2_X1 U46 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U47 ( .A(n176), .ZN(n432) );
  NAND2_X1 U48 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U49 ( .A(n177), .ZN(n434) );
  INV_X1 U50 ( .A(n178), .ZN(n433) );
  AOI22_X1 U51 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U52 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U53 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U54 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U55 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U56 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U57 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U58 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U59 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U60 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U61 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U62 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U63 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U64 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U65 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U66 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U67 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U68 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U69 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U70 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U71 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U72 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U73 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U74 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U75 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U76 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U77 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U78 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U79 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U80 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U81 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U82 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U83 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U84 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U85 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U86 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND4_X1 U87 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  NAND2_X1 U88 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U89 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U90 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U91 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U92 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U93 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U94 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U95 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U96 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U97 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U98 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U99 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U100 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U101 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U102 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U103 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U104 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U105 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U106 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND2_X1 U107 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U108 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U109 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U110 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U111 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U112 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U113 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U114 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U115 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U116 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U117 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U118 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U119 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U120 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U121 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U122 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U123 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U124 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U125 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U126 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U127 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U128 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U129 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U130 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U131 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U132 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U133 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U134 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U135 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U136 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U137 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U138 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U139 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U140 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U141 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U142 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U143 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U144 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U145 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U146 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U147 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U148 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U149 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U150 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U151 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U152 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U153 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U154 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U155 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U156 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U157 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U158 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U159 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U160 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U161 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U162 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U163 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U164 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U165 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U166 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U167 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U168 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U169 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U170 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U171 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U172 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U173 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U174 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U175 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U176 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U177 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U178 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U179 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U180 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U181 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U182 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U183 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U184 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U185 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U186 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U187 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U188 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U189 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U190 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U191 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U192 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U193 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U194 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U195 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U196 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U197 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U198 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U199 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U200 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U201 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U202 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U203 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U204 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U205 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U206 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U207 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U208 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U209 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U210 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U211 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U212 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U213 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U214 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U215 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U216 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U217 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U218 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U219 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U220 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U221 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U222 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U223 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U224 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U225 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U226 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U227 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U228 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U229 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U230 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U231 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U232 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U233 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U234 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U235 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U236 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U237 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U238 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U239 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U240 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U241 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U242 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U243 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U244 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U245 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U246 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U247 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U248 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U249 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U250 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U251 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U252 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U253 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U254 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U255 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U256 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U257 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U258 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U259 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U260 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U261 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U262 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U263 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U264 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U265 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U266 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U267 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U268 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U269 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U270 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U271 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U272 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U273 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U274 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U275 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U276 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U277 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U278 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U279 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U280 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U281 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U282 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U283 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U284 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U285 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U286 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U287 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U288 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U289 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U290 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U291 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U292 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U293 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U294 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U295 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U296 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U297 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U298 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U299 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U300 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U301 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U302 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U303 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U304 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U305 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U306 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U307 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U308 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U309 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U310 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U311 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U312 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U313 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U314 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U315 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U316 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U317 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U318 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U319 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U320 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U321 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U322 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U323 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U324 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U325 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U326 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U327 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U328 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U329 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U330 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U331 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U332 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U333 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U334 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U335 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U336 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U337 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U338 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U339 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U340 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U341 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U342 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U343 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U344 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U345 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U346 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U347 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U348 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U349 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U350 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U351 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U352 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U353 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U354 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U355 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND2_X1 U356 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U357 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U358 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U359 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_5 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X2 U1 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND4_X2 U2 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  BUF_X2 U3 ( .A(n434), .Z(n164) );
  BUF_X2 U4 ( .A(n432), .Z(n152) );
  BUF_X2 U5 ( .A(n431), .Z(n146) );
  BUF_X2 U6 ( .A(n139), .Z(n140) );
  BUF_X2 U7 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U8 ( .A(n434), .Z(n165) );
  CLKBUF_X1 U9 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U10 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U11 ( .A(n139), .Z(n141) );
  CLKBUF_X1 U12 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U13 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U14 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U15 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U16 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U17 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U18 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U19 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U20 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U21 ( .A(n433), .Z(n161) );
  CLKBUF_X1 U22 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U23 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U24 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U25 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U26 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U27 ( .A(n433), .Z(n162) );
  AND4_X1 U28 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U29 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U30 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U31 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U32 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U33 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U34 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U35 ( .A(n434), .Z(n169) );
  INV_X1 U36 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U37 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U38 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U39 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U40 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U41 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U42 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U43 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U44 ( .A(n175), .ZN(n431) );
  NAND2_X1 U45 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U46 ( .A(n176), .ZN(n432) );
  NAND2_X1 U47 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U48 ( .A(n177), .ZN(n434) );
  INV_X1 U49 ( .A(n178), .ZN(n433) );
  AOI22_X1 U50 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U51 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U52 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U53 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U54 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U55 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U56 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U57 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U58 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U59 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U60 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U61 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U62 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U63 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U64 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U65 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U66 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U67 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U68 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U69 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U70 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U71 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U72 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U73 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U74 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U75 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U76 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U77 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U78 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U79 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U80 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U81 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U82 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U83 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U84 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U85 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND2_X1 U86 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U87 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U88 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U89 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U90 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U91 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U92 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U93 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U94 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U95 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U96 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U97 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U98 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U99 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND2_X1 U100 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U101 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U102 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U103 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND4_X1 U104 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND2_X1 U105 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U106 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U107 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U108 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U109 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U110 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U111 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U112 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U113 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U114 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U115 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U116 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U117 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U118 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U119 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U120 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U121 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U122 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U123 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U124 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U125 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U126 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U127 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U128 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U129 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U130 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U131 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U132 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U133 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U134 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U135 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U136 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U137 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U138 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U139 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U140 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U141 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U142 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U143 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U144 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U145 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U146 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U147 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U148 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U149 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U150 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U151 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U152 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U153 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U154 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U155 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U156 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U157 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U158 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U159 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U160 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U161 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U162 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U163 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U164 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U165 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U166 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U167 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U168 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U169 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U170 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U171 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U172 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U173 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U174 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U175 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U176 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U177 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U178 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U179 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U180 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U181 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U182 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U183 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U184 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U185 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U186 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U187 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U188 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U189 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U190 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U191 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U192 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U193 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U194 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U195 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U196 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U197 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U198 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U199 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U200 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U201 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U202 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U203 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U204 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U205 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U206 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U207 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U208 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U209 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U210 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U211 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U212 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U213 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U214 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U215 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U216 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U217 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U218 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U219 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U220 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U221 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U222 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U223 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U224 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U225 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U226 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U227 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U228 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U229 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U230 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U231 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U232 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U233 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U234 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U235 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U236 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U237 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U238 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U239 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U240 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U241 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U242 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U243 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U244 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U245 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U246 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U247 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U248 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U249 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U250 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U251 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U252 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U253 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U254 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U255 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U256 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U257 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U258 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U259 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U260 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U261 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U262 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U263 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U264 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U265 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U266 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U267 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U268 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U269 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U270 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U271 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U272 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U273 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U274 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U275 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U276 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U277 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U278 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U279 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U280 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U281 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U282 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U283 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U284 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U285 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U286 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U287 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U288 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U289 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U290 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U291 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U292 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U293 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U294 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U295 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U296 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U297 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U298 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U299 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U300 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U301 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U302 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U303 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U304 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U305 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U306 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U307 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U308 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U309 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U310 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U311 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U312 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U313 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U314 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U315 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U316 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U317 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U318 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U319 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U320 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U321 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U322 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U323 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U324 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U325 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U326 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U327 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U328 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U329 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U330 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U331 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U332 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U333 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U334 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U335 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U336 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U337 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U338 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U339 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U340 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U341 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U342 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U343 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U344 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U345 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U346 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U347 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U348 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U349 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U350 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U351 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U352 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U353 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND4_X1 U354 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND2_X1 U355 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U356 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U357 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U358 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND4_X1 U359 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_4 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X1 U1 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND4_X2 U2 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND4_X2 U3 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  AND4_X1 U4 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  BUF_X2 U5 ( .A(n434), .Z(n164) );
  BUF_X2 U6 ( .A(n432), .Z(n152) );
  BUF_X2 U7 ( .A(n431), .Z(n146) );
  BUF_X2 U8 ( .A(n139), .Z(n140) );
  BUF_X2 U9 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U10 ( .A(n434), .Z(n165) );
  CLKBUF_X1 U11 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U12 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U13 ( .A(n139), .Z(n141) );
  CLKBUF_X1 U14 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U15 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U16 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U17 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U18 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U19 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U20 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U21 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U22 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U23 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U24 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U25 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U26 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U27 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U28 ( .A(n433), .Z(n162) );
  CLKBUF_X1 U29 ( .A(n433), .Z(n161) );
  NAND2_X1 U30 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U31 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U32 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U33 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U34 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U35 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U36 ( .A(n434), .Z(n169) );
  INV_X1 U37 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U38 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U39 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U40 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U41 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U42 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U43 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U44 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U45 ( .A(n175), .ZN(n431) );
  NAND2_X1 U46 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U47 ( .A(n176), .ZN(n432) );
  NAND2_X1 U48 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U49 ( .A(n177), .ZN(n434) );
  INV_X1 U50 ( .A(n178), .ZN(n433) );
  AOI22_X1 U51 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U52 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U53 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U54 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U55 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U56 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U57 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U58 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U59 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U60 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U61 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U62 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U63 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U64 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U65 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U66 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U67 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U68 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U69 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U70 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U71 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U72 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U73 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U74 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U75 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U76 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U77 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U78 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U79 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U80 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U81 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U82 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U83 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U84 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U85 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U86 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND4_X1 U87 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  NAND2_X1 U88 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U89 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U90 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U91 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND2_X1 U92 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U93 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U94 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U95 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U96 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U97 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U98 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U99 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U100 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U101 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U102 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U103 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U104 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U105 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND2_X1 U106 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U107 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U108 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U109 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U110 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U111 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U112 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U113 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U114 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U115 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U116 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U117 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U118 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U119 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U120 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U121 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U122 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U123 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U124 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U125 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U126 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U127 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U128 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U129 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U130 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U131 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U132 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U133 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U134 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U135 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U136 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U137 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U138 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U139 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U140 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U141 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U142 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U143 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U144 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U145 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U146 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U147 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U148 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U149 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U150 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U151 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U152 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U153 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U154 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U155 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U156 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U157 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U158 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U159 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U160 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U161 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U162 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U163 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U164 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U165 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U166 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U167 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U168 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U169 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U170 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U171 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U172 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U173 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U174 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U175 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U176 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U177 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U178 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U179 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U180 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U181 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U182 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U183 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U184 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U185 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U186 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U187 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U188 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U189 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U190 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U191 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U192 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U193 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U194 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U195 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U196 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U197 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U198 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U199 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U200 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U201 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U202 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U203 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U204 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U205 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U206 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U207 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U208 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U209 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U210 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U211 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U212 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U213 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U214 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U215 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U216 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U217 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U218 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U219 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U220 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U221 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U222 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U223 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U224 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U225 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U226 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U227 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U228 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U229 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U230 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U231 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U232 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U233 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U234 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U235 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U236 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U237 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U238 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U239 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U240 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U241 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U242 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U243 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U244 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U245 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U246 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U247 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U248 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U249 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U250 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U251 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U252 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U253 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U254 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U255 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U256 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U257 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U258 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U259 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U260 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U261 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U262 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U263 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U264 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U265 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U266 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U267 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U268 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U269 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U270 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U271 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U272 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U273 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U274 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U275 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U276 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U277 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U278 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U279 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U280 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U281 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U282 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U283 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U284 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U285 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U286 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U287 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U288 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U289 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U290 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U291 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U292 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U293 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U294 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U295 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U296 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U297 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U298 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U299 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U300 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U301 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U302 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U303 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U304 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U305 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U306 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U307 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U308 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U309 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U310 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U311 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U312 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U313 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U314 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U315 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U316 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U317 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U318 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U319 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U320 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U321 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U322 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U323 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U324 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U325 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U326 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U327 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U328 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U329 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U330 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U331 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U332 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U333 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U334 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U335 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U336 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U337 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U338 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U339 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U340 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U341 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U342 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U343 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U344 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U345 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U346 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U347 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U348 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U349 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U350 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U351 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U352 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U353 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U354 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND2_X1 U355 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U356 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U357 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U358 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND4_X1 U359 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_3 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X1 U1 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND4_X2 U2 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  BUF_X1 U3 ( .A(n434), .Z(n164) );
  BUF_X1 U4 ( .A(n432), .Z(n152) );
  BUF_X1 U5 ( .A(n431), .Z(n146) );
  BUF_X1 U6 ( .A(n139), .Z(n140) );
  BUF_X1 U7 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U8 ( .A(n434), .Z(n165) );
  CLKBUF_X1 U9 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U10 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U11 ( .A(n139), .Z(n141) );
  CLKBUF_X1 U12 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U13 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U14 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U15 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U16 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U17 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U18 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U19 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U20 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U21 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U22 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U23 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U24 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U25 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U26 ( .A(n433), .Z(n162) );
  CLKBUF_X1 U27 ( .A(n433), .Z(n161) );
  AND4_X1 U28 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U29 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U30 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U31 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U32 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U33 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U34 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U35 ( .A(n434), .Z(n169) );
  INV_X1 U36 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U37 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U38 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U39 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U40 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U41 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U42 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U43 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U44 ( .A(n175), .ZN(n431) );
  NAND2_X1 U45 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U46 ( .A(n176), .ZN(n432) );
  NAND2_X1 U47 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U48 ( .A(n177), .ZN(n434) );
  INV_X1 U49 ( .A(n178), .ZN(n433) );
  AOI22_X1 U50 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U51 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U52 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U53 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U54 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U55 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U56 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U57 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U58 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U59 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U60 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U61 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U62 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U63 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U64 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U65 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U66 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U67 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U68 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U69 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U70 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U71 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U72 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U73 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U74 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U75 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U76 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U77 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U78 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U79 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U80 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U81 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U82 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U83 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U84 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U85 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND4_X1 U86 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  NAND2_X1 U87 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U88 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U89 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U90 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U91 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U92 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U93 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U94 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U95 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U96 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U97 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U98 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U99 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U100 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U101 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U102 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U103 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U104 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U105 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND4_X1 U106 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND2_X1 U107 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U108 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U109 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U110 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U111 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U112 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U113 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U114 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U115 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U116 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U117 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U118 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U119 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U120 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U121 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U122 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U123 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U124 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U125 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U126 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U127 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U128 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U129 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U130 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U131 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U132 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U133 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U134 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U135 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U136 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U137 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U138 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U139 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U140 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U141 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U142 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U143 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U144 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U145 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U146 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U147 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U148 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U149 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U150 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U151 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U152 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U153 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U154 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U155 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U156 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U157 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U158 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U159 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U160 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U161 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U162 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U163 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U164 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U165 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U166 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U167 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U168 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U169 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U170 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U171 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U172 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U173 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U174 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U175 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U176 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U177 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U178 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U179 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U180 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U181 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U182 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U183 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U184 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U185 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U186 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U187 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U188 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U189 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U190 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U191 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U192 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U193 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U194 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U195 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U196 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U197 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U198 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U199 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U200 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U201 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U202 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U203 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U204 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U205 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U206 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U207 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U208 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U209 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U210 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U211 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U212 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U213 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U214 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U215 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U216 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U217 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U218 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U219 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U220 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U221 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U222 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U223 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U224 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U225 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U226 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U227 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U228 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U229 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U230 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U231 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U232 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U233 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U234 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U235 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U236 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U237 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U238 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U239 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U240 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U241 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U242 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U243 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U244 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U245 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U246 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U247 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U248 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U249 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U250 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U251 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U252 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U253 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U254 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U255 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U256 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U257 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U258 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U259 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U260 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U261 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U262 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U263 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U264 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U265 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U266 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U267 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U268 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U269 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U270 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U271 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U272 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U273 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U274 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U275 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U276 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U277 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U278 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U279 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U280 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U281 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U282 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U283 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U284 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U285 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U286 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U287 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U288 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U289 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U290 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U291 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U292 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U293 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U294 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U295 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U296 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U297 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U298 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U299 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U300 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U301 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U302 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U303 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U304 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U305 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U306 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U307 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U308 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U309 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U310 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U311 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U312 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U313 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U314 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U315 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U316 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U317 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U318 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U319 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U320 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U321 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U322 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U323 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U324 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U325 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U326 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U327 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U328 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U329 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U330 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U331 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U332 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U333 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U334 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U335 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U336 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U337 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U338 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U339 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U340 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U341 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U342 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U343 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U344 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U345 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U346 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U347 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U348 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U349 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U350 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND2_X1 U351 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U352 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U353 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U354 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND2_X1 U355 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U356 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U357 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U358 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND4_X1 U359 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_2 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  NAND4_X2 U1 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  CLKBUF_X1 U2 ( .A(n434), .Z(n165) );
  CLKBUF_X1 U3 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U4 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U5 ( .A(n433), .Z(n159) );
  BUF_X1 U6 ( .A(n139), .Z(n140) );
  BUF_X1 U7 ( .A(n434), .Z(n164) );
  BUF_X1 U8 ( .A(n432), .Z(n152) );
  BUF_X1 U9 ( .A(n431), .Z(n146) );
  CLKBUF_X1 U10 ( .A(n139), .Z(n141) );
  BUF_X1 U11 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U12 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U13 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U14 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U15 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U16 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U17 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U18 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U19 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U20 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U21 ( .A(n433), .Z(n161) );
  CLKBUF_X1 U22 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U23 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U24 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U25 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U26 ( .A(n433), .Z(n162) );
  AND4_X1 U27 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U28 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U29 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U30 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U31 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U32 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U33 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U34 ( .A(n434), .Z(n169) );
  INV_X1 U35 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U36 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U37 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U38 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U39 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U40 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U41 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U42 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U43 ( .A(n175), .ZN(n431) );
  NAND2_X1 U44 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U45 ( .A(n176), .ZN(n432) );
  NAND2_X1 U46 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U47 ( .A(n177), .ZN(n434) );
  INV_X1 U48 ( .A(n178), .ZN(n433) );
  AOI22_X1 U49 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U50 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U51 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U52 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U53 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U54 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U55 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U56 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U57 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U58 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U59 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U60 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U61 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U62 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U63 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U64 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U65 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U66 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U67 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U68 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U69 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U70 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U71 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U72 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U73 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U74 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U75 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U76 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U77 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U78 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U79 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U80 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U81 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U82 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U83 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U84 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND4_X1 U85 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  NAND2_X1 U86 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U87 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U88 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U89 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U90 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U91 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U92 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U93 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U94 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U95 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U96 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U97 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U98 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U99 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U100 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U101 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U102 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U103 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U104 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND4_X1 U105 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND2_X1 U106 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U107 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U108 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U109 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U110 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U111 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U112 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U113 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U114 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U115 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U116 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U117 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U118 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U119 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U120 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U121 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U122 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U123 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U124 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U125 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U126 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U127 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U128 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U129 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U130 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U131 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U132 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U133 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U134 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U135 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U136 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U137 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U138 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U139 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U140 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U141 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U142 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U143 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U144 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U145 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U146 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U147 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U148 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U149 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U150 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U151 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U152 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U153 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U154 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U155 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U156 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U157 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U158 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U159 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U160 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U161 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U162 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U163 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U164 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U165 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U166 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U167 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U168 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U169 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U170 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U171 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U172 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U173 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U174 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U175 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U176 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U177 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U178 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U179 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U180 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U181 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U182 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U183 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U184 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U185 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U186 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U187 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U188 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U189 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U190 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U191 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U192 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U193 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U194 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U195 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U196 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U197 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U198 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U199 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U200 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U201 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U202 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U203 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U204 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U205 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U206 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U207 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U208 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U209 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U210 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U211 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U212 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U213 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U214 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U215 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U216 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U217 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U218 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U219 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U220 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U221 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U222 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U223 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U224 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U225 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U226 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U227 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U228 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U229 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U230 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U231 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U232 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U233 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U234 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U235 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U236 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U237 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U238 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U239 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U240 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U241 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U242 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U243 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U244 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U245 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U246 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U247 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U248 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U249 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U250 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U251 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U252 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U253 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U254 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U255 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U256 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U257 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U258 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U259 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U260 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U261 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U262 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U263 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U264 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U265 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U266 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U267 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U268 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U269 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U270 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U271 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U272 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U273 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U274 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U275 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U276 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U277 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U278 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U279 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U280 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U281 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U282 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U283 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U284 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U285 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U286 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U287 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U288 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U289 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U290 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U291 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U292 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U293 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U294 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U295 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U296 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U297 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U298 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U299 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U300 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U301 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U302 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U303 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U304 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U305 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U306 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U307 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U308 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U309 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U310 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U311 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U312 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U313 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U314 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U315 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U316 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U317 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U318 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U319 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U320 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U321 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U322 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U323 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U324 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U325 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U326 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U327 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U328 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U329 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U330 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U331 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U332 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U333 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U334 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U335 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U336 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U337 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U338 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U339 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U340 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U341 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U342 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U343 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U344 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U345 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U346 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U347 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U348 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U349 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U350 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U351 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U352 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U353 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U354 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND2_X1 U355 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U356 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U357 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U358 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND4_X1 U359 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module MUX51_GENERIC_N64_1 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438;

  BUF_X1 U1 ( .A(n434), .Z(n164) );
  BUF_X1 U2 ( .A(n432), .Z(n152) );
  BUF_X1 U3 ( .A(n431), .Z(n146) );
  BUF_X1 U4 ( .A(n139), .Z(n140) );
  CLKBUF_X1 U5 ( .A(n139), .Z(n141) );
  BUF_X1 U6 ( .A(n433), .Z(n158) );
  CLKBUF_X1 U7 ( .A(n434), .Z(n165) );
  CLKBUF_X1 U8 ( .A(n434), .Z(n166) );
  CLKBUF_X1 U9 ( .A(n432), .Z(n153) );
  CLKBUF_X1 U10 ( .A(n432), .Z(n154) );
  CLKBUF_X1 U11 ( .A(n431), .Z(n147) );
  CLKBUF_X1 U12 ( .A(n431), .Z(n148) );
  CLKBUF_X1 U13 ( .A(n139), .Z(n142) );
  CLKBUF_X1 U14 ( .A(n433), .Z(n159) );
  CLKBUF_X1 U15 ( .A(n433), .Z(n160) );
  CLKBUF_X1 U16 ( .A(n434), .Z(n167) );
  CLKBUF_X1 U17 ( .A(n432), .Z(n155) );
  CLKBUF_X1 U18 ( .A(n431), .Z(n149) );
  CLKBUF_X1 U19 ( .A(n139), .Z(n143) );
  CLKBUF_X1 U20 ( .A(n433), .Z(n161) );
  CLKBUF_X1 U21 ( .A(n434), .Z(n168) );
  CLKBUF_X1 U22 ( .A(n432), .Z(n156) );
  CLKBUF_X1 U23 ( .A(n431), .Z(n150) );
  CLKBUF_X1 U24 ( .A(n139), .Z(n144) );
  CLKBUF_X1 U25 ( .A(n433), .Z(n162) );
  AND4_X1 U26 ( .A1(n175), .A2(n176), .A3(n178), .A4(n177), .ZN(n139) );
  NAND2_X1 U27 ( .A1(n174), .A2(n173), .ZN(n177) );
  NAND2_X1 U28 ( .A1(n174), .A2(n171), .ZN(n178) );
  CLKBUF_X1 U29 ( .A(n139), .Z(n145) );
  CLKBUF_X1 U30 ( .A(n431), .Z(n151) );
  CLKBUF_X1 U31 ( .A(n432), .Z(n157) );
  CLKBUF_X1 U32 ( .A(n433), .Z(n163) );
  CLKBUF_X1 U33 ( .A(n434), .Z(n169) );
  INV_X1 U34 ( .A(SEL[1]), .ZN(n172) );
  INV_X1 U35 ( .A(SEL[2]), .ZN(n170) );
  NAND3_X1 U36 ( .A1(SEL[0]), .A2(n172), .A3(n170), .ZN(n175) );
  NAND3_X1 U37 ( .A1(SEL[0]), .A2(SEL[1]), .A3(n170), .ZN(n176) );
  INV_X1 U38 ( .A(SEL[0]), .ZN(n174) );
  NOR2_X1 U39 ( .A1(SEL[1]), .A2(SEL[2]), .ZN(n171) );
  NOR2_X1 U40 ( .A1(n172), .A2(SEL[2]), .ZN(n173) );
  NAND2_X1 U41 ( .A1(E[0]), .A2(n140), .ZN(n182) );
  INV_X1 U42 ( .A(n175), .ZN(n431) );
  NAND2_X1 U43 ( .A1(B[0]), .A2(n146), .ZN(n181) );
  INV_X1 U44 ( .A(n176), .ZN(n432) );
  NAND2_X1 U45 ( .A1(D[0]), .A2(n152), .ZN(n180) );
  INV_X1 U46 ( .A(n177), .ZN(n434) );
  INV_X1 U47 ( .A(n178), .ZN(n433) );
  AOI22_X1 U48 ( .A1(C[0]), .A2(n164), .B1(A[0]), .B2(n158), .ZN(n179) );
  NAND4_X1 U49 ( .A1(n182), .A2(n181), .A3(n180), .A4(n179), .ZN(Y[0]) );
  NAND2_X1 U50 ( .A1(E[1]), .A2(n140), .ZN(n186) );
  NAND2_X1 U51 ( .A1(B[1]), .A2(n146), .ZN(n185) );
  NAND2_X1 U52 ( .A1(D[1]), .A2(n152), .ZN(n184) );
  AOI22_X1 U53 ( .A1(C[1]), .A2(n164), .B1(A[1]), .B2(n158), .ZN(n183) );
  NAND4_X1 U54 ( .A1(n186), .A2(n185), .A3(n184), .A4(n183), .ZN(Y[1]) );
  NAND2_X1 U55 ( .A1(E[2]), .A2(n140), .ZN(n190) );
  NAND2_X1 U56 ( .A1(B[2]), .A2(n146), .ZN(n189) );
  NAND2_X1 U57 ( .A1(D[2]), .A2(n152), .ZN(n188) );
  AOI22_X1 U58 ( .A1(C[2]), .A2(n164), .B1(A[2]), .B2(n158), .ZN(n187) );
  NAND4_X1 U59 ( .A1(n190), .A2(n189), .A3(n188), .A4(n187), .ZN(Y[2]) );
  NAND2_X1 U60 ( .A1(E[3]), .A2(n140), .ZN(n194) );
  NAND2_X1 U61 ( .A1(B[3]), .A2(n146), .ZN(n193) );
  NAND2_X1 U62 ( .A1(D[3]), .A2(n152), .ZN(n192) );
  AOI22_X1 U63 ( .A1(C[3]), .A2(n164), .B1(A[3]), .B2(n158), .ZN(n191) );
  NAND4_X1 U64 ( .A1(n194), .A2(n193), .A3(n192), .A4(n191), .ZN(Y[3]) );
  NAND2_X1 U65 ( .A1(E[4]), .A2(n140), .ZN(n198) );
  NAND2_X1 U66 ( .A1(B[4]), .A2(n146), .ZN(n197) );
  NAND2_X1 U67 ( .A1(D[4]), .A2(n152), .ZN(n196) );
  AOI22_X1 U68 ( .A1(C[4]), .A2(n164), .B1(A[4]), .B2(n158), .ZN(n195) );
  NAND4_X1 U69 ( .A1(n198), .A2(n197), .A3(n196), .A4(n195), .ZN(Y[4]) );
  NAND2_X1 U70 ( .A1(E[5]), .A2(n140), .ZN(n202) );
  NAND2_X1 U71 ( .A1(B[5]), .A2(n146), .ZN(n201) );
  NAND2_X1 U72 ( .A1(D[5]), .A2(n152), .ZN(n200) );
  AOI22_X1 U73 ( .A1(C[5]), .A2(n164), .B1(A[5]), .B2(n158), .ZN(n199) );
  NAND4_X1 U74 ( .A1(n202), .A2(n201), .A3(n200), .A4(n199), .ZN(Y[5]) );
  NAND2_X1 U75 ( .A1(E[6]), .A2(n140), .ZN(n206) );
  NAND2_X1 U76 ( .A1(B[6]), .A2(n146), .ZN(n205) );
  NAND2_X1 U77 ( .A1(D[6]), .A2(n152), .ZN(n204) );
  AOI22_X1 U78 ( .A1(C[6]), .A2(n164), .B1(A[6]), .B2(n158), .ZN(n203) );
  NAND4_X1 U79 ( .A1(n206), .A2(n205), .A3(n204), .A4(n203), .ZN(Y[6]) );
  NAND2_X1 U80 ( .A1(E[7]), .A2(n140), .ZN(n210) );
  NAND2_X1 U81 ( .A1(B[7]), .A2(n146), .ZN(n209) );
  NAND2_X1 U82 ( .A1(D[7]), .A2(n152), .ZN(n208) );
  AOI22_X1 U83 ( .A1(C[7]), .A2(n164), .B1(A[7]), .B2(n158), .ZN(n207) );
  NAND4_X1 U84 ( .A1(n210), .A2(n209), .A3(n208), .A4(n207), .ZN(Y[7]) );
  NAND2_X1 U85 ( .A1(E[8]), .A2(n140), .ZN(n214) );
  NAND2_X1 U86 ( .A1(B[8]), .A2(n146), .ZN(n213) );
  NAND2_X1 U87 ( .A1(D[8]), .A2(n152), .ZN(n212) );
  AOI22_X1 U88 ( .A1(C[8]), .A2(n164), .B1(A[8]), .B2(n158), .ZN(n211) );
  NAND4_X1 U89 ( .A1(n214), .A2(n213), .A3(n212), .A4(n211), .ZN(Y[8]) );
  NAND2_X1 U90 ( .A1(E[9]), .A2(n140), .ZN(n218) );
  NAND2_X1 U91 ( .A1(B[9]), .A2(n146), .ZN(n217) );
  NAND2_X1 U92 ( .A1(D[9]), .A2(n152), .ZN(n216) );
  AOI22_X1 U93 ( .A1(C[9]), .A2(n164), .B1(A[9]), .B2(n158), .ZN(n215) );
  NAND4_X1 U94 ( .A1(n218), .A2(n217), .A3(n216), .A4(n215), .ZN(Y[9]) );
  NAND2_X1 U95 ( .A1(E[10]), .A2(n140), .ZN(n222) );
  NAND2_X1 U96 ( .A1(B[10]), .A2(n146), .ZN(n221) );
  NAND2_X1 U97 ( .A1(D[10]), .A2(n152), .ZN(n220) );
  AOI22_X1 U98 ( .A1(C[10]), .A2(n164), .B1(A[10]), .B2(n158), .ZN(n219) );
  NAND4_X1 U99 ( .A1(n222), .A2(n221), .A3(n220), .A4(n219), .ZN(Y[10]) );
  NAND2_X1 U100 ( .A1(E[11]), .A2(n140), .ZN(n226) );
  NAND2_X1 U101 ( .A1(B[11]), .A2(n146), .ZN(n225) );
  NAND2_X1 U102 ( .A1(D[11]), .A2(n152), .ZN(n224) );
  AOI22_X1 U103 ( .A1(C[11]), .A2(n164), .B1(A[11]), .B2(n158), .ZN(n223) );
  NAND4_X1 U104 ( .A1(n226), .A2(n225), .A3(n224), .A4(n223), .ZN(Y[11]) );
  NAND2_X1 U105 ( .A1(E[12]), .A2(n141), .ZN(n230) );
  NAND2_X1 U106 ( .A1(B[12]), .A2(n147), .ZN(n229) );
  NAND2_X1 U107 ( .A1(D[12]), .A2(n153), .ZN(n228) );
  AOI22_X1 U108 ( .A1(C[12]), .A2(n165), .B1(A[12]), .B2(n159), .ZN(n227) );
  NAND4_X1 U109 ( .A1(n230), .A2(n229), .A3(n228), .A4(n227), .ZN(Y[12]) );
  NAND2_X1 U110 ( .A1(E[13]), .A2(n141), .ZN(n234) );
  NAND2_X1 U111 ( .A1(B[13]), .A2(n147), .ZN(n233) );
  NAND2_X1 U112 ( .A1(D[13]), .A2(n153), .ZN(n232) );
  AOI22_X1 U113 ( .A1(C[13]), .A2(n165), .B1(A[13]), .B2(n159), .ZN(n231) );
  NAND4_X1 U114 ( .A1(n234), .A2(n233), .A3(n232), .A4(n231), .ZN(Y[13]) );
  NAND2_X1 U115 ( .A1(E[14]), .A2(n141), .ZN(n238) );
  NAND2_X1 U116 ( .A1(B[14]), .A2(n147), .ZN(n237) );
  NAND2_X1 U117 ( .A1(D[14]), .A2(n153), .ZN(n236) );
  AOI22_X1 U118 ( .A1(C[14]), .A2(n165), .B1(A[14]), .B2(n159), .ZN(n235) );
  NAND4_X1 U119 ( .A1(n238), .A2(n237), .A3(n236), .A4(n235), .ZN(Y[14]) );
  NAND2_X1 U120 ( .A1(E[15]), .A2(n141), .ZN(n242) );
  NAND2_X1 U121 ( .A1(B[15]), .A2(n147), .ZN(n241) );
  NAND2_X1 U122 ( .A1(D[15]), .A2(n153), .ZN(n240) );
  AOI22_X1 U123 ( .A1(C[15]), .A2(n165), .B1(A[15]), .B2(n159), .ZN(n239) );
  NAND4_X1 U124 ( .A1(n242), .A2(n241), .A3(n240), .A4(n239), .ZN(Y[15]) );
  NAND2_X1 U125 ( .A1(E[16]), .A2(n141), .ZN(n246) );
  NAND2_X1 U126 ( .A1(B[16]), .A2(n147), .ZN(n245) );
  NAND2_X1 U127 ( .A1(D[16]), .A2(n153), .ZN(n244) );
  AOI22_X1 U128 ( .A1(C[16]), .A2(n165), .B1(A[16]), .B2(n159), .ZN(n243) );
  NAND4_X1 U129 ( .A1(n246), .A2(n245), .A3(n244), .A4(n243), .ZN(Y[16]) );
  NAND2_X1 U130 ( .A1(E[17]), .A2(n141), .ZN(n250) );
  NAND2_X1 U131 ( .A1(B[17]), .A2(n147), .ZN(n249) );
  NAND2_X1 U132 ( .A1(D[17]), .A2(n153), .ZN(n248) );
  AOI22_X1 U133 ( .A1(C[17]), .A2(n165), .B1(A[17]), .B2(n159), .ZN(n247) );
  NAND4_X1 U134 ( .A1(n250), .A2(n249), .A3(n248), .A4(n247), .ZN(Y[17]) );
  NAND2_X1 U135 ( .A1(E[18]), .A2(n141), .ZN(n254) );
  NAND2_X1 U136 ( .A1(B[18]), .A2(n147), .ZN(n253) );
  NAND2_X1 U137 ( .A1(D[18]), .A2(n153), .ZN(n252) );
  AOI22_X1 U138 ( .A1(C[18]), .A2(n165), .B1(A[18]), .B2(n159), .ZN(n251) );
  NAND4_X1 U139 ( .A1(n254), .A2(n253), .A3(n252), .A4(n251), .ZN(Y[18]) );
  NAND2_X1 U140 ( .A1(E[19]), .A2(n141), .ZN(n258) );
  NAND2_X1 U141 ( .A1(B[19]), .A2(n147), .ZN(n257) );
  NAND2_X1 U142 ( .A1(D[19]), .A2(n153), .ZN(n256) );
  AOI22_X1 U143 ( .A1(C[19]), .A2(n165), .B1(A[19]), .B2(n159), .ZN(n255) );
  NAND4_X1 U144 ( .A1(n258), .A2(n257), .A3(n256), .A4(n255), .ZN(Y[19]) );
  NAND2_X1 U145 ( .A1(E[20]), .A2(n141), .ZN(n262) );
  NAND2_X1 U146 ( .A1(B[20]), .A2(n147), .ZN(n261) );
  NAND2_X1 U147 ( .A1(D[20]), .A2(n153), .ZN(n260) );
  AOI22_X1 U148 ( .A1(C[20]), .A2(n165), .B1(A[20]), .B2(n159), .ZN(n259) );
  NAND4_X1 U149 ( .A1(n262), .A2(n261), .A3(n260), .A4(n259), .ZN(Y[20]) );
  NAND2_X1 U150 ( .A1(E[21]), .A2(n141), .ZN(n266) );
  NAND2_X1 U151 ( .A1(B[21]), .A2(n147), .ZN(n265) );
  NAND2_X1 U152 ( .A1(D[21]), .A2(n153), .ZN(n264) );
  AOI22_X1 U153 ( .A1(C[21]), .A2(n165), .B1(A[21]), .B2(n159), .ZN(n263) );
  NAND4_X1 U154 ( .A1(n266), .A2(n265), .A3(n264), .A4(n263), .ZN(Y[21]) );
  NAND2_X1 U155 ( .A1(E[22]), .A2(n141), .ZN(n270) );
  NAND2_X1 U156 ( .A1(B[22]), .A2(n147), .ZN(n269) );
  NAND2_X1 U157 ( .A1(D[22]), .A2(n153), .ZN(n268) );
  AOI22_X1 U158 ( .A1(C[22]), .A2(n165), .B1(A[22]), .B2(n159), .ZN(n267) );
  NAND4_X1 U159 ( .A1(n270), .A2(n269), .A3(n268), .A4(n267), .ZN(Y[22]) );
  NAND2_X1 U160 ( .A1(E[23]), .A2(n141), .ZN(n274) );
  NAND2_X1 U161 ( .A1(B[23]), .A2(n147), .ZN(n273) );
  NAND2_X1 U162 ( .A1(D[23]), .A2(n153), .ZN(n272) );
  AOI22_X1 U163 ( .A1(C[23]), .A2(n165), .B1(A[23]), .B2(n159), .ZN(n271) );
  NAND4_X1 U164 ( .A1(n274), .A2(n273), .A3(n272), .A4(n271), .ZN(Y[23]) );
  NAND2_X1 U165 ( .A1(E[24]), .A2(n142), .ZN(n278) );
  NAND2_X1 U166 ( .A1(B[24]), .A2(n148), .ZN(n277) );
  NAND2_X1 U167 ( .A1(D[24]), .A2(n154), .ZN(n276) );
  AOI22_X1 U168 ( .A1(C[24]), .A2(n166), .B1(A[24]), .B2(n160), .ZN(n275) );
  NAND4_X1 U169 ( .A1(n278), .A2(n277), .A3(n276), .A4(n275), .ZN(Y[24]) );
  NAND2_X1 U170 ( .A1(E[25]), .A2(n142), .ZN(n282) );
  NAND2_X1 U171 ( .A1(B[25]), .A2(n148), .ZN(n281) );
  NAND2_X1 U172 ( .A1(D[25]), .A2(n154), .ZN(n280) );
  AOI22_X1 U173 ( .A1(C[25]), .A2(n166), .B1(A[25]), .B2(n160), .ZN(n279) );
  NAND4_X1 U174 ( .A1(n282), .A2(n281), .A3(n280), .A4(n279), .ZN(Y[25]) );
  NAND2_X1 U175 ( .A1(E[26]), .A2(n142), .ZN(n286) );
  NAND2_X1 U176 ( .A1(B[26]), .A2(n148), .ZN(n285) );
  NAND2_X1 U177 ( .A1(D[26]), .A2(n154), .ZN(n284) );
  AOI22_X1 U178 ( .A1(C[26]), .A2(n166), .B1(A[26]), .B2(n160), .ZN(n283) );
  NAND4_X1 U179 ( .A1(n286), .A2(n285), .A3(n284), .A4(n283), .ZN(Y[26]) );
  NAND2_X1 U180 ( .A1(E[27]), .A2(n142), .ZN(n290) );
  NAND2_X1 U181 ( .A1(B[27]), .A2(n148), .ZN(n289) );
  NAND2_X1 U182 ( .A1(D[27]), .A2(n154), .ZN(n288) );
  AOI22_X1 U183 ( .A1(C[27]), .A2(n166), .B1(A[27]), .B2(n160), .ZN(n287) );
  NAND4_X1 U184 ( .A1(n290), .A2(n289), .A3(n288), .A4(n287), .ZN(Y[27]) );
  NAND2_X1 U185 ( .A1(E[28]), .A2(n142), .ZN(n294) );
  NAND2_X1 U186 ( .A1(B[28]), .A2(n148), .ZN(n293) );
  NAND2_X1 U187 ( .A1(D[28]), .A2(n154), .ZN(n292) );
  AOI22_X1 U188 ( .A1(C[28]), .A2(n166), .B1(A[28]), .B2(n160), .ZN(n291) );
  NAND4_X1 U189 ( .A1(n294), .A2(n293), .A3(n292), .A4(n291), .ZN(Y[28]) );
  NAND2_X1 U190 ( .A1(E[29]), .A2(n142), .ZN(n298) );
  NAND2_X1 U191 ( .A1(B[29]), .A2(n148), .ZN(n297) );
  NAND2_X1 U192 ( .A1(D[29]), .A2(n154), .ZN(n296) );
  AOI22_X1 U193 ( .A1(C[29]), .A2(n166), .B1(A[29]), .B2(n160), .ZN(n295) );
  NAND4_X1 U194 ( .A1(n298), .A2(n297), .A3(n296), .A4(n295), .ZN(Y[29]) );
  NAND2_X1 U195 ( .A1(E[30]), .A2(n142), .ZN(n302) );
  NAND2_X1 U196 ( .A1(B[30]), .A2(n148), .ZN(n301) );
  NAND2_X1 U197 ( .A1(D[30]), .A2(n154), .ZN(n300) );
  AOI22_X1 U198 ( .A1(C[30]), .A2(n166), .B1(A[30]), .B2(n160), .ZN(n299) );
  NAND4_X1 U199 ( .A1(n302), .A2(n301), .A3(n300), .A4(n299), .ZN(Y[30]) );
  NAND2_X1 U200 ( .A1(E[31]), .A2(n142), .ZN(n306) );
  NAND2_X1 U201 ( .A1(B[31]), .A2(n148), .ZN(n305) );
  NAND2_X1 U202 ( .A1(D[31]), .A2(n154), .ZN(n304) );
  AOI22_X1 U203 ( .A1(C[31]), .A2(n166), .B1(A[31]), .B2(n160), .ZN(n303) );
  NAND4_X1 U204 ( .A1(n306), .A2(n305), .A3(n304), .A4(n303), .ZN(Y[31]) );
  NAND2_X1 U205 ( .A1(E[32]), .A2(n142), .ZN(n310) );
  NAND2_X1 U206 ( .A1(B[32]), .A2(n148), .ZN(n309) );
  NAND2_X1 U207 ( .A1(D[32]), .A2(n154), .ZN(n308) );
  AOI22_X1 U208 ( .A1(C[32]), .A2(n166), .B1(A[32]), .B2(n160), .ZN(n307) );
  NAND4_X1 U209 ( .A1(n310), .A2(n309), .A3(n308), .A4(n307), .ZN(Y[32]) );
  NAND2_X1 U210 ( .A1(E[33]), .A2(n142), .ZN(n314) );
  NAND2_X1 U211 ( .A1(B[33]), .A2(n148), .ZN(n313) );
  NAND2_X1 U212 ( .A1(D[33]), .A2(n154), .ZN(n312) );
  AOI22_X1 U213 ( .A1(C[33]), .A2(n166), .B1(A[33]), .B2(n160), .ZN(n311) );
  NAND4_X1 U214 ( .A1(n314), .A2(n313), .A3(n312), .A4(n311), .ZN(Y[33]) );
  NAND2_X1 U215 ( .A1(E[34]), .A2(n142), .ZN(n318) );
  NAND2_X1 U216 ( .A1(B[34]), .A2(n148), .ZN(n317) );
  NAND2_X1 U217 ( .A1(D[34]), .A2(n154), .ZN(n316) );
  AOI22_X1 U218 ( .A1(C[34]), .A2(n166), .B1(A[34]), .B2(n160), .ZN(n315) );
  NAND4_X1 U219 ( .A1(n318), .A2(n317), .A3(n316), .A4(n315), .ZN(Y[34]) );
  NAND2_X1 U220 ( .A1(E[35]), .A2(n142), .ZN(n322) );
  NAND2_X1 U221 ( .A1(B[35]), .A2(n148), .ZN(n321) );
  NAND2_X1 U222 ( .A1(D[35]), .A2(n154), .ZN(n320) );
  AOI22_X1 U223 ( .A1(C[35]), .A2(n166), .B1(A[35]), .B2(n160), .ZN(n319) );
  NAND4_X1 U224 ( .A1(n322), .A2(n321), .A3(n320), .A4(n319), .ZN(Y[35]) );
  NAND2_X1 U225 ( .A1(E[36]), .A2(n143), .ZN(n326) );
  NAND2_X1 U226 ( .A1(B[36]), .A2(n149), .ZN(n325) );
  NAND2_X1 U227 ( .A1(D[36]), .A2(n155), .ZN(n324) );
  AOI22_X1 U228 ( .A1(C[36]), .A2(n167), .B1(A[36]), .B2(n161), .ZN(n323) );
  NAND4_X1 U229 ( .A1(n326), .A2(n325), .A3(n324), .A4(n323), .ZN(Y[36]) );
  NAND2_X1 U230 ( .A1(E[37]), .A2(n143), .ZN(n330) );
  NAND2_X1 U231 ( .A1(B[37]), .A2(n149), .ZN(n329) );
  NAND2_X1 U232 ( .A1(D[37]), .A2(n155), .ZN(n328) );
  AOI22_X1 U233 ( .A1(C[37]), .A2(n167), .B1(A[37]), .B2(n161), .ZN(n327) );
  NAND4_X1 U234 ( .A1(n330), .A2(n329), .A3(n328), .A4(n327), .ZN(Y[37]) );
  NAND2_X1 U235 ( .A1(E[38]), .A2(n143), .ZN(n334) );
  NAND2_X1 U236 ( .A1(B[38]), .A2(n149), .ZN(n333) );
  NAND2_X1 U237 ( .A1(D[38]), .A2(n155), .ZN(n332) );
  AOI22_X1 U238 ( .A1(C[38]), .A2(n167), .B1(A[38]), .B2(n161), .ZN(n331) );
  NAND4_X1 U239 ( .A1(n334), .A2(n333), .A3(n332), .A4(n331), .ZN(Y[38]) );
  NAND2_X1 U240 ( .A1(E[39]), .A2(n143), .ZN(n338) );
  NAND2_X1 U241 ( .A1(B[39]), .A2(n149), .ZN(n337) );
  NAND2_X1 U242 ( .A1(D[39]), .A2(n155), .ZN(n336) );
  AOI22_X1 U243 ( .A1(C[39]), .A2(n167), .B1(A[39]), .B2(n161), .ZN(n335) );
  NAND4_X1 U244 ( .A1(n338), .A2(n337), .A3(n336), .A4(n335), .ZN(Y[39]) );
  NAND2_X1 U245 ( .A1(E[40]), .A2(n143), .ZN(n342) );
  NAND2_X1 U246 ( .A1(B[40]), .A2(n149), .ZN(n341) );
  NAND2_X1 U247 ( .A1(D[40]), .A2(n155), .ZN(n340) );
  AOI22_X1 U248 ( .A1(C[40]), .A2(n167), .B1(A[40]), .B2(n161), .ZN(n339) );
  NAND4_X1 U249 ( .A1(n342), .A2(n341), .A3(n340), .A4(n339), .ZN(Y[40]) );
  NAND2_X1 U250 ( .A1(E[41]), .A2(n143), .ZN(n346) );
  NAND2_X1 U251 ( .A1(B[41]), .A2(n149), .ZN(n345) );
  NAND2_X1 U252 ( .A1(D[41]), .A2(n155), .ZN(n344) );
  AOI22_X1 U253 ( .A1(C[41]), .A2(n167), .B1(A[41]), .B2(n161), .ZN(n343) );
  NAND4_X1 U254 ( .A1(n346), .A2(n345), .A3(n344), .A4(n343), .ZN(Y[41]) );
  NAND2_X1 U255 ( .A1(E[42]), .A2(n143), .ZN(n350) );
  NAND2_X1 U256 ( .A1(B[42]), .A2(n149), .ZN(n349) );
  NAND2_X1 U257 ( .A1(D[42]), .A2(n155), .ZN(n348) );
  AOI22_X1 U258 ( .A1(C[42]), .A2(n167), .B1(A[42]), .B2(n161), .ZN(n347) );
  NAND4_X1 U259 ( .A1(n350), .A2(n349), .A3(n348), .A4(n347), .ZN(Y[42]) );
  NAND2_X1 U260 ( .A1(E[43]), .A2(n143), .ZN(n354) );
  NAND2_X1 U261 ( .A1(B[43]), .A2(n149), .ZN(n353) );
  NAND2_X1 U262 ( .A1(D[43]), .A2(n155), .ZN(n352) );
  AOI22_X1 U263 ( .A1(C[43]), .A2(n167), .B1(A[43]), .B2(n161), .ZN(n351) );
  NAND4_X1 U264 ( .A1(n354), .A2(n353), .A3(n352), .A4(n351), .ZN(Y[43]) );
  NAND2_X1 U265 ( .A1(E[44]), .A2(n143), .ZN(n358) );
  NAND2_X1 U266 ( .A1(B[44]), .A2(n149), .ZN(n357) );
  NAND2_X1 U267 ( .A1(D[44]), .A2(n155), .ZN(n356) );
  AOI22_X1 U268 ( .A1(C[44]), .A2(n167), .B1(A[44]), .B2(n161), .ZN(n355) );
  NAND4_X1 U269 ( .A1(n358), .A2(n357), .A3(n356), .A4(n355), .ZN(Y[44]) );
  NAND2_X1 U270 ( .A1(E[45]), .A2(n143), .ZN(n362) );
  NAND2_X1 U271 ( .A1(B[45]), .A2(n149), .ZN(n361) );
  NAND2_X1 U272 ( .A1(D[45]), .A2(n155), .ZN(n360) );
  AOI22_X1 U273 ( .A1(C[45]), .A2(n167), .B1(A[45]), .B2(n161), .ZN(n359) );
  NAND4_X1 U274 ( .A1(n362), .A2(n361), .A3(n360), .A4(n359), .ZN(Y[45]) );
  NAND2_X1 U275 ( .A1(E[46]), .A2(n143), .ZN(n366) );
  NAND2_X1 U276 ( .A1(B[46]), .A2(n149), .ZN(n365) );
  NAND2_X1 U277 ( .A1(D[46]), .A2(n155), .ZN(n364) );
  AOI22_X1 U278 ( .A1(C[46]), .A2(n167), .B1(A[46]), .B2(n161), .ZN(n363) );
  NAND4_X1 U279 ( .A1(n366), .A2(n365), .A3(n364), .A4(n363), .ZN(Y[46]) );
  NAND2_X1 U280 ( .A1(E[47]), .A2(n143), .ZN(n370) );
  NAND2_X1 U281 ( .A1(B[47]), .A2(n149), .ZN(n369) );
  NAND2_X1 U282 ( .A1(D[47]), .A2(n155), .ZN(n368) );
  AOI22_X1 U283 ( .A1(C[47]), .A2(n167), .B1(A[47]), .B2(n161), .ZN(n367) );
  NAND4_X1 U284 ( .A1(n370), .A2(n369), .A3(n368), .A4(n367), .ZN(Y[47]) );
  NAND2_X1 U285 ( .A1(E[48]), .A2(n144), .ZN(n374) );
  NAND2_X1 U286 ( .A1(B[48]), .A2(n150), .ZN(n373) );
  NAND2_X1 U287 ( .A1(D[48]), .A2(n156), .ZN(n372) );
  AOI22_X1 U288 ( .A1(C[48]), .A2(n168), .B1(A[48]), .B2(n162), .ZN(n371) );
  NAND4_X1 U289 ( .A1(n374), .A2(n373), .A3(n372), .A4(n371), .ZN(Y[48]) );
  NAND2_X1 U290 ( .A1(E[49]), .A2(n144), .ZN(n378) );
  NAND2_X1 U291 ( .A1(B[49]), .A2(n150), .ZN(n377) );
  NAND2_X1 U292 ( .A1(D[49]), .A2(n156), .ZN(n376) );
  AOI22_X1 U293 ( .A1(C[49]), .A2(n168), .B1(A[49]), .B2(n162), .ZN(n375) );
  NAND4_X1 U294 ( .A1(n378), .A2(n377), .A3(n376), .A4(n375), .ZN(Y[49]) );
  NAND2_X1 U295 ( .A1(E[50]), .A2(n144), .ZN(n382) );
  NAND2_X1 U296 ( .A1(B[50]), .A2(n150), .ZN(n381) );
  NAND2_X1 U297 ( .A1(D[50]), .A2(n156), .ZN(n380) );
  AOI22_X1 U298 ( .A1(C[50]), .A2(n168), .B1(A[50]), .B2(n162), .ZN(n379) );
  NAND4_X1 U299 ( .A1(n382), .A2(n381), .A3(n380), .A4(n379), .ZN(Y[50]) );
  NAND2_X1 U300 ( .A1(E[51]), .A2(n144), .ZN(n386) );
  NAND2_X1 U301 ( .A1(B[51]), .A2(n150), .ZN(n385) );
  NAND2_X1 U302 ( .A1(D[51]), .A2(n156), .ZN(n384) );
  AOI22_X1 U303 ( .A1(C[51]), .A2(n168), .B1(A[51]), .B2(n162), .ZN(n383) );
  NAND4_X1 U304 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(Y[51]) );
  NAND2_X1 U305 ( .A1(E[52]), .A2(n144), .ZN(n390) );
  NAND2_X1 U306 ( .A1(B[52]), .A2(n150), .ZN(n389) );
  NAND2_X1 U307 ( .A1(D[52]), .A2(n156), .ZN(n388) );
  AOI22_X1 U308 ( .A1(C[52]), .A2(n168), .B1(A[52]), .B2(n162), .ZN(n387) );
  NAND4_X1 U309 ( .A1(n390), .A2(n389), .A3(n388), .A4(n387), .ZN(Y[52]) );
  NAND2_X1 U310 ( .A1(E[53]), .A2(n144), .ZN(n394) );
  NAND2_X1 U311 ( .A1(B[53]), .A2(n150), .ZN(n393) );
  NAND2_X1 U312 ( .A1(D[53]), .A2(n156), .ZN(n392) );
  AOI22_X1 U313 ( .A1(C[53]), .A2(n168), .B1(A[53]), .B2(n162), .ZN(n391) );
  NAND4_X1 U314 ( .A1(n394), .A2(n393), .A3(n392), .A4(n391), .ZN(Y[53]) );
  NAND2_X1 U315 ( .A1(E[54]), .A2(n144), .ZN(n398) );
  NAND2_X1 U316 ( .A1(B[54]), .A2(n150), .ZN(n397) );
  NAND2_X1 U317 ( .A1(D[54]), .A2(n156), .ZN(n396) );
  AOI22_X1 U318 ( .A1(C[54]), .A2(n168), .B1(A[54]), .B2(n162), .ZN(n395) );
  NAND4_X1 U319 ( .A1(n398), .A2(n397), .A3(n396), .A4(n395), .ZN(Y[54]) );
  NAND2_X1 U320 ( .A1(E[55]), .A2(n144), .ZN(n402) );
  NAND2_X1 U321 ( .A1(B[55]), .A2(n150), .ZN(n401) );
  NAND2_X1 U322 ( .A1(D[55]), .A2(n156), .ZN(n400) );
  AOI22_X1 U323 ( .A1(C[55]), .A2(n168), .B1(A[55]), .B2(n162), .ZN(n399) );
  NAND4_X1 U324 ( .A1(n402), .A2(n401), .A3(n400), .A4(n399), .ZN(Y[55]) );
  NAND2_X1 U325 ( .A1(E[56]), .A2(n144), .ZN(n406) );
  NAND2_X1 U326 ( .A1(B[56]), .A2(n150), .ZN(n405) );
  NAND2_X1 U327 ( .A1(D[56]), .A2(n156), .ZN(n404) );
  AOI22_X1 U328 ( .A1(C[56]), .A2(n168), .B1(A[56]), .B2(n162), .ZN(n403) );
  NAND4_X1 U329 ( .A1(n406), .A2(n405), .A3(n404), .A4(n403), .ZN(Y[56]) );
  NAND2_X1 U330 ( .A1(E[57]), .A2(n144), .ZN(n410) );
  NAND2_X1 U331 ( .A1(B[57]), .A2(n150), .ZN(n409) );
  NAND2_X1 U332 ( .A1(D[57]), .A2(n156), .ZN(n408) );
  AOI22_X1 U333 ( .A1(C[57]), .A2(n168), .B1(A[57]), .B2(n162), .ZN(n407) );
  NAND4_X1 U334 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(Y[57]) );
  NAND2_X1 U335 ( .A1(E[58]), .A2(n144), .ZN(n414) );
  NAND2_X1 U336 ( .A1(B[58]), .A2(n150), .ZN(n413) );
  NAND2_X1 U337 ( .A1(D[58]), .A2(n156), .ZN(n412) );
  AOI22_X1 U338 ( .A1(C[58]), .A2(n168), .B1(A[58]), .B2(n162), .ZN(n411) );
  NAND4_X1 U339 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(Y[58]) );
  NAND2_X1 U340 ( .A1(E[59]), .A2(n144), .ZN(n418) );
  NAND2_X1 U341 ( .A1(B[59]), .A2(n150), .ZN(n417) );
  NAND2_X1 U342 ( .A1(D[59]), .A2(n156), .ZN(n416) );
  AOI22_X1 U343 ( .A1(C[59]), .A2(n168), .B1(A[59]), .B2(n162), .ZN(n415) );
  NAND4_X1 U344 ( .A1(n418), .A2(n417), .A3(n416), .A4(n415), .ZN(Y[59]) );
  NAND2_X1 U345 ( .A1(E[60]), .A2(n145), .ZN(n422) );
  NAND2_X1 U346 ( .A1(B[60]), .A2(n151), .ZN(n421) );
  NAND2_X1 U347 ( .A1(D[60]), .A2(n157), .ZN(n420) );
  AOI22_X1 U348 ( .A1(C[60]), .A2(n169), .B1(A[60]), .B2(n163), .ZN(n419) );
  NAND4_X1 U349 ( .A1(n422), .A2(n421), .A3(n420), .A4(n419), .ZN(Y[60]) );
  NAND2_X1 U350 ( .A1(E[61]), .A2(n145), .ZN(n426) );
  NAND2_X1 U351 ( .A1(B[61]), .A2(n151), .ZN(n425) );
  NAND2_X1 U352 ( .A1(D[61]), .A2(n157), .ZN(n424) );
  AOI22_X1 U353 ( .A1(C[61]), .A2(n169), .B1(A[61]), .B2(n163), .ZN(n423) );
  NAND4_X1 U354 ( .A1(n426), .A2(n425), .A3(n424), .A4(n423), .ZN(Y[61]) );
  NAND2_X1 U355 ( .A1(E[62]), .A2(n145), .ZN(n430) );
  NAND2_X1 U356 ( .A1(B[62]), .A2(n151), .ZN(n429) );
  NAND2_X1 U357 ( .A1(D[62]), .A2(n157), .ZN(n428) );
  AOI22_X1 U358 ( .A1(C[62]), .A2(n169), .B1(A[62]), .B2(n163), .ZN(n427) );
  NAND4_X1 U359 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(Y[62]) );
  NAND2_X1 U360 ( .A1(E[63]), .A2(n145), .ZN(n438) );
  NAND2_X1 U361 ( .A1(B[63]), .A2(n151), .ZN(n437) );
  NAND2_X1 U362 ( .A1(D[63]), .A2(n157), .ZN(n436) );
  AOI22_X1 U363 ( .A1(C[63]), .A2(n169), .B1(A[63]), .B2(n163), .ZN(n435) );
  NAND4_X1 U364 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(Y[63]) );
endmodule


module BOOTH_ENCODER_19 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7, n8, n9, n10, n11, n12, n14;

  OR2_X1 U1 ( .A1(I[1]), .A2(I[0]), .ZN(n9) );
  MUX2_X2 U2 ( .A(n5), .B(n6), .S(I[2]), .Z(O[1]) );
  AND2_X1 U3 ( .A1(I[1]), .A2(I[0]), .ZN(n5) );
  AND2_X1 U4 ( .A1(n12), .A2(n14), .ZN(n6) );
  AOI21_X1 U5 ( .B1(n10), .B2(n14), .A(I[2]), .ZN(O[0]) );
  INV_X1 U6 ( .A(I[1]), .ZN(n7) );
  INV_X1 U7 ( .A(I[0]), .ZN(n8) );
  AND3_X2 U8 ( .A1(n10), .A2(I[2]), .A3(n11), .ZN(O[2]) );
  NAND2_X1 U9 ( .A1(n9), .A2(n14), .ZN(n10) );
  NAND2_X1 U10 ( .A1(I[1]), .A2(I[0]), .ZN(n11) );
  NAND2_X1 U11 ( .A1(n7), .A2(n8), .ZN(n12) );
  NAND2_X1 U12 ( .A1(I[1]), .A2(I[0]), .ZN(n14) );
endmodule


module BOOTH_ENCODER_18 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n4, n5, n6, n7, n9, n10, n11;

  BUF_X1 U1 ( .A(n11), .Z(n4) );
  NAND2_X1 U2 ( .A1(n5), .A2(n6), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n7), .A2(n11), .ZN(n10) );
  INV_X1 U4 ( .A(I[0]), .ZN(n5) );
  INV_X1 U5 ( .A(I[1]), .ZN(n6) );
  NAND2_X1 U6 ( .A1(I[1]), .A2(I[0]), .ZN(n11) );
  AND3_X1 U7 ( .A1(n4), .A2(I[2]), .A3(n10), .ZN(O[2]) );
  AOI21_X1 U8 ( .B1(n10), .B2(n4), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U9 ( .A(n4), .B(n10), .S(I[2]), .Z(n9) );
  INV_X1 U10 ( .A(n9), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_17 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_16 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_15 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_14 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_13 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_12 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_11 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_10 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_9 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_8 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_7 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_6 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module BOOTH_ENCODER_5 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   n5, n6, n7;

  OAI21_X1 U1 ( .B1(I[0]), .B2(I[1]), .A(n7), .ZN(n6) );
  NAND2_X1 U2 ( .A1(I[1]), .A2(I[0]), .ZN(n7) );
  AND3_X1 U3 ( .A1(n7), .A2(I[2]), .A3(n6), .ZN(O[2]) );
  AOI21_X1 U4 ( .B1(n7), .B2(n6), .A(I[2]), .ZN(O[0]) );
  MUX2_X1 U5 ( .A(n7), .B(n6), .S(I[2]), .Z(n5) );
  INV_X1 U6 ( .A(n5), .ZN(O[1]) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net46712, net148457, net148418, net138085, net138084, n3;
  assign Co = net46712;

  OAI21_X1 U1 ( .B1(n3), .B2(net138084), .A(net138085), .ZN(net46712) );
  NAND2_X1 U2 ( .A1(net148418), .A2(net148457), .ZN(net138085) );
  CLKBUF_X1 U3 ( .A(B), .Z(net148457) );
  CLKBUF_X1 U4 ( .A(A), .Z(net148418) );
  INV_X1 U5 ( .A(Ci), .ZN(net138084) );
  XNOR2_X1 U6 ( .A(A), .B(B), .ZN(n3) );
  XNOR2_X1 U7 ( .A(n3), .B(Ci), .ZN(S) );
endmodule


module BOOTHMUL_N32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [63:0] A;
  input [63:0] B;
  output [63:0] SUM;
  input CI;
  output CO;
  wire   \carry[61] , \carry[60] , \carry[59] , \carry[58] , \carry[57] ,
         \carry[56] , \carry[55] , \carry[54] , \carry[53] , \carry[52] ,
         \carry[51] , \carry[50] , \carry[49] , \carry[48] , \carry[47] ,
         \carry[46] , \carry[45] , \carry[44] , \carry[43] , \carry[42] ,
         \carry[41] , \carry[40] , \carry[39] , \carry[38] , \carry[37] ,
         \carry[36] , \carry[35] , \carry[34] , \carry[33] , \carry[32] ,
         \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] , \carry[62] , n1;

  XOR2_X1 U7 ( .A(A[60]), .B(\carry[60] ), .Z(SUM[60]) );
  XOR2_X1 U9 ( .A(A[59]), .B(\carry[59] ), .Z(SUM[59]) );
  XOR2_X1 U11 ( .A(A[58]), .B(\carry[58] ), .Z(SUM[58]) );
  XOR2_X1 U13 ( .A(A[57]), .B(\carry[57] ), .Z(SUM[57]) );
  XOR2_X1 U15 ( .A(A[56]), .B(\carry[56] ), .Z(SUM[56]) );
  XOR2_X1 U17 ( .A(A[55]), .B(\carry[55] ), .Z(SUM[55]) );
  XOR2_X1 U19 ( .A(A[54]), .B(\carry[54] ), .Z(SUM[54]) );
  XOR2_X1 U21 ( .A(A[53]), .B(\carry[53] ), .Z(SUM[53]) );
  XOR2_X1 U23 ( .A(A[52]), .B(\carry[52] ), .Z(SUM[52]) );
  XOR2_X1 U25 ( .A(A[51]), .B(\carry[51] ), .Z(SUM[51]) );
  XOR2_X1 U27 ( .A(A[50]), .B(\carry[50] ), .Z(SUM[50]) );
  XOR2_X1 U29 ( .A(A[49]), .B(\carry[49] ), .Z(SUM[49]) );
  XOR2_X1 U31 ( .A(A[48]), .B(\carry[48] ), .Z(SUM[48]) );
  XOR2_X1 U33 ( .A(A[47]), .B(\carry[47] ), .Z(SUM[47]) );
  XOR2_X1 U35 ( .A(A[46]), .B(\carry[46] ), .Z(SUM[46]) );
  XOR2_X1 U37 ( .A(A[45]), .B(\carry[45] ), .Z(SUM[45]) );
  XOR2_X1 U39 ( .A(A[44]), .B(\carry[44] ), .Z(SUM[44]) );
  XOR2_X1 U41 ( .A(A[43]), .B(\carry[43] ), .Z(SUM[43]) );
  XOR2_X1 U43 ( .A(A[42]), .B(\carry[42] ), .Z(SUM[42]) );
  XOR2_X1 U45 ( .A(A[41]), .B(\carry[41] ), .Z(SUM[41]) );
  XOR2_X1 U47 ( .A(A[40]), .B(\carry[40] ), .Z(SUM[40]) );
  XOR2_X1 U49 ( .A(A[39]), .B(\carry[39] ), .Z(SUM[39]) );
  XOR2_X1 U51 ( .A(A[38]), .B(\carry[38] ), .Z(SUM[38]) );
  XOR2_X1 U53 ( .A(A[37]), .B(\carry[37] ), .Z(SUM[37]) );
  XOR2_X1 U55 ( .A(A[36]), .B(\carry[36] ), .Z(SUM[36]) );
  XOR2_X1 U57 ( .A(A[35]), .B(\carry[35] ), .Z(SUM[35]) );
  XOR2_X1 U59 ( .A(A[34]), .B(\carry[34] ), .Z(SUM[34]) );
  XOR2_X1 U61 ( .A(A[33]), .B(\carry[33] ), .Z(SUM[33]) );
  XOR2_X1 U63 ( .A(A[32]), .B(\carry[32] ), .Z(SUM[32]) );
  XOR2_X1 U65 ( .A(A[31]), .B(\carry[31] ), .Z(SUM[31]) );
  XOR2_X1 U67 ( .A(A[30]), .B(\carry[30] ), .Z(SUM[30]) );
  XOR2_X1 U69 ( .A(A[29]), .B(\carry[29] ), .Z(SUM[29]) );
  XOR2_X1 U71 ( .A(A[28]), .B(\carry[28] ), .Z(SUM[28]) );
  XOR2_X1 U73 ( .A(A[27]), .B(\carry[27] ), .Z(SUM[27]) );
  XOR2_X1 U75 ( .A(A[26]), .B(\carry[26] ), .Z(SUM[26]) );
  XOR2_X1 U77 ( .A(A[25]), .B(\carry[25] ), .Z(SUM[25]) );
  XOR2_X1 U79 ( .A(A[24]), .B(\carry[24] ), .Z(SUM[24]) );
  XOR2_X1 U81 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  XOR2_X1 U83 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  XOR2_X1 U85 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  XOR2_X1 U87 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  XOR2_X1 U89 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  XOR2_X1 U91 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  XOR2_X1 U93 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  XOR2_X1 U95 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  XOR2_X1 U97 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  XOR2_X1 U99 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  XOR2_X1 U101 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  XOR2_X1 U103 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  XOR2_X1 U105 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  XOR2_X1 U107 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  XOR2_X1 U109 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
  XOR2_X1 U111 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  XOR2_X1 U113 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  XOR2_X1 U115 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  XOR2_X1 U117 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  XOR2_X1 U119 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  XOR2_X1 U121 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  XOR2_X1 U123 ( .A(A[2]), .B(\carry[2] ), .Z(SUM[2]) );
  XOR2_X1 U125 ( .A(A[1]), .B(\carry[1] ), .Z(SUM[1]) );
  XOR2_X1 U127 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  XOR2_X1 U5 ( .A(A[61]), .B(\carry[61] ), .Z(SUM[61]) );
  XOR2_X1 U3 ( .A(\carry[62] ), .B(A[62]), .Z(SUM[62]) );
  AND2_X1 U1 ( .A1(A[61]), .A2(\carry[61] ), .ZN(\carry[62] ) );
  XNOR2_X1 U2 ( .A(A[63]), .B(n1), .ZN(SUM[63]) );
  NAND2_X1 U4 ( .A1(\carry[62] ), .A2(A[62]), .ZN(n1) );
  AND2_X1 U6 ( .A1(\carry[57] ), .A2(A[57]), .ZN(\carry[58] ) );
  AND2_X1 U8 ( .A1(A[56]), .A2(\carry[56] ), .ZN(\carry[57] ) );
  AND2_X1 U10 ( .A1(A[54]), .A2(\carry[54] ), .ZN(\carry[55] ) );
  AND2_X1 U12 ( .A1(A[55]), .A2(\carry[55] ), .ZN(\carry[56] ) );
  AND2_X1 U14 ( .A1(\carry[53] ), .A2(A[53]), .ZN(\carry[54] ) );
  AND2_X1 U16 ( .A1(\carry[52] ), .A2(A[52]), .ZN(\carry[53] ) );
  AND2_X1 U18 ( .A1(\carry[51] ), .A2(A[51]), .ZN(\carry[52] ) );
  AND2_X1 U20 ( .A1(A[50]), .A2(\carry[50] ), .ZN(\carry[51] ) );
  AND2_X1 U22 ( .A1(\carry[49] ), .A2(A[49]), .ZN(\carry[50] ) );
  AND2_X1 U24 ( .A1(\carry[46] ), .A2(A[46]), .ZN(\carry[47] ) );
  AND2_X1 U26 ( .A1(\carry[41] ), .A2(A[41]), .ZN(\carry[42] ) );
  AND2_X1 U28 ( .A1(\carry[40] ), .A2(A[40]), .ZN(\carry[41] ) );
  AND2_X1 U30 ( .A1(\carry[39] ), .A2(A[39]), .ZN(\carry[40] ) );
  AND2_X1 U32 ( .A1(\carry[37] ), .A2(A[37]), .ZN(\carry[38] ) );
  AND2_X1 U34 ( .A1(\carry[35] ), .A2(A[35]), .ZN(\carry[36] ) );
  AND2_X1 U36 ( .A1(\carry[25] ), .A2(A[25]), .ZN(\carry[26] ) );
  AND2_X1 U38 ( .A1(\carry[24] ), .A2(A[24]), .ZN(\carry[25] ) );
  AND2_X1 U40 ( .A1(\carry[60] ), .A2(A[60]), .ZN(\carry[61] ) );
  AND2_X1 U42 ( .A1(A[58]), .A2(\carry[58] ), .ZN(\carry[59] ) );
  AND2_X1 U44 ( .A1(\carry[59] ), .A2(A[59]), .ZN(\carry[60] ) );
  AND2_X1 U46 ( .A1(\carry[48] ), .A2(A[48]), .ZN(\carry[49] ) );
  AND2_X1 U48 ( .A1(A[47]), .A2(\carry[47] ), .ZN(\carry[48] ) );
  AND2_X1 U50 ( .A1(\carry[45] ), .A2(A[45]), .ZN(\carry[46] ) );
  AND2_X1 U52 ( .A1(\carry[44] ), .A2(A[44]), .ZN(\carry[45] ) );
  AND2_X1 U54 ( .A1(\carry[43] ), .A2(A[43]), .ZN(\carry[44] ) );
  AND2_X1 U56 ( .A1(\carry[42] ), .A2(A[42]), .ZN(\carry[43] ) );
  AND2_X1 U58 ( .A1(\carry[38] ), .A2(A[38]), .ZN(\carry[39] ) );
  AND2_X1 U60 ( .A1(\carry[36] ), .A2(A[36]), .ZN(\carry[37] ) );
  AND2_X1 U62 ( .A1(\carry[34] ), .A2(A[34]), .ZN(\carry[35] ) );
  AND2_X1 U64 ( .A1(\carry[33] ), .A2(A[33]), .ZN(\carry[34] ) );
  AND2_X1 U66 ( .A1(\carry[32] ), .A2(A[32]), .ZN(\carry[33] ) );
  AND2_X1 U68 ( .A1(\carry[31] ), .A2(A[31]), .ZN(\carry[32] ) );
  AND2_X1 U70 ( .A1(\carry[29] ), .A2(A[29]), .ZN(\carry[30] ) );
  AND2_X1 U72 ( .A1(\carry[30] ), .A2(A[30]), .ZN(\carry[31] ) );
  AND2_X1 U74 ( .A1(\carry[28] ), .A2(A[28]), .ZN(\carry[29] ) );
  AND2_X1 U76 ( .A1(\carry[27] ), .A2(A[27]), .ZN(\carry[28] ) );
  AND2_X1 U78 ( .A1(\carry[26] ), .A2(A[26]), .ZN(\carry[27] ) );
  AND2_X1 U80 ( .A1(\carry[23] ), .A2(A[23]), .ZN(\carry[24] ) );
  AND2_X1 U82 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  AND2_X1 U84 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  AND2_X1 U86 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  AND2_X1 U88 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  AND2_X1 U90 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  AND2_X1 U92 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  AND2_X1 U94 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  AND2_X1 U96 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  AND2_X1 U98 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  AND2_X1 U100 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  AND2_X1 U102 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  AND2_X1 U104 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  AND2_X1 U106 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  AND2_X1 U108 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  AND2_X1 U110 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  AND2_X1 U112 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  AND2_X1 U114 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  AND2_X1 U116 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  AND2_X1 U118 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
  AND2_X1 U120 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  AND2_X1 U122 ( .A1(\carry[2] ), .A2(A[2]), .ZN(\carry[3] ) );
  AND2_X1 U124 ( .A1(\carry[1] ), .A2(A[1]), .ZN(\carry[2] ) );
  AND2_X1 U126 ( .A1(A[0]), .A2(B[0]), .ZN(\carry[1] ) );
endmodule


module RCA_generic_N64_0 ( A, B, Ci, S, Co );
  input [63:0] A;
  input [63:0] B;
  output [63:0] S;
  input Ci;
  output Co;

  wire   [63:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1007 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1006 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1005 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_1004 FAI_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_1003 FAI_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_1002 FAI_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_1001 FAI_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_1000 FAI_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_999 FAI_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_998 FAI_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11]) );
  FA_997 FAI_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12]) );
  FA_996 FAI_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13]) );
  FA_995 FAI_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14]) );
  FA_994 FAI_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15]) );
  FA_993 FAI_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16]) );
  FA_992 FAI_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17]) );
  FA_991 FAI_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18]) );
  FA_990 FAI_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19]) );
  FA_989 FAI_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20]) );
  FA_988 FAI_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21]) );
  FA_987 FAI_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22]) );
  FA_986 FAI_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23]) );
  FA_985 FAI_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24]) );
  FA_984 FAI_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25]) );
  FA_983 FAI_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26]) );
  FA_982 FAI_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27]) );
  FA_981 FAI_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28]) );
  FA_980 FAI_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29]) );
  FA_979 FAI_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30]) );
  FA_978 FAI_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31]) );
  FA_977 FAI_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(CTMP[32]) );
  FA_976 FAI_33 ( .A(A[32]), .B(B[32]), .Ci(CTMP[32]), .S(S[32]), .Co(CTMP[33]) );
  FA_975 FAI_34 ( .A(A[33]), .B(B[33]), .Ci(CTMP[33]), .S(S[33]), .Co(CTMP[34]) );
  FA_974 FAI_35 ( .A(A[34]), .B(B[34]), .Ci(CTMP[34]), .S(S[34]), .Co(CTMP[35]) );
  FA_973 FAI_36 ( .A(A[35]), .B(B[35]), .Ci(CTMP[35]), .S(S[35]), .Co(CTMP[36]) );
  FA_972 FAI_37 ( .A(A[36]), .B(B[36]), .Ci(CTMP[36]), .S(S[36]), .Co(CTMP[37]) );
  FA_971 FAI_38 ( .A(A[37]), .B(B[37]), .Ci(CTMP[37]), .S(S[37]), .Co(CTMP[38]) );
  FA_970 FAI_39 ( .A(A[38]), .B(B[38]), .Ci(CTMP[38]), .S(S[38]), .Co(CTMP[39]) );
  FA_969 FAI_40 ( .A(A[39]), .B(B[39]), .Ci(CTMP[39]), .S(S[39]), .Co(CTMP[40]) );
  FA_968 FAI_41 ( .A(A[40]), .B(B[40]), .Ci(CTMP[40]), .S(S[40]), .Co(CTMP[41]) );
  FA_967 FAI_42 ( .A(A[41]), .B(B[41]), .Ci(CTMP[41]), .S(S[41]), .Co(CTMP[42]) );
  FA_966 FAI_43 ( .A(A[42]), .B(B[42]), .Ci(CTMP[42]), .S(S[42]), .Co(CTMP[43]) );
  FA_965 FAI_44 ( .A(A[43]), .B(B[43]), .Ci(CTMP[43]), .S(S[43]), .Co(CTMP[44]) );
  FA_964 FAI_45 ( .A(A[44]), .B(B[44]), .Ci(CTMP[44]), .S(S[44]), .Co(CTMP[45]) );
  FA_963 FAI_46 ( .A(A[45]), .B(B[45]), .Ci(CTMP[45]), .S(S[45]), .Co(CTMP[46]) );
  FA_962 FAI_47 ( .A(A[46]), .B(B[46]), .Ci(CTMP[46]), .S(S[46]), .Co(CTMP[47]) );
  FA_961 FAI_48 ( .A(A[47]), .B(B[47]), .Ci(CTMP[47]), .S(S[47]), .Co(CTMP[48]) );
  FA_960 FAI_49 ( .A(A[48]), .B(B[48]), .Ci(CTMP[48]), .S(S[48]), .Co(CTMP[49]) );
  FA_959 FAI_50 ( .A(A[49]), .B(B[49]), .Ci(CTMP[49]), .S(S[49]), .Co(CTMP[50]) );
  FA_958 FAI_51 ( .A(A[50]), .B(B[50]), .Ci(CTMP[50]), .S(S[50]), .Co(CTMP[51]) );
  FA_957 FAI_52 ( .A(A[51]), .B(B[51]), .Ci(CTMP[51]), .S(S[51]), .Co(CTMP[52]) );
  FA_956 FAI_53 ( .A(A[52]), .B(B[52]), .Ci(CTMP[52]), .S(S[52]), .Co(CTMP[53]) );
  FA_955 FAI_54 ( .A(A[53]), .B(B[53]), .Ci(CTMP[53]), .S(S[53]), .Co(CTMP[54]) );
  FA_954 FAI_55 ( .A(A[54]), .B(B[54]), .Ci(CTMP[54]), .S(S[54]), .Co(CTMP[55]) );
  FA_953 FAI_56 ( .A(A[55]), .B(B[55]), .Ci(CTMP[55]), .S(S[55]), .Co(CTMP[56]) );
  FA_952 FAI_57 ( .A(A[56]), .B(B[56]), .Ci(CTMP[56]), .S(S[56]), .Co(CTMP[57]) );
  FA_951 FAI_58 ( .A(A[57]), .B(B[57]), .Ci(CTMP[57]), .S(S[57]), .Co(CTMP[58]) );
  FA_950 FAI_59 ( .A(A[58]), .B(B[58]), .Ci(CTMP[58]), .S(S[58]), .Co(CTMP[59]) );
  FA_949 FAI_60 ( .A(A[59]), .B(B[59]), .Ci(CTMP[59]), .S(S[59]), .Co(CTMP[60]) );
  FA_948 FAI_61 ( .A(A[60]), .B(B[60]), .Ci(CTMP[60]), .S(S[60]), .Co(CTMP[61]) );
  FA_947 FAI_62 ( .A(A[61]), .B(B[61]), .Ci(CTMP[61]), .S(S[61]), .Co(CTMP[62]) );
  FA_946 FAI_63 ( .A(A[62]), .B(B[62]), .Ci(CTMP[62]), .S(S[62]), .Co(CTMP[63]) );
  FA_945 FAI_64 ( .A(A[63]), .B(B[63]), .Ci(CTMP[63]), .S(S[63]), .Co(Co) );
endmodule


module MUX51_GENERIC_N64_0 ( A, B, C, D, E, SEL, Y );
  input [63:0] A;
  input [63:0] B;
  input [63:0] C;
  input [63:0] D;
  input [63:0] E;
  input [2:0] SEL;
  output [63:0] Y;
  wire   net142158, net142406, net145869, net145867, net145865, net145863,
         net145879, net145875, net145893, net145891, net145889, net145887,
         net145885, net145903, net145901, net145899, net145897, net145917,
         net145915, net145909, net148517, net148599, net158795, net157198,
         net148598, net145883, net142411, net142410, net142409, net149357,
         net148545, net148525, net148524, net142421, net142420, net142417,
         net142415, net142414, net142412, net142408, net149341, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395;

  BUF_X2 U1 ( .A(n142), .Z(net145903) );
  INV_X1 U2 ( .A(net142412), .ZN(n139) );
  CLKBUF_X1 U3 ( .A(SEL[0]), .Z(net149357) );
  BUF_X1 U4 ( .A(n140), .Z(net145875) );
  AND2_X1 U5 ( .A1(net142420), .A2(net142417), .ZN(n140) );
  OR2_X1 U6 ( .A1(net148525), .A2(n143), .ZN(n144) );
  CLKBUF_X1 U7 ( .A(SEL[1]), .Z(n141) );
  INV_X1 U8 ( .A(net142415), .ZN(n142) );
  CLKBUF_X1 U9 ( .A(net142158), .Z(net145897) );
  AND2_X1 U10 ( .A1(net157198), .A2(E[0]), .ZN(net149341) );
  NAND2_X1 U11 ( .A1(net148545), .A2(net149341), .ZN(net142408) );
  AND4_X1 U12 ( .A1(net157198), .A2(net142415), .A3(net142412), .A4(net142414), 
        .ZN(net148517) );
  INV_X1 U13 ( .A(n144), .ZN(net148599) );
  INV_X1 U14 ( .A(SEL[1]), .ZN(n143) );
  OR2_X1 U15 ( .A1(n143), .A2(net148525), .ZN(net157198) );
  NAND3_X1 U16 ( .A1(n143), .A2(net149357), .A3(net142421), .ZN(net142415) );
  AND3_X1 U17 ( .A1(SEL[1]), .A2(net149357), .A3(net142421), .ZN(net158795) );
  NAND3_X1 U18 ( .A1(n141), .A2(net149357), .A3(net142421), .ZN(net142414) );
  NOR2_X1 U19 ( .A1(SEL[2]), .A2(SEL[1]), .ZN(net142420) );
  NAND4_X1 U20 ( .A1(net142408), .A2(net142411), .A3(net142410), .A4(net142409), .ZN(Y[0]) );
  AND3_X1 U21 ( .A1(net142415), .A2(net142412), .A3(net142414), .ZN(net148545)
         );
  INV_X1 U22 ( .A(SEL[2]), .ZN(net142421) );
  INV_X1 U23 ( .A(net142415), .ZN(net142158) );
  NAND2_X1 U24 ( .A1(net142420), .A2(net142417), .ZN(net142412) );
  INV_X1 U25 ( .A(SEL[0]), .ZN(net142417) );
  NAND2_X1 U26 ( .A1(net142417), .A2(net148524), .ZN(net148525) );
  INV_X1 U27 ( .A(SEL[2]), .ZN(net148524) );
  NAND2_X1 U28 ( .A1(B[0]), .A2(net142158), .ZN(net142409) );
  NAND2_X1 U29 ( .A1(D[0]), .A2(net145883), .ZN(net142410) );
  BUF_X1 U30 ( .A(net158795), .Z(net145883) );
  NAND2_X1 U31 ( .A1(D[1]), .A2(net145883), .ZN(net142406) );
  AOI22_X1 U32 ( .A1(net148598), .A2(C[0]), .B1(n139), .B2(A[0]), .ZN(
        net142411) );
  INV_X1 U33 ( .A(n144), .ZN(net148598) );
  CLKBUF_X1 U34 ( .A(net148599), .Z(net145867) );
  BUF_X4 U35 ( .A(net148599), .Z(net145865) );
  CLKBUF_X3 U36 ( .A(net148517), .Z(net145909) );
  BUF_X4 U37 ( .A(n140), .Z(net145879) );
  BUF_X1 U38 ( .A(net158795), .Z(net145885) );
  BUF_X1 U39 ( .A(net158795), .Z(net145887) );
  CLKBUF_X2 U40 ( .A(net148517), .Z(net145915) );
  CLKBUF_X1 U41 ( .A(n142), .Z(net145901) );
  CLKBUF_X1 U42 ( .A(net158795), .Z(net145889) );
  CLKBUF_X1 U43 ( .A(net158795), .Z(net145891) );
  CLKBUF_X1 U44 ( .A(n142), .Z(net145899) );
  CLKBUF_X1 U45 ( .A(net148599), .Z(net145863) );
  CLKBUF_X1 U46 ( .A(net148517), .Z(net145917) );
  CLKBUF_X1 U47 ( .A(net158795), .Z(net145893) );
  CLKBUF_X1 U48 ( .A(net148599), .Z(net145869) );
  NAND2_X1 U49 ( .A1(E[1]), .A2(net148517), .ZN(n147) );
  NAND2_X1 U50 ( .A1(B[1]), .A2(net142158), .ZN(n146) );
  AOI22_X1 U51 ( .A1(C[1]), .A2(net148599), .B1(A[1]), .B2(n140), .ZN(n145) );
  NAND4_X1 U52 ( .A1(n147), .A2(n146), .A3(net142406), .A4(n145), .ZN(Y[1]) );
  NAND2_X1 U53 ( .A1(E[2]), .A2(net145917), .ZN(n151) );
  NAND2_X1 U54 ( .A1(B[2]), .A2(n142), .ZN(n150) );
  NAND2_X1 U55 ( .A1(D[2]), .A2(net145887), .ZN(n149) );
  AOI22_X1 U56 ( .A1(C[2]), .A2(net145867), .B1(A[2]), .B2(n140), .ZN(n148) );
  NAND4_X1 U57 ( .A1(n151), .A2(n150), .A3(n149), .A4(n148), .ZN(Y[2]) );
  NAND2_X1 U58 ( .A1(E[3]), .A2(net145909), .ZN(n155) );
  NAND2_X1 U59 ( .A1(B[3]), .A2(net145897), .ZN(n154) );
  NAND2_X1 U60 ( .A1(D[3]), .A2(net145885), .ZN(n153) );
  AOI22_X1 U61 ( .A1(C[3]), .A2(net145863), .B1(A[3]), .B2(net145875), .ZN(
        n152) );
  NAND4_X1 U62 ( .A1(n155), .A2(n154), .A3(n153), .A4(n152), .ZN(Y[3]) );
  NAND2_X1 U63 ( .A1(E[4]), .A2(net145909), .ZN(n159) );
  NAND2_X1 U64 ( .A1(B[4]), .A2(net145899), .ZN(n158) );
  NAND2_X1 U65 ( .A1(D[4]), .A2(net145893), .ZN(n157) );
  AOI22_X1 U66 ( .A1(C[4]), .A2(net145863), .B1(A[4]), .B2(net145875), .ZN(
        n156) );
  NAND4_X1 U67 ( .A1(n159), .A2(n158), .A3(n157), .A4(n156), .ZN(Y[4]) );
  NAND2_X1 U68 ( .A1(E[5]), .A2(net145909), .ZN(n163) );
  NAND2_X1 U69 ( .A1(B[5]), .A2(net145901), .ZN(n162) );
  NAND2_X1 U70 ( .A1(D[5]), .A2(net145891), .ZN(n161) );
  AOI22_X1 U71 ( .A1(C[5]), .A2(net145865), .B1(A[5]), .B2(net145875), .ZN(
        n160) );
  NAND4_X1 U72 ( .A1(n163), .A2(n162), .A3(n161), .A4(n160), .ZN(Y[5]) );
  NAND2_X1 U73 ( .A1(E[6]), .A2(net145915), .ZN(n167) );
  NAND2_X1 U74 ( .A1(B[6]), .A2(net145903), .ZN(n166) );
  NAND2_X1 U75 ( .A1(D[6]), .A2(net145889), .ZN(n165) );
  AOI22_X1 U76 ( .A1(C[6]), .A2(net145869), .B1(A[6]), .B2(net145875), .ZN(
        n164) );
  NAND4_X1 U77 ( .A1(n167), .A2(n166), .A3(n165), .A4(n164), .ZN(Y[6]) );
  NAND2_X1 U78 ( .A1(E[7]), .A2(net145915), .ZN(n171) );
  NAND2_X1 U79 ( .A1(B[7]), .A2(net145903), .ZN(n170) );
  NAND2_X1 U80 ( .A1(D[7]), .A2(net145887), .ZN(n169) );
  AOI22_X1 U81 ( .A1(C[7]), .A2(net145865), .B1(A[7]), .B2(net145875), .ZN(
        n168) );
  NAND4_X1 U82 ( .A1(n171), .A2(n170), .A3(n169), .A4(n168), .ZN(Y[7]) );
  NAND2_X1 U83 ( .A1(E[8]), .A2(net145915), .ZN(n175) );
  NAND2_X1 U84 ( .A1(B[8]), .A2(net145903), .ZN(n174) );
  NAND2_X1 U85 ( .A1(D[8]), .A2(net145885), .ZN(n173) );
  AOI22_X1 U86 ( .A1(C[8]), .A2(net145865), .B1(A[8]), .B2(net145879), .ZN(
        n172) );
  NAND4_X1 U87 ( .A1(n175), .A2(n174), .A3(n173), .A4(n172), .ZN(Y[8]) );
  NAND2_X1 U88 ( .A1(E[9]), .A2(net145915), .ZN(n179) );
  NAND2_X1 U89 ( .A1(B[9]), .A2(net145903), .ZN(n178) );
  NAND2_X1 U90 ( .A1(D[9]), .A2(net145893), .ZN(n177) );
  AOI22_X1 U91 ( .A1(C[9]), .A2(net145865), .B1(A[9]), .B2(net145879), .ZN(
        n176) );
  NAND4_X1 U92 ( .A1(n179), .A2(n178), .A3(n177), .A4(n176), .ZN(Y[9]) );
  NAND2_X1 U93 ( .A1(E[10]), .A2(net145915), .ZN(n183) );
  NAND2_X1 U94 ( .A1(B[10]), .A2(net145903), .ZN(n182) );
  NAND2_X1 U95 ( .A1(D[10]), .A2(net145891), .ZN(n181) );
  AOI22_X1 U96 ( .A1(C[10]), .A2(net145865), .B1(A[10]), .B2(net145879), .ZN(
        n180) );
  NAND4_X1 U97 ( .A1(n183), .A2(n182), .A3(n181), .A4(n180), .ZN(Y[10]) );
  NAND2_X1 U98 ( .A1(E[11]), .A2(net145915), .ZN(n187) );
  NAND2_X1 U99 ( .A1(B[11]), .A2(net145903), .ZN(n186) );
  NAND2_X1 U100 ( .A1(D[11]), .A2(net145889), .ZN(n185) );
  AOI22_X1 U101 ( .A1(C[11]), .A2(net145865), .B1(A[11]), .B2(net145879), .ZN(
        n184) );
  NAND4_X1 U102 ( .A1(n187), .A2(n186), .A3(n185), .A4(n184), .ZN(Y[11]) );
  NAND2_X1 U103 ( .A1(E[12]), .A2(net145915), .ZN(n191) );
  NAND2_X1 U104 ( .A1(B[12]), .A2(net145897), .ZN(n190) );
  NAND2_X1 U105 ( .A1(D[12]), .A2(net145887), .ZN(n189) );
  AOI22_X1 U106 ( .A1(C[12]), .A2(net145865), .B1(A[12]), .B2(net145879), .ZN(
        n188) );
  NAND4_X1 U107 ( .A1(n191), .A2(n190), .A3(n189), .A4(n188), .ZN(Y[12]) );
  NAND2_X1 U108 ( .A1(E[13]), .A2(net145915), .ZN(n195) );
  NAND2_X1 U109 ( .A1(B[13]), .A2(net145897), .ZN(n194) );
  NAND2_X1 U110 ( .A1(D[13]), .A2(net145885), .ZN(n193) );
  AOI22_X1 U111 ( .A1(C[13]), .A2(net145865), .B1(A[13]), .B2(net145879), .ZN(
        n192) );
  NAND4_X1 U112 ( .A1(n195), .A2(n194), .A3(n193), .A4(n192), .ZN(Y[13]) );
  NAND2_X1 U113 ( .A1(E[14]), .A2(net145915), .ZN(n199) );
  NAND2_X1 U114 ( .A1(B[14]), .A2(net145897), .ZN(n198) );
  NAND2_X1 U115 ( .A1(D[14]), .A2(net145893), .ZN(n197) );
  AOI22_X1 U116 ( .A1(C[14]), .A2(net145865), .B1(A[14]), .B2(net145879), .ZN(
        n196) );
  NAND4_X1 U117 ( .A1(n199), .A2(n198), .A3(n197), .A4(n196), .ZN(Y[14]) );
  NAND2_X1 U118 ( .A1(E[15]), .A2(net145915), .ZN(n203) );
  NAND2_X1 U119 ( .A1(B[15]), .A2(net145897), .ZN(n202) );
  NAND2_X1 U120 ( .A1(D[15]), .A2(net145891), .ZN(n201) );
  AOI22_X1 U121 ( .A1(C[15]), .A2(net145865), .B1(A[15]), .B2(net145879), .ZN(
        n200) );
  NAND4_X1 U122 ( .A1(n203), .A2(n202), .A3(n201), .A4(n200), .ZN(Y[15]) );
  NAND2_X1 U123 ( .A1(E[16]), .A2(net145915), .ZN(n207) );
  NAND2_X1 U124 ( .A1(B[16]), .A2(net145897), .ZN(n206) );
  NAND2_X1 U125 ( .A1(D[16]), .A2(net145889), .ZN(n205) );
  AOI22_X1 U126 ( .A1(C[16]), .A2(net145865), .B1(A[16]), .B2(net145879), .ZN(
        n204) );
  NAND4_X1 U127 ( .A1(n207), .A2(n206), .A3(n205), .A4(n204), .ZN(Y[16]) );
  NAND2_X1 U128 ( .A1(E[17]), .A2(net145915), .ZN(n211) );
  NAND2_X1 U129 ( .A1(B[17]), .A2(net145897), .ZN(n210) );
  NAND2_X1 U130 ( .A1(D[17]), .A2(net145887), .ZN(n209) );
  AOI22_X1 U131 ( .A1(C[17]), .A2(net145865), .B1(A[17]), .B2(net145879), .ZN(
        n208) );
  NAND4_X1 U132 ( .A1(n211), .A2(n210), .A3(n209), .A4(n208), .ZN(Y[17]) );
  NAND2_X1 U133 ( .A1(E[18]), .A2(net145915), .ZN(n215) );
  NAND2_X1 U134 ( .A1(B[18]), .A2(net145897), .ZN(n214) );
  NAND2_X1 U135 ( .A1(D[18]), .A2(net145885), .ZN(n213) );
  AOI22_X1 U136 ( .A1(C[18]), .A2(net145869), .B1(A[18]), .B2(net145879), .ZN(
        n212) );
  NAND4_X1 U137 ( .A1(n215), .A2(n214), .A3(n213), .A4(n212), .ZN(Y[18]) );
  NAND2_X1 U138 ( .A1(E[19]), .A2(net145915), .ZN(n219) );
  NAND2_X1 U139 ( .A1(B[19]), .A2(net145897), .ZN(n218) );
  NAND2_X1 U140 ( .A1(D[19]), .A2(net145893), .ZN(n217) );
  AOI22_X1 U141 ( .A1(C[19]), .A2(net145869), .B1(A[19]), .B2(net145879), .ZN(
        n216) );
  NAND4_X1 U142 ( .A1(n219), .A2(n218), .A3(n217), .A4(n216), .ZN(Y[19]) );
  NAND2_X1 U143 ( .A1(E[20]), .A2(net145915), .ZN(n223) );
  NAND2_X1 U144 ( .A1(B[20]), .A2(net145897), .ZN(n222) );
  NAND2_X1 U145 ( .A1(D[20]), .A2(net145891), .ZN(n221) );
  AOI22_X1 U146 ( .A1(C[20]), .A2(net145865), .B1(A[20]), .B2(net145879), .ZN(
        n220) );
  NAND4_X1 U147 ( .A1(n223), .A2(n222), .A3(n221), .A4(n220), .ZN(Y[20]) );
  NAND2_X1 U148 ( .A1(E[21]), .A2(net145915), .ZN(n227) );
  NAND2_X1 U149 ( .A1(B[21]), .A2(net145897), .ZN(n226) );
  NAND2_X1 U150 ( .A1(D[21]), .A2(net145889), .ZN(n225) );
  AOI22_X1 U151 ( .A1(C[21]), .A2(net145869), .B1(A[21]), .B2(net145879), .ZN(
        n224) );
  NAND4_X1 U152 ( .A1(n227), .A2(n226), .A3(n225), .A4(n224), .ZN(Y[21]) );
  NAND2_X1 U153 ( .A1(E[22]), .A2(net145915), .ZN(n231) );
  NAND2_X1 U154 ( .A1(B[22]), .A2(net145897), .ZN(n230) );
  NAND2_X1 U155 ( .A1(D[22]), .A2(net145887), .ZN(n229) );
  AOI22_X1 U156 ( .A1(C[22]), .A2(net145865), .B1(A[22]), .B2(net145879), .ZN(
        n228) );
  NAND4_X1 U157 ( .A1(n231), .A2(n230), .A3(n229), .A4(n228), .ZN(Y[22]) );
  NAND2_X1 U158 ( .A1(E[23]), .A2(net145915), .ZN(n235) );
  NAND2_X1 U159 ( .A1(B[23]), .A2(net145897), .ZN(n234) );
  NAND2_X1 U160 ( .A1(D[23]), .A2(net145885), .ZN(n233) );
  AOI22_X1 U161 ( .A1(C[23]), .A2(net145869), .B1(A[23]), .B2(net145879), .ZN(
        n232) );
  NAND4_X1 U162 ( .A1(n235), .A2(n234), .A3(n233), .A4(n232), .ZN(Y[23]) );
  NAND2_X1 U163 ( .A1(E[24]), .A2(net145915), .ZN(n239) );
  NAND2_X1 U164 ( .A1(B[24]), .A2(net145899), .ZN(n238) );
  NAND2_X1 U165 ( .A1(D[24]), .A2(net145893), .ZN(n237) );
  AOI22_X1 U166 ( .A1(C[24]), .A2(net145865), .B1(A[24]), .B2(net145879), .ZN(
        n236) );
  NAND4_X1 U167 ( .A1(n239), .A2(n238), .A3(n237), .A4(n236), .ZN(Y[24]) );
  NAND2_X1 U168 ( .A1(E[25]), .A2(net145915), .ZN(n243) );
  NAND2_X1 U169 ( .A1(B[25]), .A2(net145899), .ZN(n242) );
  NAND2_X1 U170 ( .A1(D[25]), .A2(net145891), .ZN(n241) );
  AOI22_X1 U171 ( .A1(C[25]), .A2(net145869), .B1(A[25]), .B2(net145879), .ZN(
        n240) );
  NAND4_X1 U172 ( .A1(n243), .A2(n242), .A3(n241), .A4(n240), .ZN(Y[25]) );
  NAND2_X1 U173 ( .A1(E[26]), .A2(net145915), .ZN(n247) );
  NAND2_X1 U174 ( .A1(B[26]), .A2(net145899), .ZN(n246) );
  NAND2_X1 U175 ( .A1(D[26]), .A2(net145889), .ZN(n245) );
  AOI22_X1 U176 ( .A1(C[26]), .A2(net145865), .B1(A[26]), .B2(net145879), .ZN(
        n244) );
  NAND4_X1 U177 ( .A1(n247), .A2(n246), .A3(n245), .A4(n244), .ZN(Y[26]) );
  NAND2_X1 U178 ( .A1(E[27]), .A2(net145915), .ZN(n251) );
  NAND2_X1 U179 ( .A1(B[27]), .A2(net145899), .ZN(n250) );
  NAND2_X1 U180 ( .A1(D[27]), .A2(net145887), .ZN(n249) );
  AOI22_X1 U181 ( .A1(C[27]), .A2(net145869), .B1(A[27]), .B2(net145879), .ZN(
        n248) );
  NAND4_X1 U182 ( .A1(n251), .A2(n250), .A3(n249), .A4(n248), .ZN(Y[27]) );
  NAND2_X1 U183 ( .A1(E[28]), .A2(net145915), .ZN(n255) );
  NAND2_X1 U184 ( .A1(B[28]), .A2(net145899), .ZN(n254) );
  NAND2_X1 U185 ( .A1(D[28]), .A2(net145885), .ZN(n253) );
  AOI22_X1 U186 ( .A1(C[28]), .A2(net145865), .B1(A[28]), .B2(net145879), .ZN(
        n252) );
  NAND4_X1 U187 ( .A1(n255), .A2(n254), .A3(n253), .A4(n252), .ZN(Y[28]) );
  NAND2_X1 U188 ( .A1(E[29]), .A2(net145915), .ZN(n259) );
  NAND2_X1 U189 ( .A1(B[29]), .A2(net145899), .ZN(n258) );
  NAND2_X1 U190 ( .A1(D[29]), .A2(net145893), .ZN(n257) );
  AOI22_X1 U191 ( .A1(C[29]), .A2(net145869), .B1(A[29]), .B2(net145879), .ZN(
        n256) );
  NAND4_X1 U192 ( .A1(n259), .A2(n258), .A3(n257), .A4(n256), .ZN(Y[29]) );
  NAND2_X1 U193 ( .A1(E[30]), .A2(net145915), .ZN(n263) );
  NAND2_X1 U194 ( .A1(B[30]), .A2(net145899), .ZN(n262) );
  NAND2_X1 U195 ( .A1(D[30]), .A2(net145891), .ZN(n261) );
  AOI22_X1 U196 ( .A1(C[30]), .A2(net145865), .B1(A[30]), .B2(net145879), .ZN(
        n260) );
  NAND4_X1 U197 ( .A1(n263), .A2(n262), .A3(n261), .A4(n260), .ZN(Y[30]) );
  NAND2_X1 U198 ( .A1(E[31]), .A2(net145915), .ZN(n267) );
  NAND2_X1 U199 ( .A1(B[31]), .A2(net145899), .ZN(n266) );
  NAND2_X1 U200 ( .A1(D[31]), .A2(net145889), .ZN(n265) );
  AOI22_X1 U201 ( .A1(C[31]), .A2(net145869), .B1(A[31]), .B2(net145879), .ZN(
        n264) );
  NAND4_X1 U202 ( .A1(n267), .A2(n266), .A3(n265), .A4(n264), .ZN(Y[31]) );
  NAND2_X1 U203 ( .A1(E[32]), .A2(net145915), .ZN(n271) );
  NAND2_X1 U204 ( .A1(B[32]), .A2(net145899), .ZN(n270) );
  NAND2_X1 U205 ( .A1(D[32]), .A2(net145887), .ZN(n269) );
  AOI22_X1 U206 ( .A1(C[32]), .A2(net145865), .B1(A[32]), .B2(net145879), .ZN(
        n268) );
  NAND4_X1 U207 ( .A1(n271), .A2(n270), .A3(n269), .A4(n268), .ZN(Y[32]) );
  NAND2_X1 U208 ( .A1(E[33]), .A2(net145909), .ZN(n275) );
  NAND2_X1 U209 ( .A1(B[33]), .A2(net145899), .ZN(n274) );
  NAND2_X1 U210 ( .A1(D[33]), .A2(net145885), .ZN(n273) );
  AOI22_X1 U211 ( .A1(C[33]), .A2(net145869), .B1(A[33]), .B2(net145879), .ZN(
        n272) );
  NAND4_X1 U212 ( .A1(n275), .A2(n274), .A3(n273), .A4(n272), .ZN(Y[33]) );
  NAND2_X1 U213 ( .A1(E[34]), .A2(net145915), .ZN(n279) );
  NAND2_X1 U214 ( .A1(B[34]), .A2(net145899), .ZN(n278) );
  NAND2_X1 U215 ( .A1(D[34]), .A2(net145893), .ZN(n277) );
  AOI22_X1 U216 ( .A1(C[34]), .A2(net145869), .B1(A[34]), .B2(net145879), .ZN(
        n276) );
  NAND4_X1 U217 ( .A1(n279), .A2(n278), .A3(n277), .A4(n276), .ZN(Y[34]) );
  NAND2_X1 U218 ( .A1(E[35]), .A2(net145909), .ZN(n283) );
  NAND2_X1 U219 ( .A1(B[35]), .A2(net145899), .ZN(n282) );
  NAND2_X1 U220 ( .A1(D[35]), .A2(net145891), .ZN(n281) );
  AOI22_X1 U221 ( .A1(C[35]), .A2(net145865), .B1(A[35]), .B2(net145879), .ZN(
        n280) );
  NAND4_X1 U222 ( .A1(n283), .A2(n282), .A3(n281), .A4(n280), .ZN(Y[35]) );
  NAND2_X1 U223 ( .A1(E[36]), .A2(net145915), .ZN(n287) );
  NAND2_X1 U224 ( .A1(B[36]), .A2(net145901), .ZN(n286) );
  NAND2_X1 U225 ( .A1(D[36]), .A2(net145889), .ZN(n285) );
  AOI22_X1 U226 ( .A1(C[36]), .A2(net145865), .B1(A[36]), .B2(net145879), .ZN(
        n284) );
  NAND4_X1 U227 ( .A1(n287), .A2(n286), .A3(n285), .A4(n284), .ZN(Y[36]) );
  NAND2_X1 U228 ( .A1(E[37]), .A2(net145909), .ZN(n291) );
  NAND2_X1 U229 ( .A1(B[37]), .A2(net145901), .ZN(n290) );
  NAND2_X1 U230 ( .A1(D[37]), .A2(net145887), .ZN(n289) );
  AOI22_X1 U231 ( .A1(C[37]), .A2(net145865), .B1(A[37]), .B2(net145879), .ZN(
        n288) );
  NAND4_X1 U232 ( .A1(n291), .A2(n290), .A3(n289), .A4(n288), .ZN(Y[37]) );
  NAND2_X1 U233 ( .A1(E[38]), .A2(net145915), .ZN(n295) );
  NAND2_X1 U234 ( .A1(B[38]), .A2(net145901), .ZN(n294) );
  NAND2_X1 U235 ( .A1(D[38]), .A2(net145885), .ZN(n293) );
  AOI22_X1 U236 ( .A1(C[38]), .A2(net145869), .B1(A[38]), .B2(net145879), .ZN(
        n292) );
  NAND4_X1 U237 ( .A1(n295), .A2(n294), .A3(n293), .A4(n292), .ZN(Y[38]) );
  NAND2_X1 U238 ( .A1(E[39]), .A2(net145909), .ZN(n299) );
  NAND2_X1 U239 ( .A1(B[39]), .A2(net145901), .ZN(n298) );
  NAND2_X1 U240 ( .A1(D[39]), .A2(net145893), .ZN(n297) );
  AOI22_X1 U241 ( .A1(C[39]), .A2(net145865), .B1(A[39]), .B2(net145879), .ZN(
        n296) );
  NAND4_X1 U242 ( .A1(n299), .A2(n298), .A3(n297), .A4(n296), .ZN(Y[39]) );
  NAND2_X1 U243 ( .A1(E[40]), .A2(net145915), .ZN(n303) );
  NAND2_X1 U244 ( .A1(B[40]), .A2(net145901), .ZN(n302) );
  NAND2_X1 U245 ( .A1(D[40]), .A2(net145891), .ZN(n301) );
  AOI22_X1 U246 ( .A1(C[40]), .A2(net145865), .B1(A[40]), .B2(net145879), .ZN(
        n300) );
  NAND4_X1 U247 ( .A1(n303), .A2(n302), .A3(n301), .A4(n300), .ZN(Y[40]) );
  NAND2_X1 U248 ( .A1(E[41]), .A2(net145909), .ZN(n307) );
  NAND2_X1 U249 ( .A1(B[41]), .A2(net145901), .ZN(n306) );
  NAND2_X1 U250 ( .A1(D[41]), .A2(net145889), .ZN(n305) );
  AOI22_X1 U251 ( .A1(C[41]), .A2(net145865), .B1(A[41]), .B2(net145879), .ZN(
        n304) );
  NAND4_X1 U252 ( .A1(n307), .A2(n306), .A3(n305), .A4(n304), .ZN(Y[41]) );
  NAND2_X1 U253 ( .A1(E[42]), .A2(net145915), .ZN(n311) );
  NAND2_X1 U254 ( .A1(B[42]), .A2(net145901), .ZN(n310) );
  NAND2_X1 U255 ( .A1(D[42]), .A2(net145887), .ZN(n309) );
  AOI22_X1 U256 ( .A1(C[42]), .A2(net145869), .B1(A[42]), .B2(net145879), .ZN(
        n308) );
  NAND4_X1 U257 ( .A1(n311), .A2(n310), .A3(n309), .A4(n308), .ZN(Y[42]) );
  NAND2_X1 U258 ( .A1(E[43]), .A2(net145909), .ZN(n315) );
  NAND2_X1 U259 ( .A1(B[43]), .A2(net145901), .ZN(n314) );
  NAND2_X1 U260 ( .A1(D[43]), .A2(net145885), .ZN(n313) );
  AOI22_X1 U261 ( .A1(C[43]), .A2(net145865), .B1(A[43]), .B2(net145879), .ZN(
        n312) );
  NAND4_X1 U262 ( .A1(n315), .A2(n314), .A3(n313), .A4(n312), .ZN(Y[43]) );
  NAND2_X1 U263 ( .A1(E[44]), .A2(net145915), .ZN(n319) );
  NAND2_X1 U264 ( .A1(B[44]), .A2(net145901), .ZN(n318) );
  NAND2_X1 U265 ( .A1(D[44]), .A2(net145893), .ZN(n317) );
  AOI22_X1 U266 ( .A1(C[44]), .A2(net145865), .B1(A[44]), .B2(net145879), .ZN(
        n316) );
  NAND4_X1 U267 ( .A1(n319), .A2(n318), .A3(n317), .A4(n316), .ZN(Y[44]) );
  NAND2_X1 U268 ( .A1(E[45]), .A2(net145915), .ZN(n323) );
  NAND2_X1 U269 ( .A1(B[45]), .A2(net145901), .ZN(n322) );
  NAND2_X1 U270 ( .A1(D[45]), .A2(net145891), .ZN(n321) );
  AOI22_X1 U271 ( .A1(C[45]), .A2(net145869), .B1(A[45]), .B2(net145879), .ZN(
        n320) );
  NAND4_X1 U272 ( .A1(n323), .A2(n322), .A3(n321), .A4(n320), .ZN(Y[45]) );
  NAND2_X1 U273 ( .A1(E[46]), .A2(net145909), .ZN(n327) );
  NAND2_X1 U274 ( .A1(B[46]), .A2(net145901), .ZN(n326) );
  NAND2_X1 U275 ( .A1(D[46]), .A2(net145889), .ZN(n325) );
  AOI22_X1 U276 ( .A1(C[46]), .A2(net145865), .B1(A[46]), .B2(net145879), .ZN(
        n324) );
  NAND4_X1 U277 ( .A1(n327), .A2(n326), .A3(n325), .A4(n324), .ZN(Y[46]) );
  NAND2_X1 U278 ( .A1(E[47]), .A2(net145909), .ZN(n331) );
  NAND2_X1 U279 ( .A1(B[47]), .A2(net145901), .ZN(n330) );
  NAND2_X1 U280 ( .A1(D[47]), .A2(net145887), .ZN(n329) );
  AOI22_X1 U281 ( .A1(C[47]), .A2(net145865), .B1(A[47]), .B2(net145875), .ZN(
        n328) );
  NAND4_X1 U282 ( .A1(n331), .A2(n330), .A3(n329), .A4(n328), .ZN(Y[47]) );
  NAND2_X1 U283 ( .A1(E[48]), .A2(net145909), .ZN(n335) );
  NAND2_X1 U284 ( .A1(B[48]), .A2(net145903), .ZN(n334) );
  NAND2_X1 U285 ( .A1(D[48]), .A2(net145885), .ZN(n333) );
  AOI22_X1 U286 ( .A1(C[48]), .A2(net145869), .B1(A[48]), .B2(net145879), .ZN(
        n332) );
  NAND4_X1 U287 ( .A1(n335), .A2(n334), .A3(n333), .A4(n332), .ZN(Y[48]) );
  NAND2_X1 U288 ( .A1(E[49]), .A2(net145909), .ZN(n339) );
  NAND2_X1 U289 ( .A1(B[49]), .A2(net145903), .ZN(n338) );
  NAND2_X1 U290 ( .A1(D[49]), .A2(net145893), .ZN(n337) );
  AOI22_X1 U291 ( .A1(C[49]), .A2(net145865), .B1(A[49]), .B2(net145879), .ZN(
        n336) );
  NAND4_X1 U292 ( .A1(n339), .A2(n338), .A3(n337), .A4(n336), .ZN(Y[49]) );
  NAND2_X1 U293 ( .A1(E[50]), .A2(net145915), .ZN(n343) );
  NAND2_X1 U294 ( .A1(B[50]), .A2(net145903), .ZN(n342) );
  NAND2_X1 U295 ( .A1(D[50]), .A2(net145891), .ZN(n341) );
  AOI22_X1 U296 ( .A1(C[50]), .A2(net145865), .B1(A[50]), .B2(net145879), .ZN(
        n340) );
  NAND4_X1 U297 ( .A1(n343), .A2(n342), .A3(n341), .A4(n340), .ZN(Y[50]) );
  NAND2_X1 U298 ( .A1(E[51]), .A2(net145909), .ZN(n347) );
  NAND2_X1 U299 ( .A1(B[51]), .A2(net145903), .ZN(n346) );
  NAND2_X1 U300 ( .A1(D[51]), .A2(net145889), .ZN(n345) );
  AOI22_X1 U301 ( .A1(C[51]), .A2(net145869), .B1(A[51]), .B2(net145879), .ZN(
        n344) );
  NAND4_X1 U302 ( .A1(n347), .A2(n346), .A3(n345), .A4(n344), .ZN(Y[51]) );
  NAND2_X1 U303 ( .A1(E[52]), .A2(net145915), .ZN(n351) );
  NAND2_X1 U304 ( .A1(B[52]), .A2(net145903), .ZN(n350) );
  NAND2_X1 U305 ( .A1(D[52]), .A2(net145887), .ZN(n349) );
  AOI22_X1 U306 ( .A1(C[52]), .A2(net145865), .B1(A[52]), .B2(net145875), .ZN(
        n348) );
  NAND4_X1 U307 ( .A1(n351), .A2(n350), .A3(n349), .A4(n348), .ZN(Y[52]) );
  NAND2_X1 U308 ( .A1(E[53]), .A2(net145915), .ZN(n355) );
  NAND2_X1 U309 ( .A1(B[53]), .A2(net145903), .ZN(n354) );
  NAND2_X1 U310 ( .A1(D[53]), .A2(net145885), .ZN(n353) );
  AOI22_X1 U311 ( .A1(C[53]), .A2(net145865), .B1(A[53]), .B2(net145879), .ZN(
        n352) );
  NAND4_X1 U312 ( .A1(n355), .A2(n354), .A3(n353), .A4(n352), .ZN(Y[53]) );
  NAND2_X1 U313 ( .A1(E[54]), .A2(net145909), .ZN(n359) );
  NAND2_X1 U314 ( .A1(B[54]), .A2(net145903), .ZN(n358) );
  NAND2_X1 U315 ( .A1(D[54]), .A2(net145893), .ZN(n357) );
  AOI22_X1 U316 ( .A1(C[54]), .A2(net145863), .B1(A[54]), .B2(net145879), .ZN(
        n356) );
  NAND4_X1 U317 ( .A1(n359), .A2(n358), .A3(n357), .A4(n356), .ZN(Y[54]) );
  NAND2_X1 U318 ( .A1(E[55]), .A2(net145915), .ZN(n363) );
  NAND2_X1 U319 ( .A1(B[55]), .A2(net145903), .ZN(n362) );
  NAND2_X1 U320 ( .A1(D[55]), .A2(net145891), .ZN(n361) );
  AOI22_X1 U321 ( .A1(C[55]), .A2(net145865), .B1(A[55]), .B2(net145879), .ZN(
        n360) );
  NAND4_X1 U322 ( .A1(n363), .A2(n362), .A3(n361), .A4(n360), .ZN(Y[55]) );
  NAND2_X1 U323 ( .A1(E[56]), .A2(net145909), .ZN(n367) );
  NAND2_X1 U324 ( .A1(B[56]), .A2(net145903), .ZN(n366) );
  NAND2_X1 U325 ( .A1(D[56]), .A2(net145889), .ZN(n365) );
  AOI22_X1 U326 ( .A1(C[56]), .A2(net145869), .B1(A[56]), .B2(net145879), .ZN(
        n364) );
  NAND4_X1 U327 ( .A1(n367), .A2(n366), .A3(n365), .A4(n364), .ZN(Y[56]) );
  NAND2_X1 U328 ( .A1(E[57]), .A2(net145915), .ZN(n371) );
  NAND2_X1 U329 ( .A1(B[57]), .A2(net145903), .ZN(n370) );
  NAND2_X1 U330 ( .A1(D[57]), .A2(net145887), .ZN(n369) );
  AOI22_X1 U331 ( .A1(C[57]), .A2(net145865), .B1(A[57]), .B2(net145879), .ZN(
        n368) );
  NAND4_X1 U332 ( .A1(n371), .A2(n370), .A3(n369), .A4(n368), .ZN(Y[57]) );
  NAND2_X1 U333 ( .A1(E[58]), .A2(net145909), .ZN(n375) );
  NAND2_X1 U334 ( .A1(B[58]), .A2(net145903), .ZN(n374) );
  NAND2_X1 U335 ( .A1(D[58]), .A2(net145885), .ZN(n373) );
  AOI22_X1 U336 ( .A1(C[58]), .A2(net145865), .B1(A[58]), .B2(net145879), .ZN(
        n372) );
  NAND4_X1 U337 ( .A1(n375), .A2(n374), .A3(n373), .A4(n372), .ZN(Y[58]) );
  NAND2_X1 U338 ( .A1(E[59]), .A2(net145915), .ZN(n379) );
  NAND2_X1 U339 ( .A1(B[59]), .A2(net145903), .ZN(n378) );
  NAND2_X1 U340 ( .A1(D[59]), .A2(net145893), .ZN(n377) );
  AOI22_X1 U341 ( .A1(C[59]), .A2(net145863), .B1(A[59]), .B2(net145875), .ZN(
        n376) );
  NAND4_X1 U342 ( .A1(n379), .A2(n378), .A3(n377), .A4(n376), .ZN(Y[59]) );
  NAND2_X1 U343 ( .A1(E[60]), .A2(net145909), .ZN(n383) );
  NAND2_X1 U344 ( .A1(B[60]), .A2(net145903), .ZN(n382) );
  NAND2_X1 U345 ( .A1(D[60]), .A2(net145891), .ZN(n381) );
  AOI22_X1 U346 ( .A1(C[60]), .A2(net145869), .B1(A[60]), .B2(net145879), .ZN(
        n380) );
  NAND4_X1 U347 ( .A1(n383), .A2(n382), .A3(n381), .A4(n380), .ZN(Y[60]) );
  NAND2_X1 U348 ( .A1(E[61]), .A2(net145915), .ZN(n387) );
  NAND2_X1 U349 ( .A1(B[61]), .A2(net145903), .ZN(n386) );
  NAND2_X1 U350 ( .A1(D[61]), .A2(net145889), .ZN(n385) );
  AOI22_X1 U351 ( .A1(C[61]), .A2(net145863), .B1(A[61]), .B2(net145879), .ZN(
        n384) );
  NAND4_X1 U352 ( .A1(n387), .A2(n386), .A3(n385), .A4(n384), .ZN(Y[61]) );
  NAND2_X1 U353 ( .A1(E[62]), .A2(net145909), .ZN(n391) );
  NAND2_X1 U354 ( .A1(B[62]), .A2(net145903), .ZN(n390) );
  NAND2_X1 U355 ( .A1(D[62]), .A2(net145887), .ZN(n389) );
  AOI22_X1 U356 ( .A1(C[62]), .A2(net145865), .B1(A[62]), .B2(net145879), .ZN(
        n388) );
  NAND4_X1 U357 ( .A1(n391), .A2(n390), .A3(n389), .A4(n388), .ZN(Y[62]) );
  NAND2_X1 U358 ( .A1(E[63]), .A2(net145915), .ZN(n395) );
  NAND2_X1 U359 ( .A1(B[63]), .A2(net145901), .ZN(n394) );
  NAND2_X1 U360 ( .A1(D[63]), .A2(net145885), .ZN(n393) );
  AOI22_X1 U361 ( .A1(C[63]), .A2(net145865), .B1(A[63]), .B2(net145879), .ZN(
        n392) );
  NAND4_X1 U362 ( .A1(n395), .A2(n394), .A3(n393), .A4(n392), .ZN(Y[63]) );
endmodule


module BOOTH_ENCODER_4 ( I, O );
  input [2:0] I;
  output [2:0] O;
  wire   net142483, net147588, net156612, net158600, net158628, net158612,
         net158610, net158606, net158605, n4;
  assign O[2] = net147588;
  assign O[1] = net158628;

  NAND2_X1 U1 ( .A1(net158610), .A2(net158612), .ZN(net158606) );
  INV_X1 U2 ( .A(I[0]), .ZN(net158612) );
  NAND2_X1 U3 ( .A1(I[1]), .A2(I[0]), .ZN(n4) );
  XNOR2_X1 U4 ( .A(n4), .B(I[2]), .ZN(net158605) );
  AND2_X2 U5 ( .A1(net158605), .A2(net158606), .ZN(net158628) );
  INV_X1 U6 ( .A(I[1]), .ZN(net158610) );
  AOI21_X1 U7 ( .B1(net156612), .B2(net142483), .A(I[2]), .ZN(O[0]) );
  AND3_X2 U8 ( .A1(net158600), .A2(I[2]), .A3(net142483), .ZN(net147588) );
  NAND2_X1 U9 ( .A1(I[0]), .A2(I[1]), .ZN(net142483) );
  XNOR2_X1 U10 ( .A(I[1]), .B(I[0]), .ZN(net158600) );
  XNOR2_X1 U11 ( .A(I[1]), .B(I[0]), .ZN(net156612) );
endmodule


module BOOTHMUL_N32 ( A, B, P );
  input [31:0] A;
  input [31:0] B;
  output [63:0] P;
  wire   \mux_out[7][63] , \mux_out[7][62] , \mux_out[7][61] ,
         \mux_out[7][60] , \mux_out[7][59] , \mux_out[7][58] ,
         \mux_out[7][57] , \mux_out[7][56] , \mux_out[7][55] ,
         \mux_out[7][54] , \mux_out[7][53] , \mux_out[7][52] ,
         \mux_out[7][51] , \mux_out[7][50] , \mux_out[7][49] ,
         \mux_out[7][48] , \mux_out[7][47] , \mux_out[7][46] ,
         \mux_out[7][45] , \mux_out[7][44] , \mux_out[7][43] ,
         \mux_out[7][42] , \mux_out[7][41] , \mux_out[7][40] ,
         \mux_out[7][39] , \mux_out[7][38] , \mux_out[7][37] ,
         \mux_out[7][36] , \mux_out[7][35] , \mux_out[7][34] ,
         \mux_out[7][33] , \mux_out[7][32] , \mux_out[7][31] ,
         \mux_out[7][30] , \mux_out[7][29] , \mux_out[7][28] ,
         \mux_out[7][27] , \mux_out[7][26] , \mux_out[7][25] ,
         \mux_out[7][24] , \mux_out[7][23] , \mux_out[7][22] ,
         \mux_out[7][21] , \mux_out[7][20] , \mux_out[7][19] ,
         \mux_out[7][18] , \mux_out[7][17] , \mux_out[7][16] ,
         \mux_out[7][15] , \mux_out[7][14] , \mux_out[7][13] ,
         \mux_out[7][12] , \mux_out[7][11] , \mux_out[7][10] , \mux_out[7][9] ,
         \mux_out[7][8] , \mux_out[7][7] , \mux_out[7][6] , \mux_out[7][5] ,
         \mux_out[7][4] , \mux_out[7][3] , \mux_out[7][2] , \mux_out[7][1] ,
         \mux_out[7][0] , \mux_out[6][63] , \mux_out[6][62] , \mux_out[6][61] ,
         \mux_out[6][60] , \mux_out[6][59] , \mux_out[6][58] ,
         \mux_out[6][57] , \mux_out[6][56] , \mux_out[6][55] ,
         \mux_out[6][54] , \mux_out[6][53] , \mux_out[6][52] ,
         \mux_out[6][51] , \mux_out[6][50] , \mux_out[6][49] ,
         \mux_out[6][48] , \mux_out[6][47] , \mux_out[6][46] ,
         \mux_out[6][45] , \mux_out[6][44] , \mux_out[6][43] ,
         \mux_out[6][42] , \mux_out[6][41] , \mux_out[6][40] ,
         \mux_out[6][39] , \mux_out[6][38] , \mux_out[6][37] ,
         \mux_out[6][36] , \mux_out[6][35] , \mux_out[6][34] ,
         \mux_out[6][33] , \mux_out[6][32] , \mux_out[6][31] ,
         \mux_out[6][30] , \mux_out[6][29] , \mux_out[6][28] ,
         \mux_out[6][27] , \mux_out[6][26] , \mux_out[6][25] ,
         \mux_out[6][24] , \mux_out[6][23] , \mux_out[6][22] ,
         \mux_out[6][21] , \mux_out[6][20] , \mux_out[6][19] ,
         \mux_out[6][18] , \mux_out[6][17] , \mux_out[6][16] ,
         \mux_out[6][15] , \mux_out[6][14] , \mux_out[6][13] ,
         \mux_out[6][12] , \mux_out[6][11] , \mux_out[6][10] , \mux_out[6][9] ,
         \mux_out[6][8] , \mux_out[6][7] , \mux_out[6][6] , \mux_out[6][5] ,
         \mux_out[6][4] , \mux_out[6][3] , \mux_out[6][2] , \mux_out[6][1] ,
         \mux_out[6][0] , \mux_out[5][63] , \mux_out[5][62] , \mux_out[5][61] ,
         \mux_out[5][60] , \mux_out[5][59] , \mux_out[5][58] ,
         \mux_out[5][57] , \mux_out[5][56] , \mux_out[5][55] ,
         \mux_out[5][54] , \mux_out[5][53] , \mux_out[5][52] ,
         \mux_out[5][51] , \mux_out[5][50] , \mux_out[5][49] ,
         \mux_out[5][48] , \mux_out[5][47] , \mux_out[5][46] ,
         \mux_out[5][45] , \mux_out[5][44] , \mux_out[5][43] ,
         \mux_out[5][42] , \mux_out[5][41] , \mux_out[5][40] ,
         \mux_out[5][39] , \mux_out[5][38] , \mux_out[5][37] ,
         \mux_out[5][36] , \mux_out[5][35] , \mux_out[5][34] ,
         \mux_out[5][33] , \mux_out[5][32] , \mux_out[5][31] ,
         \mux_out[5][30] , \mux_out[5][29] , \mux_out[5][28] ,
         \mux_out[5][27] , \mux_out[5][26] , \mux_out[5][25] ,
         \mux_out[5][24] , \mux_out[5][23] , \mux_out[5][22] ,
         \mux_out[5][21] , \mux_out[5][20] , \mux_out[5][19] ,
         \mux_out[5][18] , \mux_out[5][17] , \mux_out[5][16] ,
         \mux_out[5][15] , \mux_out[5][14] , \mux_out[5][13] ,
         \mux_out[5][12] , \mux_out[5][11] , \mux_out[5][10] , \mux_out[5][9] ,
         \mux_out[5][8] , \mux_out[5][7] , \mux_out[5][6] , \mux_out[5][5] ,
         \mux_out[5][4] , \mux_out[5][3] , \mux_out[5][2] , \mux_out[5][1] ,
         \mux_out[5][0] , \mux_out[4][63] , \mux_out[4][62] , \mux_out[4][61] ,
         \mux_out[4][60] , \mux_out[4][59] , \mux_out[4][58] ,
         \mux_out[4][57] , \mux_out[4][56] , \mux_out[4][55] ,
         \mux_out[4][54] , \mux_out[4][53] , \mux_out[4][52] ,
         \mux_out[4][51] , \mux_out[4][50] , \mux_out[4][49] ,
         \mux_out[4][48] , \mux_out[4][47] , \mux_out[4][46] ,
         \mux_out[4][45] , \mux_out[4][44] , \mux_out[4][43] ,
         \mux_out[4][42] , \mux_out[4][41] , \mux_out[4][40] ,
         \mux_out[4][39] , \mux_out[4][38] , \mux_out[4][37] ,
         \mux_out[4][36] , \mux_out[4][35] , \mux_out[4][34] ,
         \mux_out[4][33] , \mux_out[4][32] , \mux_out[4][31] ,
         \mux_out[4][30] , \mux_out[4][29] , \mux_out[4][28] ,
         \mux_out[4][27] , \mux_out[4][26] , \mux_out[4][25] ,
         \mux_out[4][24] , \mux_out[4][23] , \mux_out[4][22] ,
         \mux_out[4][21] , \mux_out[4][20] , \mux_out[4][19] ,
         \mux_out[4][18] , \mux_out[4][17] , \mux_out[4][16] ,
         \mux_out[4][15] , \mux_out[4][14] , \mux_out[4][13] ,
         \mux_out[4][12] , \mux_out[4][11] , \mux_out[4][10] , \mux_out[4][9] ,
         \mux_out[4][8] , \mux_out[4][7] , \mux_out[4][6] , \mux_out[4][5] ,
         \mux_out[4][4] , \mux_out[4][3] , \mux_out[4][2] , \mux_out[4][1] ,
         \mux_out[4][0] , \mux_out[3][63] , \mux_out[3][62] , \mux_out[3][61] ,
         \mux_out[3][60] , \mux_out[3][59] , \mux_out[3][58] ,
         \mux_out[3][57] , \mux_out[3][56] , \mux_out[3][55] ,
         \mux_out[3][54] , \mux_out[3][53] , \mux_out[3][52] ,
         \mux_out[3][51] , \mux_out[3][50] , \mux_out[3][49] ,
         \mux_out[3][48] , \mux_out[3][47] , \mux_out[3][46] ,
         \mux_out[3][45] , \mux_out[3][44] , \mux_out[3][43] ,
         \mux_out[3][42] , \mux_out[3][41] , \mux_out[3][40] ,
         \mux_out[3][39] , \mux_out[3][38] , \mux_out[3][37] ,
         \mux_out[3][36] , \mux_out[3][35] , \mux_out[3][34] ,
         \mux_out[3][33] , \mux_out[3][32] , \mux_out[3][31] ,
         \mux_out[3][30] , \mux_out[3][29] , \mux_out[3][28] ,
         \mux_out[3][27] , \mux_out[3][26] , \mux_out[3][25] ,
         \mux_out[3][24] , \mux_out[3][23] , \mux_out[3][22] ,
         \mux_out[3][21] , \mux_out[3][20] , \mux_out[3][19] ,
         \mux_out[3][18] , \mux_out[3][17] , \mux_out[3][16] ,
         \mux_out[3][15] , \mux_out[3][14] , \mux_out[3][13] ,
         \mux_out[3][12] , \mux_out[3][11] , \mux_out[3][10] , \mux_out[3][9] ,
         \mux_out[3][8] , \mux_out[3][7] , \mux_out[3][6] , \mux_out[3][5] ,
         \mux_out[3][4] , \mux_out[3][3] , \mux_out[3][2] , \mux_out[3][1] ,
         \mux_out[3][0] , \mux_out[2][63] , \mux_out[2][62] , \mux_out[2][61] ,
         \mux_out[2][60] , \mux_out[2][59] , \mux_out[2][58] ,
         \mux_out[2][57] , \mux_out[2][56] , \mux_out[2][55] ,
         \mux_out[2][54] , \mux_out[2][53] , \mux_out[2][52] ,
         \mux_out[2][51] , \mux_out[2][50] , \mux_out[2][49] ,
         \mux_out[2][48] , \mux_out[2][47] , \mux_out[2][46] ,
         \mux_out[2][45] , \mux_out[2][44] , \mux_out[2][43] ,
         \mux_out[2][42] , \mux_out[2][41] , \mux_out[2][40] ,
         \mux_out[2][39] , \mux_out[2][38] , \mux_out[2][37] ,
         \mux_out[2][36] , \mux_out[2][35] , \mux_out[2][34] ,
         \mux_out[2][33] , \mux_out[2][32] , \mux_out[2][31] ,
         \mux_out[2][30] , \mux_out[2][29] , \mux_out[2][28] ,
         \mux_out[2][27] , \mux_out[2][26] , \mux_out[2][25] ,
         \mux_out[2][24] , \mux_out[2][23] , \mux_out[2][22] ,
         \mux_out[2][21] , \mux_out[2][20] , \mux_out[2][19] ,
         \mux_out[2][18] , \mux_out[2][17] , \mux_out[2][16] ,
         \mux_out[2][15] , \mux_out[2][14] , \mux_out[2][13] ,
         \mux_out[2][12] , \mux_out[2][11] , \mux_out[2][10] , \mux_out[2][9] ,
         \mux_out[2][8] , \mux_out[2][7] , \mux_out[2][6] , \mux_out[2][5] ,
         \mux_out[2][4] , \mux_out[2][3] , \mux_out[2][2] , \mux_out[2][1] ,
         \mux_out[2][0] , \mux_out[1][63] , \mux_out[1][62] , \mux_out[1][61] ,
         \mux_out[1][60] , \mux_out[1][59] , \mux_out[1][58] ,
         \mux_out[1][57] , \mux_out[1][56] , \mux_out[1][55] ,
         \mux_out[1][54] , \mux_out[1][53] , \mux_out[1][52] ,
         \mux_out[1][51] , \mux_out[1][50] , \mux_out[1][49] ,
         \mux_out[1][48] , \mux_out[1][47] , \mux_out[1][46] ,
         \mux_out[1][45] , \mux_out[1][44] , \mux_out[1][43] ,
         \mux_out[1][42] , \mux_out[1][41] , \mux_out[1][40] ,
         \mux_out[1][39] , \mux_out[1][38] , \mux_out[1][37] ,
         \mux_out[1][36] , \mux_out[1][35] , \mux_out[1][34] ,
         \mux_out[1][33] , \mux_out[1][32] , \mux_out[1][31] ,
         \mux_out[1][30] , \mux_out[1][29] , \mux_out[1][28] ,
         \mux_out[1][27] , \mux_out[1][26] , \mux_out[1][25] ,
         \mux_out[1][24] , \mux_out[1][23] , \mux_out[1][22] ,
         \mux_out[1][21] , \mux_out[1][20] , \mux_out[1][19] ,
         \mux_out[1][18] , \mux_out[1][17] , \mux_out[1][16] ,
         \mux_out[1][15] , \mux_out[1][14] , \mux_out[1][13] ,
         \mux_out[1][12] , \mux_out[1][11] , \mux_out[1][10] , \mux_out[1][9] ,
         \mux_out[1][8] , \mux_out[1][7] , \mux_out[1][6] , \mux_out[1][5] ,
         \mux_out[1][4] , \mux_out[1][3] , \mux_out[1][2] , \mux_out[1][1] ,
         \mux_out[1][0] , \mux_out[15][63] , \mux_out[15][62] ,
         \mux_out[15][61] , \mux_out[15][60] , \mux_out[15][59] ,
         \mux_out[15][58] , \mux_out[15][57] , \mux_out[15][56] ,
         \mux_out[15][55] , \mux_out[15][54] , \mux_out[15][53] ,
         \mux_out[15][52] , \mux_out[15][51] , \mux_out[15][50] ,
         \mux_out[15][49] , \mux_out[15][48] , \mux_out[15][47] ,
         \mux_out[15][46] , \mux_out[15][45] , \mux_out[15][44] ,
         \mux_out[15][43] , \mux_out[15][42] , \mux_out[15][41] ,
         \mux_out[15][40] , \mux_out[15][39] , \mux_out[15][38] ,
         \mux_out[15][37] , \mux_out[15][36] , \mux_out[15][35] ,
         \mux_out[15][34] , \mux_out[15][33] , \mux_out[15][32] ,
         \mux_out[15][31] , \mux_out[15][30] , \mux_out[15][29] ,
         \mux_out[15][28] , \mux_out[15][27] , \mux_out[15][26] ,
         \mux_out[15][25] , \mux_out[15][24] , \mux_out[15][23] ,
         \mux_out[15][22] , \mux_out[15][21] , \mux_out[15][20] ,
         \mux_out[15][19] , \mux_out[15][18] , \mux_out[15][17] ,
         \mux_out[15][16] , \mux_out[15][15] , \mux_out[15][14] ,
         \mux_out[15][13] , \mux_out[15][12] , \mux_out[15][11] ,
         \mux_out[15][10] , \mux_out[15][9] , \mux_out[15][8] ,
         \mux_out[15][7] , \mux_out[15][6] , \mux_out[15][5] ,
         \mux_out[15][4] , \mux_out[15][3] , \mux_out[15][2] ,
         \mux_out[15][1] , \mux_out[15][0] , \mux_out[14][63] ,
         \mux_out[14][62] , \mux_out[14][61] , \mux_out[14][60] ,
         \mux_out[14][59] , \mux_out[14][58] , \mux_out[14][57] ,
         \mux_out[14][56] , \mux_out[14][55] , \mux_out[14][54] ,
         \mux_out[14][53] , \mux_out[14][52] , \mux_out[14][51] ,
         \mux_out[14][50] , \mux_out[14][49] , \mux_out[14][48] ,
         \mux_out[14][47] , \mux_out[14][46] , \mux_out[14][45] ,
         \mux_out[14][44] , \mux_out[14][43] , \mux_out[14][42] ,
         \mux_out[14][41] , \mux_out[14][40] , \mux_out[14][39] ,
         \mux_out[14][38] , \mux_out[14][37] , \mux_out[14][36] ,
         \mux_out[14][35] , \mux_out[14][34] , \mux_out[14][33] ,
         \mux_out[14][32] , \mux_out[14][31] , \mux_out[14][30] ,
         \mux_out[14][29] , \mux_out[14][28] , \mux_out[14][27] ,
         \mux_out[14][26] , \mux_out[14][25] , \mux_out[14][24] ,
         \mux_out[14][23] , \mux_out[14][22] , \mux_out[14][21] ,
         \mux_out[14][20] , \mux_out[14][19] , \mux_out[14][18] ,
         \mux_out[14][17] , \mux_out[14][16] , \mux_out[14][15] ,
         \mux_out[14][14] , \mux_out[14][13] , \mux_out[14][12] ,
         \mux_out[14][11] , \mux_out[14][10] , \mux_out[14][9] ,
         \mux_out[14][8] , \mux_out[14][7] , \mux_out[14][6] ,
         \mux_out[14][5] , \mux_out[14][4] , \mux_out[14][3] ,
         \mux_out[14][2] , \mux_out[14][1] , \mux_out[14][0] ,
         \mux_out[13][63] , \mux_out[13][62] , \mux_out[13][61] ,
         \mux_out[13][60] , \mux_out[13][59] , \mux_out[13][58] ,
         \mux_out[13][57] , \mux_out[13][56] , \mux_out[13][55] ,
         \mux_out[13][54] , \mux_out[13][53] , \mux_out[13][52] ,
         \mux_out[13][51] , \mux_out[13][50] , \mux_out[13][49] ,
         \mux_out[13][48] , \mux_out[13][47] , \mux_out[13][46] ,
         \mux_out[13][45] , \mux_out[13][44] , \mux_out[13][43] ,
         \mux_out[13][42] , \mux_out[13][41] , \mux_out[13][40] ,
         \mux_out[13][39] , \mux_out[13][38] , \mux_out[13][37] ,
         \mux_out[13][36] , \mux_out[13][35] , \mux_out[13][34] ,
         \mux_out[13][33] , \mux_out[13][32] , \mux_out[13][31] ,
         \mux_out[13][30] , \mux_out[13][29] , \mux_out[13][28] ,
         \mux_out[13][27] , \mux_out[13][26] , \mux_out[13][25] ,
         \mux_out[13][24] , \mux_out[13][23] , \mux_out[13][22] ,
         \mux_out[13][21] , \mux_out[13][20] , \mux_out[13][19] ,
         \mux_out[13][18] , \mux_out[13][17] , \mux_out[13][16] ,
         \mux_out[13][15] , \mux_out[13][14] , \mux_out[13][13] ,
         \mux_out[13][12] , \mux_out[13][11] , \mux_out[13][10] ,
         \mux_out[13][9] , \mux_out[13][8] , \mux_out[13][7] ,
         \mux_out[13][6] , \mux_out[13][5] , \mux_out[13][4] ,
         \mux_out[13][3] , \mux_out[13][2] , \mux_out[13][1] ,
         \mux_out[13][0] , \mux_out[12][63] , \mux_out[12][62] ,
         \mux_out[12][61] , \mux_out[12][60] , \mux_out[12][59] ,
         \mux_out[12][58] , \mux_out[12][57] , \mux_out[12][56] ,
         \mux_out[12][55] , \mux_out[12][54] , \mux_out[12][53] ,
         \mux_out[12][52] , \mux_out[12][51] , \mux_out[12][50] ,
         \mux_out[12][49] , \mux_out[12][48] , \mux_out[12][47] ,
         \mux_out[12][46] , \mux_out[12][45] , \mux_out[12][44] ,
         \mux_out[12][43] , \mux_out[12][42] , \mux_out[12][41] ,
         \mux_out[12][40] , \mux_out[12][39] , \mux_out[12][38] ,
         \mux_out[12][37] , \mux_out[12][36] , \mux_out[12][35] ,
         \mux_out[12][34] , \mux_out[12][33] , \mux_out[12][32] ,
         \mux_out[12][31] , \mux_out[12][30] , \mux_out[12][29] ,
         \mux_out[12][28] , \mux_out[12][27] , \mux_out[12][26] ,
         \mux_out[12][25] , \mux_out[12][24] , \mux_out[12][23] ,
         \mux_out[12][22] , \mux_out[12][21] , \mux_out[12][20] ,
         \mux_out[12][19] , \mux_out[12][18] , \mux_out[12][17] ,
         \mux_out[12][16] , \mux_out[12][15] , \mux_out[12][14] ,
         \mux_out[12][13] , \mux_out[12][12] , \mux_out[12][11] ,
         \mux_out[12][10] , \mux_out[12][9] , \mux_out[12][8] ,
         \mux_out[12][7] , \mux_out[12][6] , \mux_out[12][5] ,
         \mux_out[12][4] , \mux_out[12][3] , \mux_out[12][2] ,
         \mux_out[12][1] , \mux_out[12][0] , \mux_out[11][63] ,
         \mux_out[11][62] , \mux_out[11][61] , \mux_out[11][60] ,
         \mux_out[11][59] , \mux_out[11][58] , \mux_out[11][57] ,
         \mux_out[11][56] , \mux_out[11][55] , \mux_out[11][54] ,
         \mux_out[11][53] , \mux_out[11][52] , \mux_out[11][51] ,
         \mux_out[11][50] , \mux_out[11][49] , \mux_out[11][48] ,
         \mux_out[11][47] , \mux_out[11][46] , \mux_out[11][45] ,
         \mux_out[11][44] , \mux_out[11][43] , \mux_out[11][42] ,
         \mux_out[11][41] , \mux_out[11][40] , \mux_out[11][39] ,
         \mux_out[11][38] , \mux_out[11][37] , \mux_out[11][36] ,
         \mux_out[11][35] , \mux_out[11][34] , \mux_out[11][33] ,
         \mux_out[11][32] , \mux_out[11][31] , \mux_out[11][30] ,
         \mux_out[11][29] , \mux_out[11][28] , \mux_out[11][27] ,
         \mux_out[11][26] , \mux_out[11][25] , \mux_out[11][24] ,
         \mux_out[11][23] , \mux_out[11][22] , \mux_out[11][21] ,
         \mux_out[11][20] , \mux_out[11][19] , \mux_out[11][18] ,
         \mux_out[11][17] , \mux_out[11][16] , \mux_out[11][15] ,
         \mux_out[11][14] , \mux_out[11][13] , \mux_out[11][12] ,
         \mux_out[11][11] , \mux_out[11][10] , \mux_out[11][9] ,
         \mux_out[11][8] , \mux_out[11][7] , \mux_out[11][6] ,
         \mux_out[11][5] , \mux_out[11][4] , \mux_out[11][3] ,
         \mux_out[11][2] , \mux_out[11][1] , \mux_out[11][0] ,
         \mux_out[10][63] , \mux_out[10][62] , \mux_out[10][61] ,
         \mux_out[10][60] , \mux_out[10][59] , \mux_out[10][58] ,
         \mux_out[10][57] , \mux_out[10][56] , \mux_out[10][55] ,
         \mux_out[10][54] , \mux_out[10][53] , \mux_out[10][52] ,
         \mux_out[10][51] , \mux_out[10][50] , \mux_out[10][49] ,
         \mux_out[10][48] , \mux_out[10][47] , \mux_out[10][46] ,
         \mux_out[10][45] , \mux_out[10][44] , \mux_out[10][43] ,
         \mux_out[10][42] , \mux_out[10][41] , \mux_out[10][40] ,
         \mux_out[10][39] , \mux_out[10][38] , \mux_out[10][37] ,
         \mux_out[10][36] , \mux_out[10][35] , \mux_out[10][34] ,
         \mux_out[10][33] , \mux_out[10][32] , \mux_out[10][31] ,
         \mux_out[10][30] , \mux_out[10][29] , \mux_out[10][28] ,
         \mux_out[10][27] , \mux_out[10][26] , \mux_out[10][25] ,
         \mux_out[10][24] , \mux_out[10][23] , \mux_out[10][22] ,
         \mux_out[10][21] , \mux_out[10][20] , \mux_out[10][19] ,
         \mux_out[10][18] , \mux_out[10][17] , \mux_out[10][16] ,
         \mux_out[10][15] , \mux_out[10][14] , \mux_out[10][13] ,
         \mux_out[10][12] , \mux_out[10][11] , \mux_out[10][10] ,
         \mux_out[10][9] , \mux_out[10][8] , \mux_out[10][7] ,
         \mux_out[10][6] , \mux_out[10][5] , \mux_out[10][4] ,
         \mux_out[10][3] , \mux_out[10][2] , \mux_out[10][1] ,
         \mux_out[10][0] , \mux_out[9][63] , \mux_out[9][62] ,
         \mux_out[9][61] , \mux_out[9][60] , \mux_out[9][59] ,
         \mux_out[9][58] , \mux_out[9][57] , \mux_out[9][56] ,
         \mux_out[9][55] , \mux_out[9][54] , \mux_out[9][53] ,
         \mux_out[9][52] , \mux_out[9][51] , \mux_out[9][50] ,
         \mux_out[9][49] , \mux_out[9][48] , \mux_out[9][47] ,
         \mux_out[9][46] , \mux_out[9][45] , \mux_out[9][44] ,
         \mux_out[9][43] , \mux_out[9][42] , \mux_out[9][41] ,
         \mux_out[9][40] , \mux_out[9][39] , \mux_out[9][38] ,
         \mux_out[9][37] , \mux_out[9][36] , \mux_out[9][35] ,
         \mux_out[9][34] , \mux_out[9][33] , \mux_out[9][32] ,
         \mux_out[9][31] , \mux_out[9][30] , \mux_out[9][29] ,
         \mux_out[9][28] , \mux_out[9][27] , \mux_out[9][26] ,
         \mux_out[9][25] , \mux_out[9][24] , \mux_out[9][23] ,
         \mux_out[9][22] , \mux_out[9][21] , \mux_out[9][20] ,
         \mux_out[9][19] , \mux_out[9][18] , \mux_out[9][17] ,
         \mux_out[9][16] , \mux_out[9][15] , \mux_out[9][14] ,
         \mux_out[9][13] , \mux_out[9][12] , \mux_out[9][11] ,
         \mux_out[9][10] , \mux_out[9][9] , \mux_out[9][8] , \mux_out[9][7] ,
         \mux_out[9][6] , \mux_out[9][5] , \mux_out[9][4] , \mux_out[9][3] ,
         \mux_out[9][2] , \mux_out[9][1] , \mux_out[9][0] , \mux_out[8][63] ,
         \mux_out[8][62] , \mux_out[8][61] , \mux_out[8][60] ,
         \mux_out[8][59] , \mux_out[8][58] , \mux_out[8][57] ,
         \mux_out[8][56] , \mux_out[8][55] , \mux_out[8][54] ,
         \mux_out[8][53] , \mux_out[8][52] , \mux_out[8][51] ,
         \mux_out[8][50] , \mux_out[8][49] , \mux_out[8][48] ,
         \mux_out[8][47] , \mux_out[8][46] , \mux_out[8][45] ,
         \mux_out[8][44] , \mux_out[8][43] , \mux_out[8][42] ,
         \mux_out[8][41] , \mux_out[8][40] , \mux_out[8][39] ,
         \mux_out[8][38] , \mux_out[8][37] , \mux_out[8][36] ,
         \mux_out[8][35] , \mux_out[8][34] , \mux_out[8][33] ,
         \mux_out[8][32] , \mux_out[8][31] , \mux_out[8][30] ,
         \mux_out[8][29] , \mux_out[8][28] , \mux_out[8][27] ,
         \mux_out[8][26] , \mux_out[8][25] , \mux_out[8][24] ,
         \mux_out[8][23] , \mux_out[8][22] , \mux_out[8][21] ,
         \mux_out[8][20] , \mux_out[8][19] , \mux_out[8][18] ,
         \mux_out[8][17] , \mux_out[8][16] , \mux_out[8][15] ,
         \mux_out[8][14] , \mux_out[8][13] , \mux_out[8][12] ,
         \mux_out[8][11] , \mux_out[8][10] , \mux_out[8][9] , \mux_out[8][8] ,
         \mux_out[8][7] , \mux_out[8][6] , \mux_out[8][5] , \mux_out[8][4] ,
         \mux_out[8][3] , \mux_out[8][2] , \mux_out[8][1] , \mux_out[8][0] ,
         \add_in[15][63] , \add_in[15][62] , \add_in[15][61] ,
         \add_in[15][60] , \add_in[15][59] , \add_in[15][58] ,
         \add_in[15][57] , \add_in[15][56] , \add_in[15][55] ,
         \add_in[15][54] , \add_in[15][53] , \add_in[15][52] ,
         \add_in[15][51] , \add_in[15][50] , \add_in[15][49] ,
         \add_in[15][48] , \add_in[15][47] , \add_in[15][46] ,
         \add_in[15][45] , \add_in[15][44] , \add_in[15][43] ,
         \add_in[15][42] , \add_in[15][41] , \add_in[15][40] ,
         \add_in[15][39] , \add_in[15][38] , \add_in[15][37] ,
         \add_in[15][36] , \add_in[15][35] , \add_in[15][34] ,
         \add_in[15][33] , \add_in[15][32] , \add_in[15][31] ,
         \add_in[15][30] , \add_in[15][29] , \add_in[15][28] ,
         \add_in[15][27] , \add_in[15][26] , \add_in[15][25] ,
         \add_in[15][24] , \add_in[15][23] , \add_in[15][22] ,
         \add_in[15][21] , \add_in[15][20] , \add_in[15][19] ,
         \add_in[15][18] , \add_in[15][17] , \add_in[15][16] ,
         \add_in[15][15] , \add_in[15][14] , \add_in[15][13] ,
         \add_in[15][12] , \add_in[15][11] , \add_in[15][10] , \add_in[15][9] ,
         \add_in[15][8] , \add_in[15][7] , \add_in[15][6] , \add_in[15][5] ,
         \add_in[15][4] , \add_in[15][3] , \add_in[15][2] , \add_in[15][1] ,
         \add_in[15][0] , \add_in[14][63] , \add_in[14][62] , \add_in[14][61] ,
         \add_in[14][60] , \add_in[14][59] , \add_in[14][58] ,
         \add_in[14][57] , \add_in[14][56] , \add_in[14][55] ,
         \add_in[14][54] , \add_in[14][53] , \add_in[14][52] ,
         \add_in[14][51] , \add_in[14][50] , \add_in[14][49] ,
         \add_in[14][48] , \add_in[14][47] , \add_in[14][46] ,
         \add_in[14][45] , \add_in[14][44] , \add_in[14][43] ,
         \add_in[14][42] , \add_in[14][41] , \add_in[14][40] ,
         \add_in[14][39] , \add_in[14][38] , \add_in[14][37] ,
         \add_in[14][36] , \add_in[14][35] , \add_in[14][34] ,
         \add_in[14][33] , \add_in[14][32] , \add_in[14][31] ,
         \add_in[14][30] , \add_in[14][29] , \add_in[14][28] ,
         \add_in[14][27] , \add_in[14][26] , \add_in[14][25] ,
         \add_in[14][24] , \add_in[14][23] , \add_in[14][22] ,
         \add_in[14][21] , \add_in[14][20] , \add_in[14][19] ,
         \add_in[14][18] , \add_in[14][17] , \add_in[14][16] ,
         \add_in[14][15] , \add_in[14][14] , \add_in[14][13] ,
         \add_in[14][12] , \add_in[14][11] , \add_in[14][10] , \add_in[14][9] ,
         \add_in[14][8] , \add_in[14][7] , \add_in[14][6] , \add_in[14][5] ,
         \add_in[14][4] , \add_in[14][3] , \add_in[14][2] , \add_in[14][1] ,
         \add_in[14][0] , \add_in[13][63] , \add_in[13][62] , \add_in[13][61] ,
         \add_in[13][60] , \add_in[13][59] , \add_in[13][58] ,
         \add_in[13][57] , \add_in[13][56] , \add_in[13][55] ,
         \add_in[13][54] , \add_in[13][53] , \add_in[13][52] ,
         \add_in[13][51] , \add_in[13][50] , \add_in[13][49] ,
         \add_in[13][48] , \add_in[13][47] , \add_in[13][46] ,
         \add_in[13][45] , \add_in[13][44] , \add_in[13][43] ,
         \add_in[13][42] , \add_in[13][41] , \add_in[13][40] ,
         \add_in[13][39] , \add_in[13][38] , \add_in[13][37] ,
         \add_in[13][36] , \add_in[13][35] , \add_in[13][34] ,
         \add_in[13][33] , \add_in[13][32] , \add_in[13][31] ,
         \add_in[13][30] , \add_in[13][29] , \add_in[13][28] ,
         \add_in[13][27] , \add_in[13][26] , \add_in[13][25] ,
         \add_in[13][24] , \add_in[13][23] , \add_in[13][22] ,
         \add_in[13][21] , \add_in[13][20] , \add_in[13][19] ,
         \add_in[13][18] , \add_in[13][17] , \add_in[13][16] ,
         \add_in[13][15] , \add_in[13][14] , \add_in[13][13] ,
         \add_in[13][12] , \add_in[13][11] , \add_in[13][10] , \add_in[13][9] ,
         \add_in[13][8] , \add_in[13][7] , \add_in[13][6] , \add_in[13][5] ,
         \add_in[13][4] , \add_in[13][3] , \add_in[13][2] , \add_in[13][1] ,
         \add_in[13][0] , \add_in[12][63] , \add_in[12][62] , \add_in[12][61] ,
         \add_in[12][60] , \add_in[12][59] , \add_in[12][58] ,
         \add_in[12][57] , \add_in[12][56] , \add_in[12][55] ,
         \add_in[12][54] , \add_in[12][53] , \add_in[12][52] ,
         \add_in[12][51] , \add_in[12][50] , \add_in[12][49] ,
         \add_in[12][48] , \add_in[12][47] , \add_in[12][46] ,
         \add_in[12][45] , \add_in[12][44] , \add_in[12][43] ,
         \add_in[12][42] , \add_in[12][41] , \add_in[12][40] ,
         \add_in[12][39] , \add_in[12][38] , \add_in[12][37] ,
         \add_in[12][36] , \add_in[12][35] , \add_in[12][34] ,
         \add_in[12][33] , \add_in[12][32] , \add_in[12][31] ,
         \add_in[12][30] , \add_in[12][29] , \add_in[12][28] ,
         \add_in[12][27] , \add_in[12][26] , \add_in[12][25] ,
         \add_in[12][24] , \add_in[12][23] , \add_in[12][22] ,
         \add_in[12][21] , \add_in[12][20] , \add_in[12][19] ,
         \add_in[12][18] , \add_in[12][17] , \add_in[12][16] ,
         \add_in[12][15] , \add_in[12][14] , \add_in[12][13] ,
         \add_in[12][12] , \add_in[12][11] , \add_in[12][10] , \add_in[12][9] ,
         \add_in[12][8] , \add_in[12][7] , \add_in[12][6] , \add_in[12][5] ,
         \add_in[12][4] , \add_in[12][3] , \add_in[12][2] , \add_in[12][1] ,
         \add_in[12][0] , \add_in[11][63] , \add_in[11][62] , \add_in[11][61] ,
         \add_in[11][60] , \add_in[11][59] , \add_in[11][58] ,
         \add_in[11][57] , \add_in[11][56] , \add_in[11][55] ,
         \add_in[11][54] , \add_in[11][53] , \add_in[11][52] ,
         \add_in[11][51] , \add_in[11][50] , \add_in[11][49] ,
         \add_in[11][48] , \add_in[11][47] , \add_in[11][46] ,
         \add_in[11][45] , \add_in[11][44] , \add_in[11][43] ,
         \add_in[11][42] , \add_in[11][41] , \add_in[11][40] ,
         \add_in[11][39] , \add_in[11][38] , \add_in[11][37] ,
         \add_in[11][36] , \add_in[11][35] , \add_in[11][34] ,
         \add_in[11][33] , \add_in[11][32] , \add_in[11][31] ,
         \add_in[11][30] , \add_in[11][29] , \add_in[11][28] ,
         \add_in[11][27] , \add_in[11][26] , \add_in[11][25] ,
         \add_in[11][24] , \add_in[11][23] , \add_in[11][22] ,
         \add_in[11][21] , \add_in[11][20] , \add_in[11][19] ,
         \add_in[11][18] , \add_in[11][17] , \add_in[11][16] ,
         \add_in[11][15] , \add_in[11][14] , \add_in[11][13] ,
         \add_in[11][12] , \add_in[11][11] , \add_in[11][10] , \add_in[11][9] ,
         \add_in[11][8] , \add_in[11][7] , \add_in[11][6] , \add_in[11][5] ,
         \add_in[11][4] , \add_in[11][3] , \add_in[11][2] , \add_in[11][1] ,
         \add_in[11][0] , \add_in[10][63] , \add_in[10][62] , \add_in[10][61] ,
         \add_in[10][60] , \add_in[10][59] , \add_in[10][58] ,
         \add_in[10][57] , \add_in[10][56] , \add_in[10][55] ,
         \add_in[10][54] , \add_in[10][53] , \add_in[10][52] ,
         \add_in[10][51] , \add_in[10][50] , \add_in[10][49] ,
         \add_in[10][48] , \add_in[10][47] , \add_in[10][46] ,
         \add_in[10][45] , \add_in[10][44] , \add_in[10][43] ,
         \add_in[10][42] , \add_in[10][41] , \add_in[10][40] ,
         \add_in[10][39] , \add_in[10][38] , \add_in[10][37] ,
         \add_in[10][36] , \add_in[10][35] , \add_in[10][34] ,
         \add_in[10][33] , \add_in[10][32] , \add_in[10][31] ,
         \add_in[10][30] , \add_in[10][29] , \add_in[10][28] ,
         \add_in[10][27] , \add_in[10][26] , \add_in[10][25] ,
         \add_in[10][24] , \add_in[10][23] , \add_in[10][22] ,
         \add_in[10][21] , \add_in[10][20] , \add_in[10][19] ,
         \add_in[10][18] , \add_in[10][17] , \add_in[10][16] ,
         \add_in[10][15] , \add_in[10][14] , \add_in[10][13] ,
         \add_in[10][12] , \add_in[10][11] , \add_in[10][10] , \add_in[10][9] ,
         \add_in[10][8] , \add_in[10][7] , \add_in[10][6] , \add_in[10][5] ,
         \add_in[10][4] , \add_in[10][3] , \add_in[10][2] , \add_in[10][1] ,
         \add_in[10][0] , \add_in[9][63] , \add_in[9][62] , \add_in[9][61] ,
         \add_in[9][60] , \add_in[9][59] , \add_in[9][58] , \add_in[9][57] ,
         \add_in[9][56] , \add_in[9][55] , \add_in[9][54] , \add_in[9][53] ,
         \add_in[9][52] , \add_in[9][51] , \add_in[9][50] , \add_in[9][49] ,
         \add_in[9][48] , \add_in[9][47] , \add_in[9][46] , \add_in[9][45] ,
         \add_in[9][44] , \add_in[9][43] , \add_in[9][42] , \add_in[9][41] ,
         \add_in[9][40] , \add_in[9][39] , \add_in[9][38] , \add_in[9][37] ,
         \add_in[9][36] , \add_in[9][35] , \add_in[9][34] , \add_in[9][33] ,
         \add_in[9][32] , \add_in[9][31] , \add_in[9][30] , \add_in[9][29] ,
         \add_in[9][28] , \add_in[9][27] , \add_in[9][26] , \add_in[9][25] ,
         \add_in[9][24] , \add_in[9][23] , \add_in[9][22] , \add_in[9][21] ,
         \add_in[9][20] , \add_in[9][19] , \add_in[9][18] , \add_in[9][17] ,
         \add_in[9][16] , \add_in[9][15] , \add_in[9][14] , \add_in[9][13] ,
         \add_in[9][12] , \add_in[9][11] , \add_in[9][10] , \add_in[9][9] ,
         \add_in[9][8] , \add_in[9][7] , \add_in[9][6] , \add_in[9][5] ,
         \add_in[9][4] , \add_in[9][3] , \add_in[9][2] , \add_in[9][1] ,
         \add_in[9][0] , \add_in[8][63] , \add_in[8][62] , \add_in[8][61] ,
         \add_in[8][60] , \add_in[8][59] , \add_in[8][58] , \add_in[8][57] ,
         \add_in[8][56] , \add_in[8][55] , \add_in[8][54] , \add_in[8][53] ,
         \add_in[8][52] , \add_in[8][51] , \add_in[8][50] , \add_in[8][49] ,
         \add_in[8][48] , \add_in[8][47] , \add_in[8][46] , \add_in[8][45] ,
         \add_in[8][44] , \add_in[8][43] , \add_in[8][42] , \add_in[8][41] ,
         \add_in[8][40] , \add_in[8][39] , \add_in[8][38] , \add_in[8][37] ,
         \add_in[8][36] , \add_in[8][35] , \add_in[8][34] , \add_in[8][33] ,
         \add_in[8][32] , \add_in[8][31] , \add_in[8][30] , \add_in[8][29] ,
         \add_in[8][28] , \add_in[8][27] , \add_in[8][26] , \add_in[8][25] ,
         \add_in[8][24] , \add_in[8][23] , \add_in[8][22] , \add_in[8][21] ,
         \add_in[8][20] , \add_in[8][19] , \add_in[8][18] , \add_in[8][17] ,
         \add_in[8][16] , \add_in[8][15] , \add_in[8][14] , \add_in[8][13] ,
         \add_in[8][12] , \add_in[8][11] , \add_in[8][10] , \add_in[8][9] ,
         \add_in[8][8] , \add_in[8][7] , \add_in[8][6] , \add_in[8][5] ,
         \add_in[8][4] , \add_in[8][3] , \add_in[8][2] , \add_in[8][1] ,
         \add_in[8][0] , \add_in[7][63] , \add_in[7][62] , \add_in[7][61] ,
         \add_in[7][60] , \add_in[7][59] , \add_in[7][58] , \add_in[7][57] ,
         \add_in[7][56] , \add_in[7][55] , \add_in[7][54] , \add_in[7][53] ,
         \add_in[7][52] , \add_in[7][51] , \add_in[7][50] , \add_in[7][49] ,
         \add_in[7][48] , \add_in[7][47] , \add_in[7][46] , \add_in[7][45] ,
         \add_in[7][44] , \add_in[7][43] , \add_in[7][42] , \add_in[7][41] ,
         \add_in[7][40] , \add_in[7][39] , \add_in[7][38] , \add_in[7][37] ,
         \add_in[7][36] , \add_in[7][35] , \add_in[7][34] , \add_in[7][33] ,
         \add_in[7][32] , \add_in[7][31] , \add_in[7][30] , \add_in[7][29] ,
         \add_in[7][28] , \add_in[7][27] , \add_in[7][26] , \add_in[7][25] ,
         \add_in[7][24] , \add_in[7][23] , \add_in[7][22] , \add_in[7][21] ,
         \add_in[7][20] , \add_in[7][19] , \add_in[7][18] , \add_in[7][17] ,
         \add_in[7][16] , \add_in[7][15] , \add_in[7][14] , \add_in[7][13] ,
         \add_in[7][12] , \add_in[7][11] , \add_in[7][10] , \add_in[7][9] ,
         \add_in[7][8] , \add_in[7][7] , \add_in[7][6] , \add_in[7][5] ,
         \add_in[7][4] , \add_in[7][3] , \add_in[7][2] , \add_in[7][1] ,
         \add_in[7][0] , \add_in[6][63] , \add_in[6][62] , \add_in[6][61] ,
         \add_in[6][60] , \add_in[6][59] , \add_in[6][58] , \add_in[6][57] ,
         \add_in[6][56] , \add_in[6][55] , \add_in[6][54] , \add_in[6][53] ,
         \add_in[6][52] , \add_in[6][51] , \add_in[6][50] , \add_in[6][49] ,
         \add_in[6][48] , \add_in[6][47] , \add_in[6][46] , \add_in[6][45] ,
         \add_in[6][44] , \add_in[6][43] , \add_in[6][42] , \add_in[6][41] ,
         \add_in[6][40] , \add_in[6][39] , \add_in[6][38] , \add_in[6][37] ,
         \add_in[6][36] , \add_in[6][35] , \add_in[6][34] , \add_in[6][33] ,
         \add_in[6][32] , \add_in[6][31] , \add_in[6][30] , \add_in[6][29] ,
         \add_in[6][28] , \add_in[6][27] , \add_in[6][26] , \add_in[6][25] ,
         \add_in[6][24] , \add_in[6][23] , \add_in[6][22] , \add_in[6][21] ,
         \add_in[6][20] , \add_in[6][19] , \add_in[6][18] , \add_in[6][17] ,
         \add_in[6][16] , \add_in[6][15] , \add_in[6][14] , \add_in[6][13] ,
         \add_in[6][12] , \add_in[6][11] , \add_in[6][10] , \add_in[6][9] ,
         \add_in[6][8] , \add_in[6][7] , \add_in[6][6] , \add_in[6][5] ,
         \add_in[6][4] , \add_in[6][3] , \add_in[6][2] , \add_in[6][1] ,
         \add_in[6][0] , \add_in[5][63] , \add_in[5][62] , \add_in[5][61] ,
         \add_in[5][60] , \add_in[5][59] , \add_in[5][58] , \add_in[5][57] ,
         \add_in[5][56] , \add_in[5][55] , \add_in[5][54] , \add_in[5][53] ,
         \add_in[5][52] , \add_in[5][51] , \add_in[5][50] , \add_in[5][49] ,
         \add_in[5][48] , \add_in[5][47] , \add_in[5][46] , \add_in[5][45] ,
         \add_in[5][44] , \add_in[5][43] , \add_in[5][42] , \add_in[5][41] ,
         \add_in[5][40] , \add_in[5][39] , \add_in[5][38] , \add_in[5][37] ,
         \add_in[5][36] , \add_in[5][35] , \add_in[5][34] , \add_in[5][33] ,
         \add_in[5][32] , \add_in[5][31] , \add_in[5][30] , \add_in[5][29] ,
         \add_in[5][28] , \add_in[5][27] , \add_in[5][26] , \add_in[5][25] ,
         \add_in[5][24] , \add_in[5][23] , \add_in[5][22] , \add_in[5][21] ,
         \add_in[5][20] , \add_in[5][19] , \add_in[5][18] , \add_in[5][17] ,
         \add_in[5][16] , \add_in[5][15] , \add_in[5][14] , \add_in[5][13] ,
         \add_in[5][12] , \add_in[5][11] , \add_in[5][10] , \add_in[5][9] ,
         \add_in[5][8] , \add_in[5][7] , \add_in[5][6] , \add_in[5][5] ,
         \add_in[5][4] , \add_in[5][3] , \add_in[5][2] , \add_in[5][1] ,
         \add_in[5][0] , \add_in[4][63] , \add_in[4][62] , \add_in[4][61] ,
         \add_in[4][60] , \add_in[4][59] , \add_in[4][58] , \add_in[4][57] ,
         \add_in[4][56] , \add_in[4][55] , \add_in[4][54] , \add_in[4][53] ,
         \add_in[4][52] , \add_in[4][51] , \add_in[4][50] , \add_in[4][49] ,
         \add_in[4][48] , \add_in[4][47] , \add_in[4][46] , \add_in[4][45] ,
         \add_in[4][44] , \add_in[4][43] , \add_in[4][42] , \add_in[4][41] ,
         \add_in[4][40] , \add_in[4][39] , \add_in[4][38] , \add_in[4][37] ,
         \add_in[4][36] , \add_in[4][35] , \add_in[4][34] , \add_in[4][33] ,
         \add_in[4][32] , \add_in[4][31] , \add_in[4][30] , \add_in[4][29] ,
         \add_in[4][28] , \add_in[4][27] , \add_in[4][26] , \add_in[4][25] ,
         \add_in[4][24] , \add_in[4][23] , \add_in[4][22] , \add_in[4][21] ,
         \add_in[4][20] , \add_in[4][19] , \add_in[4][18] , \add_in[4][17] ,
         \add_in[4][16] , \add_in[4][15] , \add_in[4][14] , \add_in[4][13] ,
         \add_in[4][12] , \add_in[4][11] , \add_in[4][10] , \add_in[4][9] ,
         \add_in[4][8] , \add_in[4][7] , \add_in[4][6] , \add_in[4][5] ,
         \add_in[4][4] , \add_in[4][3] , \add_in[4][2] , \add_in[4][1] ,
         \add_in[4][0] , \add_in[3][63] , \add_in[3][62] , \add_in[3][61] ,
         \add_in[3][60] , \add_in[3][59] , \add_in[3][58] , \add_in[3][57] ,
         \add_in[3][56] , \add_in[3][55] , \add_in[3][54] , \add_in[3][53] ,
         \add_in[3][52] , \add_in[3][51] , \add_in[3][50] , \add_in[3][49] ,
         \add_in[3][48] , \add_in[3][47] , \add_in[3][46] , \add_in[3][45] ,
         \add_in[3][44] , \add_in[3][43] , \add_in[3][42] , \add_in[3][41] ,
         \add_in[3][40] , \add_in[3][39] , \add_in[3][38] , \add_in[3][37] ,
         \add_in[3][36] , \add_in[3][35] , \add_in[3][34] , \add_in[3][33] ,
         \add_in[3][32] , \add_in[3][31] , \add_in[3][30] , \add_in[3][29] ,
         \add_in[3][28] , \add_in[3][27] , \add_in[3][26] , \add_in[3][25] ,
         \add_in[3][24] , \add_in[3][23] , \add_in[3][22] , \add_in[3][21] ,
         \add_in[3][20] , \add_in[3][19] , \add_in[3][18] , \add_in[3][17] ,
         \add_in[3][16] , \add_in[3][15] , \add_in[3][14] , \add_in[3][13] ,
         \add_in[3][12] , \add_in[3][11] , \add_in[3][10] , \add_in[3][9] ,
         \add_in[3][8] , \add_in[3][7] , \add_in[3][6] , \add_in[3][5] ,
         \add_in[3][4] , \add_in[3][3] , \add_in[3][2] , \add_in[3][1] ,
         \add_in[3][0] , \add_in[2][63] , \add_in[2][62] , \add_in[2][61] ,
         \add_in[2][60] , \add_in[2][59] , \add_in[2][58] , \add_in[2][57] ,
         \add_in[2][56] , \add_in[2][55] , \add_in[2][54] , \add_in[2][53] ,
         \add_in[2][52] , \add_in[2][51] , \add_in[2][50] , \add_in[2][49] ,
         \add_in[2][48] , \add_in[2][47] , \add_in[2][46] , \add_in[2][45] ,
         \add_in[2][44] , \add_in[2][43] , \add_in[2][42] , \add_in[2][41] ,
         \add_in[2][40] , \add_in[2][39] , \add_in[2][38] , \add_in[2][37] ,
         \add_in[2][36] , \add_in[2][35] , \add_in[2][34] , \add_in[2][33] ,
         \add_in[2][32] , \add_in[2][31] , \add_in[2][30] , \add_in[2][29] ,
         \add_in[2][28] , \add_in[2][27] , \add_in[2][26] , \add_in[2][25] ,
         \add_in[2][24] , \add_in[2][23] , \add_in[2][22] , \add_in[2][21] ,
         \add_in[2][20] , \add_in[2][19] , \add_in[2][18] , \add_in[2][17] ,
         \add_in[2][16] , \add_in[2][15] , \add_in[2][14] , \add_in[2][13] ,
         \add_in[2][12] , \add_in[2][11] , \add_in[2][10] , \add_in[2][9] ,
         \add_in[2][8] , \add_in[2][7] , \add_in[2][6] , \add_in[2][5] ,
         \add_in[2][4] , \add_in[2][3] , \add_in[2][2] , \add_in[2][1] ,
         \add_in[2][0] , \add_in[1][63] , \add_in[1][62] , \add_in[1][61] ,
         \add_in[1][60] , \add_in[1][59] , \add_in[1][58] , \add_in[1][57] ,
         \add_in[1][56] , \add_in[1][55] , \add_in[1][54] , \add_in[1][53] ,
         \add_in[1][52] , \add_in[1][51] , \add_in[1][50] , \add_in[1][49] ,
         \add_in[1][48] , \add_in[1][47] , \add_in[1][46] , \add_in[1][45] ,
         \add_in[1][44] , \add_in[1][43] , \add_in[1][42] , \add_in[1][41] ,
         \add_in[1][40] , \add_in[1][39] , \add_in[1][38] , \add_in[1][37] ,
         \add_in[1][36] , \add_in[1][35] , \add_in[1][34] , \add_in[1][33] ,
         \add_in[1][32] , \add_in[1][31] , \add_in[1][30] , \add_in[1][29] ,
         \add_in[1][28] , \add_in[1][27] , \add_in[1][26] , \add_in[1][25] ,
         \add_in[1][24] , \add_in[1][23] , \add_in[1][22] , \add_in[1][21] ,
         \add_in[1][20] , \add_in[1][19] , \add_in[1][18] , \add_in[1][17] ,
         \add_in[1][16] , \add_in[1][15] , \add_in[1][14] , \add_in[1][13] ,
         \add_in[1][12] , \add_in[1][11] , \add_in[1][10] , \add_in[1][9] ,
         \add_in[1][8] , \add_in[1][7] , \add_in[1][6] , \add_in[1][5] ,
         \add_in[1][4] , \add_in[1][3] , \add_in[1][2] , \add_in[1][1] ,
         \add_in[1][0] , \add_in[0][63] , \add_in[0][62] , \add_in[0][61] ,
         \add_in[0][60] , \add_in[0][59] , \add_in[0][58] , \add_in[0][57] ,
         \add_in[0][56] , \add_in[0][55] , \add_in[0][54] , \add_in[0][53] ,
         \add_in[0][52] , \add_in[0][51] , \add_in[0][50] , \add_in[0][49] ,
         \add_in[0][48] , \add_in[0][47] , \add_in[0][46] , \add_in[0][45] ,
         \add_in[0][44] , \add_in[0][43] , \add_in[0][42] , \add_in[0][41] ,
         \add_in[0][40] , \add_in[0][39] , \add_in[0][38] , \add_in[0][37] ,
         \add_in[0][36] , \add_in[0][35] , \add_in[0][34] , \add_in[0][33] ,
         \add_in[0][32] , \add_in[0][31] , \add_in[0][30] , \add_in[0][29] ,
         \add_in[0][28] , \add_in[0][27] , \add_in[0][26] , \add_in[0][25] ,
         \add_in[0][24] , \add_in[0][23] , \add_in[0][22] , \add_in[0][21] ,
         \add_in[0][20] , \add_in[0][19] , \add_in[0][18] , \add_in[0][17] ,
         \add_in[0][16] , \add_in[0][15] , \add_in[0][14] , \add_in[0][13] ,
         \add_in[0][12] , \add_in[0][11] , \add_in[0][10] , \add_in[0][9] ,
         \add_in[0][8] , \add_in[0][7] , \add_in[0][6] , \add_in[0][5] ,
         \add_in[0][4] , \add_in[0][3] , \add_in[0][2] , \add_in[0][1] ,
         \add_in[0][0] , n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695;
  wire   [47:0] encoder_out;
  wire   [15:0] mode;
  assign mode[0] = B[1];

  BOOTH_ENCODER_4 enc_i_0 ( .I({mode[0], B[0], 1'b0}), .O(encoder_out[2:0]) );
  BOOTH_ENCODER_19 enc_i_1 ( .I({B[3:2], mode[0]}), .O(encoder_out[5:3]) );
  BOOTH_ENCODER_18 enc_i_2 ( .I(B[5:3]), .O(encoder_out[8:6]) );
  BOOTH_ENCODER_17 enc_i_3 ( .I(B[7:5]), .O(encoder_out[11:9]) );
  BOOTH_ENCODER_16 enc_i_4 ( .I(B[9:7]), .O(encoder_out[14:12]) );
  BOOTH_ENCODER_15 enc_i_5 ( .I(B[11:9]), .O(encoder_out[17:15]) );
  BOOTH_ENCODER_14 enc_i_6 ( .I(B[13:11]), .O(encoder_out[20:18]) );
  BOOTH_ENCODER_13 enc_i_7 ( .I(B[15:13]), .O(encoder_out[23:21]) );
  BOOTH_ENCODER_12 enc_i_8 ( .I(B[17:15]), .O(encoder_out[26:24]) );
  BOOTH_ENCODER_11 enc_i_9 ( .I(B[19:17]), .O(encoder_out[29:27]) );
  BOOTH_ENCODER_10 enc_i_10 ( .I(B[21:19]), .O(encoder_out[32:30]) );
  BOOTH_ENCODER_9 enc_i_11 ( .I(B[23:21]), .O(encoder_out[35:33]) );
  BOOTH_ENCODER_8 enc_i_12 ( .I(B[25:23]), .O(encoder_out[38:36]) );
  BOOTH_ENCODER_7 enc_i_13 ( .I(B[27:25]), .O(encoder_out[41:39]) );
  BOOTH_ENCODER_6 enc_i_14 ( .I(B[29:27]), .O(encoder_out[44:42]) );
  BOOTH_ENCODER_5 enc_i_15 ( .I(B[31:29]), .O(encoder_out[47:45]) );
  MUX51_GENERIC_N64_0 mux_i_0 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n587, n587, 
        n587, n587, n587, n587, n587, n586, n586, n586, n586, n586, n586, n586, 
        n585, n585, n585, n585, n585, n585, n585, n584, n584, n584, n584, n584, 
        n584, n584, n583, n583, n583, n583, n583, n502, n492, n482, n472, n462, 
        n452, n442, n432, n422, n412, n402, n392, n382, n372, n362, n352, n342, 
        n332, n322, n312, n302, n292, n282, n272, n262, n252, n242, n232, n222, 
        n212, n202}), .C({n656, n659, n659, n659, n659, n659, n659, n658, n658, 
        n658, n658, n658, n658, n658, n658, n657, n657, n657, n657, n656, n656, 
        n656, n656, n656, n656, n654, n654, n654, n654, n654, n654, n654, n654, 
        n505, n495, n485, n475, n465, n455, n445, n435, n425, n415, n405, n395, 
        n385, n375, n365, n355, n345, n335, n325, n315, n305, n295, n285, n275, 
        n265, n255, n245, n235, n225, n215, n205}), .D({n583, n583, n582, n582, 
        n582, n582, n582, n582, n582, n581, n581, n581, n581, n581, n581, n581, 
        n580, n580, n580, n580, n580, n580, n580, n579, n579, n579, n579, n579, 
        n579, n579, n578, n578, n502, n492, n482, n472, n462, n452, n442, n432, 
        n422, n412, n402, n392, n382, n372, n362, n352, n342, n332, n322, n312, 
        n302, n292, n282, n272, n262, n252, n242, n232, n222, n212, n202, 1'b0}), .E({n666, n666, n666, n665, n665, n665, n665, n665, n665, n665, n665, n664, 
        n664, n664, n664, n664, n663, n663, n663, n663, n662, n662, n662, n662, 
        n662, n662, n662, n662, n662, n662, n662, n661, n506, n496, n486, n476, 
        n466, n456, n446, n436, n426, n416, n406, n396, n386, n376, n366, n356, 
        n346, n336, n326, n316, n306, n296, n286, n276, n266, n256, n246, n236, 
        n226, n216, n206, 1'b1}), .SEL(encoder_out[2:0]), .Y({\add_in[0][63] , 
        \add_in[0][62] , \add_in[0][61] , \add_in[0][60] , \add_in[0][59] , 
        \add_in[0][58] , \add_in[0][57] , \add_in[0][56] , \add_in[0][55] , 
        \add_in[0][54] , \add_in[0][53] , \add_in[0][52] , \add_in[0][51] , 
        \add_in[0][50] , \add_in[0][49] , \add_in[0][48] , \add_in[0][47] , 
        \add_in[0][46] , \add_in[0][45] , \add_in[0][44] , \add_in[0][43] , 
        \add_in[0][42] , \add_in[0][41] , \add_in[0][40] , \add_in[0][39] , 
        \add_in[0][38] , \add_in[0][37] , \add_in[0][36] , \add_in[0][35] , 
        \add_in[0][34] , \add_in[0][33] , \add_in[0][32] , \add_in[0][31] , 
        \add_in[0][30] , \add_in[0][29] , \add_in[0][28] , \add_in[0][27] , 
        \add_in[0][26] , \add_in[0][25] , \add_in[0][24] , \add_in[0][23] , 
        \add_in[0][22] , \add_in[0][21] , \add_in[0][20] , \add_in[0][19] , 
        \add_in[0][18] , \add_in[0][17] , \add_in[0][16] , \add_in[0][15] , 
        \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , \add_in[0][11] , 
        \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , \add_in[0][7] , 
        \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , \add_in[0][3] , 
        \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }) );
  MUX51_GENERIC_N64_15 mux_i_1 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n516, n516, 
        n516, n516, n516, n515, n515, n515, n515, n515, n515, n515, n514, n514, 
        n514, n514, n514, n514, n514, n513, n513, n513, n513, n513, n513, n513, 
        n512, n512, n512, n512, n512, n498, n488, n478, n468, n458, n448, n438, 
        n428, n418, n408, n398, n388, n378, n368, n358, n348, n338, n328, n318, 
        n308, n298, n288, n278, n268, n258, n248, n238, n228, n218, n208, n198, 
        1'b0, 1'b0}), .C({n653, n653, n653, n653, n653, n653, n653, n653, n653, 
        n655, n655, n655, n655, n655, n658, n658, n658, n658, n657, n657, n657, 
        n657, n657, n657, n657, n657, n656, n656, n656, n656, n656, n505, n495, 
        n485, n475, n465, n455, n445, n435, n425, n415, n405, n395, n385, n375, 
        n365, n355, n345, n335, n325, n315, n305, n295, n285, n275, n265, n255, 
        n245, n235, n225, n215, n205, 1'b1, 1'b1}), .D({n512, n512, n511, n511, 
        n511, n511, n511, n511, n511, n510, n510, n510, n510, n510, n510, n510, 
        n509, n509, n509, n509, n509, n509, n509, n508, n508, n508, n508, n508, 
        n508, n508, n498, n488, n478, n468, n458, n448, n438, n428, n418, n408, 
        n398, n388, n378, n368, n358, n348, n338, n328, n318, n308, n298, n288, 
        n278, n268, n258, n248, n238, n228, n218, n208, n198, 1'b0, 1'b0, 1'b0}), .E({n680, n680, n680, n680, n678, n678, n678, n678, n678, n678, n678, n678, 
        n678, n678, n677, n677, n677, n677, n677, n677, n677, n677, n677, n677, 
        n677, n675, n675, n674, n674, n674, n507, n497, n487, n477, n467, n457, 
        n447, n437, n427, n417, n407, n397, n387, n377, n367, n357, n347, n337, 
        n327, n317, n307, n297, n287, n277, n267, n257, n247, n237, n227, n217, 
        n207, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[5:3]), .Y({\mux_out[1][63] , 
        \mux_out[1][62] , \mux_out[1][61] , \mux_out[1][60] , \mux_out[1][59] , 
        \mux_out[1][58] , \mux_out[1][57] , \mux_out[1][56] , \mux_out[1][55] , 
        \mux_out[1][54] , \mux_out[1][53] , \mux_out[1][52] , \mux_out[1][51] , 
        \mux_out[1][50] , \mux_out[1][49] , \mux_out[1][48] , \mux_out[1][47] , 
        \mux_out[1][46] , \mux_out[1][45] , \mux_out[1][44] , \mux_out[1][43] , 
        \mux_out[1][42] , \mux_out[1][41] , \mux_out[1][40] , \mux_out[1][39] , 
        \mux_out[1][38] , \mux_out[1][37] , \mux_out[1][36] , \mux_out[1][35] , 
        \mux_out[1][34] , \mux_out[1][33] , \mux_out[1][32] , \mux_out[1][31] , 
        \mux_out[1][30] , \mux_out[1][29] , \mux_out[1][28] , \mux_out[1][27] , 
        \mux_out[1][26] , \mux_out[1][25] , \mux_out[1][24] , \mux_out[1][23] , 
        \mux_out[1][22] , \mux_out[1][21] , \mux_out[1][20] , \mux_out[1][19] , 
        \mux_out[1][18] , \mux_out[1][17] , \mux_out[1][16] , \mux_out[1][15] , 
        \mux_out[1][14] , \mux_out[1][13] , \mux_out[1][12] , \mux_out[1][11] , 
        \mux_out[1][10] , \mux_out[1][9] , \mux_out[1][8] , \mux_out[1][7] , 
        \mux_out[1][6] , \mux_out[1][5] , \mux_out[1][4] , \mux_out[1][3] , 
        \mux_out[1][2] , \mux_out[1][1] , \mux_out[1][0] }) );
  MUX51_GENERIC_N64_14 mux_i_2 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n524, n524, 
        n524, n524, n524, n524, n523, n523, n523, n523, n523, n523, n523, n522, 
        n522, n522, n522, n522, n522, n522, n521, n521, n521, n521, n521, n521, 
        n521, n520, n520, n498, n488, n478, n468, n458, n448, n438, n428, n418, 
        n408, n398, n388, n378, n368, n358, n348, n338, n328, n318, n308, n298, 
        n288, n278, n268, n258, n248, n238, n228, n218, n208, n198, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n651, n651, n651, n652, n652, n652, n652, n652, n652, 
        n652, n652, n652, n652, n652, n652, n653, n653, n653, n654, n654, n654, 
        n654, n655, n655, n655, n655, n655, n655, n655, n505, n495, n485, n475, 
        n465, n455, n445, n435, n425, n415, n405, n395, n385, n375, n365, n355, 
        n345, n335, n325, n315, n305, n295, n285, n275, n265, n255, n245, n235, 
        n225, n215, n205, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n520, n520, n520, n520, 
        n520, n519, n519, n519, n519, n519, n519, n519, n518, n518, n518, n518, 
        n518, n518, n518, n517, n517, n517, n517, n517, n517, n517, n516, n516, 
        n498, n488, n478, n468, n458, n448, n438, n428, n418, n408, n398, n388, 
        n378, n368, n358, n348, n338, n328, n318, n308, n298, n288, n278, n268, 
        n258, n248, n238, n228, n218, n208, n198, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n668, n668, n647, n667, n666, n650, n649, n648, n651, n672, n672, n672, 
        n672, n672, n670, n670, n670, n670, n670, n669, n669, n669, n669, n669, 
        n669, n669, n675, n660, n507, n497, n487, n477, n467, n457, n447, n437, 
        n427, n417, n407, n397, n387, n377, n367, n357, n347, n337, n327, n317, 
        n307, n297, n287, n277, n267, n257, n247, n237, n227, n217, n207, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[8:6]), .Y({\mux_out[2][63] , 
        \mux_out[2][62] , \mux_out[2][61] , \mux_out[2][60] , \mux_out[2][59] , 
        \mux_out[2][58] , \mux_out[2][57] , \mux_out[2][56] , \mux_out[2][55] , 
        \mux_out[2][54] , \mux_out[2][53] , \mux_out[2][52] , \mux_out[2][51] , 
        \mux_out[2][50] , \mux_out[2][49] , \mux_out[2][48] , \mux_out[2][47] , 
        \mux_out[2][46] , \mux_out[2][45] , \mux_out[2][44] , \mux_out[2][43] , 
        \mux_out[2][42] , \mux_out[2][41] , \mux_out[2][40] , \mux_out[2][39] , 
        \mux_out[2][38] , \mux_out[2][37] , \mux_out[2][36] , \mux_out[2][35] , 
        \mux_out[2][34] , \mux_out[2][33] , \mux_out[2][32] , \mux_out[2][31] , 
        \mux_out[2][30] , \mux_out[2][29] , \mux_out[2][28] , \mux_out[2][27] , 
        \mux_out[2][26] , \mux_out[2][25] , \mux_out[2][24] , \mux_out[2][23] , 
        \mux_out[2][22] , \mux_out[2][21] , \mux_out[2][20] , \mux_out[2][19] , 
        \mux_out[2][18] , \mux_out[2][17] , \mux_out[2][16] , \mux_out[2][15] , 
        \mux_out[2][14] , \mux_out[2][13] , \mux_out[2][12] , \mux_out[2][11] , 
        \mux_out[2][10] , \mux_out[2][9] , \mux_out[2][8] , \mux_out[2][7] , 
        \mux_out[2][6] , \mux_out[2][5] , \mux_out[2][4] , \mux_out[2][3] , 
        \mux_out[2][2] , \mux_out[2][1] , \mux_out[2][0] }) );
  MUX51_GENERIC_N64_13 mux_i_3 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n532, n532, 
        n532, n531, n531, n531, n531, n531, n531, n531, n530, n530, n530, n530, 
        n530, n530, n530, n529, n529, n529, n529, n529, n529, n529, n528, n528, 
        n528, n498, n488, n478, n468, n458, n448, n438, n428, n418, n408, n398, 
        n388, n378, n368, n358, n348, n338, n328, n318, n308, n298, n288, n278, 
        n268, n258, n248, n238, n228, n218, n208, n198, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n659, n659, n659, n659, n659, n659, n643, n636, n636, 
        n636, n636, n636, n636, n636, n636, n636, n636, n636, n637, n637, n637, 
        n637, n637, n637, n637, n637, n637, n505, n495, n485, n475, n465, n455, 
        n445, n435, n425, n415, n405, n395, n385, n375, n365, n355, n345, n335, 
        n325, n315, n305, n295, n285, n275, n265, n255, n245, n235, n225, n215, 
        n205, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n528, n528, n528, n528, 
        n527, n527, n527, n527, n527, n527, n527, n526, n526, n526, n526, n526, 
        n526, n526, n525, n525, n525, n525, n525, n525, n525, n524, n498, n488, 
        n478, n468, n458, n448, n438, n428, n418, n408, n398, n388, n378, n368, 
        n358, n348, n338, n328, n318, n308, n298, n288, n278, n268, n258, n248, 
        n238, n228, n218, n208, n198, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n670, n670, n670, n670, n670, n670, n670, n671, n671, n671, n671, n671, 
        n671, n671, n671, n671, n671, n671, n671, n672, n672, n672, n672, n672, 
        n672, n672, n507, n497, n487, n477, n467, n457, n447, n437, n427, n417, 
        n407, n397, n387, n377, n367, n357, n347, n337, n327, n317, n307, n297, 
        n287, n277, n267, n257, n247, n237, n227, n217, n207, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[11:9]), .Y({
        \mux_out[3][63] , \mux_out[3][62] , \mux_out[3][61] , \mux_out[3][60] , 
        \mux_out[3][59] , \mux_out[3][58] , \mux_out[3][57] , \mux_out[3][56] , 
        \mux_out[3][55] , \mux_out[3][54] , \mux_out[3][53] , \mux_out[3][52] , 
        \mux_out[3][51] , \mux_out[3][50] , \mux_out[3][49] , \mux_out[3][48] , 
        \mux_out[3][47] , \mux_out[3][46] , \mux_out[3][45] , \mux_out[3][44] , 
        \mux_out[3][43] , \mux_out[3][42] , \mux_out[3][41] , \mux_out[3][40] , 
        \mux_out[3][39] , \mux_out[3][38] , \mux_out[3][37] , \mux_out[3][36] , 
        \mux_out[3][35] , \mux_out[3][34] , \mux_out[3][33] , \mux_out[3][32] , 
        \mux_out[3][31] , \mux_out[3][30] , \mux_out[3][29] , \mux_out[3][28] , 
        \mux_out[3][27] , \mux_out[3][26] , \mux_out[3][25] , \mux_out[3][24] , 
        \mux_out[3][23] , \mux_out[3][22] , \mux_out[3][21] , \mux_out[3][20] , 
        \mux_out[3][19] , \mux_out[3][18] , \mux_out[3][17] , \mux_out[3][16] , 
        \mux_out[3][15] , \mux_out[3][14] , \mux_out[3][13] , \mux_out[3][12] , 
        \mux_out[3][11] , \mux_out[3][10] , \mux_out[3][9] , \mux_out[3][8] , 
        \mux_out[3][7] , \mux_out[3][6] , \mux_out[3][5] , \mux_out[3][4] , 
        \mux_out[3][3] , \mux_out[3][2] , \mux_out[3][1] , \mux_out[3][0] })
         );
  MUX51_GENERIC_N64_12 mux_i_4 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n539, n539, 
        n539, n538, n538, n538, n538, n538, n538, n538, n537, n537, n537, n537, 
        n537, n537, n537, n536, n536, n536, n536, n536, n536, n536, n535, n499, 
        n489, n479, n469, n459, n449, n439, n429, n419, n409, n399, n389, n379, 
        n369, n359, n349, n339, n329, n319, n309, n299, n289, n279, n269, n259, 
        n249, n239, n229, n219, n209, n199, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n637, n637, n637, n638, n638, n638, n638, n638, n638, 
        n638, n638, n638, n638, n638, n638, n639, n639, n639, n639, n639, n639, 
        n639, n639, n639, n639, n505, n495, n485, n475, n465, n455, n445, n435, 
        n425, n415, n405, n395, n385, n375, n365, n355, n345, n335, n325, n315, 
        n305, n295, n285, n275, n265, n255, n245, n235, n225, n215, n205, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n535, n535, n535, n535, 
        n535, n535, n534, n534, n534, n534, n534, n534, n534, n533, n533, n533, 
        n533, n533, n533, n533, n532, n532, n532, n532, n498, n488, n478, n468, 
        n458, n448, n438, n428, n418, n408, n398, n388, n378, n368, n358, n348, 
        n338, n328, n318, n308, n298, n288, n278, n268, n258, n248, n238, n228, 
        n218, n208, n198, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n668, n668, n668, n673, n673, n673, n673, n673, n673, n673, n673, n673, 
        n673, n673, n673, n674, n674, n674, n674, n674, n674, n674, n674, n674, 
        n507, n497, n487, n477, n467, n457, n447, n437, n427, n417, n407, n397, 
        n387, n377, n367, n357, n347, n337, n327, n317, n307, n297, n287, n277, 
        n267, n257, n247, n237, n227, n217, n207, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[14:12]), .Y({
        \mux_out[4][63] , \mux_out[4][62] , \mux_out[4][61] , \mux_out[4][60] , 
        \mux_out[4][59] , \mux_out[4][58] , \mux_out[4][57] , \mux_out[4][56] , 
        \mux_out[4][55] , \mux_out[4][54] , \mux_out[4][53] , \mux_out[4][52] , 
        \mux_out[4][51] , \mux_out[4][50] , \mux_out[4][49] , \mux_out[4][48] , 
        \mux_out[4][47] , \mux_out[4][46] , \mux_out[4][45] , \mux_out[4][44] , 
        \mux_out[4][43] , \mux_out[4][42] , \mux_out[4][41] , \mux_out[4][40] , 
        \mux_out[4][39] , \mux_out[4][38] , \mux_out[4][37] , \mux_out[4][36] , 
        \mux_out[4][35] , \mux_out[4][34] , \mux_out[4][33] , \mux_out[4][32] , 
        \mux_out[4][31] , \mux_out[4][30] , \mux_out[4][29] , \mux_out[4][28] , 
        \mux_out[4][27] , \mux_out[4][26] , \mux_out[4][25] , \mux_out[4][24] , 
        \mux_out[4][23] , \mux_out[4][22] , \mux_out[4][21] , \mux_out[4][20] , 
        \mux_out[4][19] , \mux_out[4][18] , \mux_out[4][17] , \mux_out[4][16] , 
        \mux_out[4][15] , \mux_out[4][14] , \mux_out[4][13] , \mux_out[4][12] , 
        \mux_out[4][11] , \mux_out[4][10] , \mux_out[4][9] , \mux_out[4][8] , 
        \mux_out[4][7] , \mux_out[4][6] , \mux_out[4][5] , \mux_out[4][4] , 
        \mux_out[4][3] , \mux_out[4][2] , \mux_out[4][1] , \mux_out[4][0] })
         );
  MUX51_GENERIC_N64_11 mux_i_5 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n545, n545, 
        n545, n545, n545, n545, n544, n544, n544, n544, n544, n544, n544, n543, 
        n543, n543, n543, n543, n543, n543, n542, n542, n542, n499, n489, n479, 
        n469, n459, n449, n439, n429, n419, n409, n399, n389, n379, n369, n359, 
        n349, n339, n329, n319, n309, n299, n289, n279, n269, n259, n249, n239, 
        n229, n219, n209, n199, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n639, n639, n640, n640, n640, n640, n640, n640, n640, 
        n640, n640, n640, n640, n640, n641, n641, n641, n641, n641, n641, n641, 
        n641, n641, n505, n495, n485, n475, n465, n455, n445, n435, n425, n415, 
        n405, n395, n385, n375, n365, n355, n345, n335, n325, n315, n305, n295, 
        n285, n275, n265, n255, n245, n235, n225, n215, n205, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n542, n542, n542, n542, 
        n541, n541, n541, n541, n541, n541, n541, n540, n540, n540, n540, n540, 
        n540, n540, n539, n539, n539, n539, n499, n489, n479, n469, n459, n449, 
        n439, n429, n419, n409, n399, n389, n379, n369, n359, n349, n339, n329, 
        n319, n309, n299, n289, n279, n269, n259, n249, n239, n229, n219, n209, 
        n199, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n675, n675, n675, n675, n675, n675, n675, n675, n675, n676, n676, n676, 
        n676, n676, n676, n676, n676, n676, n676, n676, n676, n677, n507, n497, 
        n487, n477, n467, n457, n447, n437, n427, n417, n407, n397, n387, n377, 
        n367, n357, n347, n337, n327, n317, n307, n297, n287, n277, n267, n257, 
        n247, n237, n227, n217, n207, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[17:15]), .Y({
        \mux_out[5][63] , \mux_out[5][62] , \mux_out[5][61] , \mux_out[5][60] , 
        \mux_out[5][59] , \mux_out[5][58] , \mux_out[5][57] , \mux_out[5][56] , 
        \mux_out[5][55] , \mux_out[5][54] , \mux_out[5][53] , \mux_out[5][52] , 
        \mux_out[5][51] , \mux_out[5][50] , \mux_out[5][49] , \mux_out[5][48] , 
        \mux_out[5][47] , \mux_out[5][46] , \mux_out[5][45] , \mux_out[5][44] , 
        \mux_out[5][43] , \mux_out[5][42] , \mux_out[5][41] , \mux_out[5][40] , 
        \mux_out[5][39] , \mux_out[5][38] , \mux_out[5][37] , \mux_out[5][36] , 
        \mux_out[5][35] , \mux_out[5][34] , \mux_out[5][33] , \mux_out[5][32] , 
        \mux_out[5][31] , \mux_out[5][30] , \mux_out[5][29] , \mux_out[5][28] , 
        \mux_out[5][27] , \mux_out[5][26] , \mux_out[5][25] , \mux_out[5][24] , 
        \mux_out[5][23] , \mux_out[5][22] , \mux_out[5][21] , \mux_out[5][20] , 
        \mux_out[5][19] , \mux_out[5][18] , \mux_out[5][17] , \mux_out[5][16] , 
        \mux_out[5][15] , \mux_out[5][14] , \mux_out[5][13] , \mux_out[5][12] , 
        \mux_out[5][11] , \mux_out[5][10] , \mux_out[5][9] , \mux_out[5][8] , 
        \mux_out[5][7] , \mux_out[5][6] , \mux_out[5][5] , \mux_out[5][4] , 
        \mux_out[5][3] , \mux_out[5][2] , \mux_out[5][1] , \mux_out[5][0] })
         );
  MUX51_GENERIC_N64_10 mux_i_6 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n551, n551, 
        n551, n551, n551, n550, n550, n550, n550, n550, n550, n550, n549, n549, 
        n549, n549, n549, n549, n549, n548, n548, n499, n489, n479, n469, n459, 
        n449, n439, n429, n419, n409, n399, n389, n379, n369, n359, n349, n339, 
        n329, n319, n309, n299, n289, n279, n269, n259, n249, n239, n229, n219, 
        n209, n199, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n641, n641, n641, n642, n642, n642, n642, n642, n642, 
        n642, n642, n642, n642, n642, n642, n643, n643, n643, n643, n643, n643, 
        n505, n495, n485, n475, n465, n455, n445, n435, n425, n415, n405, n395, 
        n385, n375, n365, n355, n345, n335, n325, n315, n305, n295, n285, n275, 
        n265, n255, n245, n235, n225, n215, n205, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n548, n548, n548, n548, 
        n548, n547, n547, n547, n547, n547, n547, n547, n546, n546, n546, n546, 
        n546, n546, n546, n545, n499, n489, n479, n469, n459, n449, n439, n429, 
        n419, n409, n399, n389, n379, n369, n359, n349, n339, n329, n319, n309, 
        n299, n289, n279, n269, n259, n249, n239, n229, n219, n209, n199, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n678, n678, n679, n679, n679, n679, n679, n679, n679, n679, n679, n679, 
        n679, n679, n680, n680, n680, n680, n680, n680, n507, n497, n487, n477, 
        n467, n457, n447, n437, n427, n417, n407, n397, n387, n377, n367, n357, 
        n347, n337, n327, n317, n307, n297, n287, n277, n267, n257, n247, n237, 
        n227, n217, n207, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[20:18]), .Y({
        \mux_out[6][63] , \mux_out[6][62] , \mux_out[6][61] , \mux_out[6][60] , 
        \mux_out[6][59] , \mux_out[6][58] , \mux_out[6][57] , \mux_out[6][56] , 
        \mux_out[6][55] , \mux_out[6][54] , \mux_out[6][53] , \mux_out[6][52] , 
        \mux_out[6][51] , \mux_out[6][50] , \mux_out[6][49] , \mux_out[6][48] , 
        \mux_out[6][47] , \mux_out[6][46] , \mux_out[6][45] , \mux_out[6][44] , 
        \mux_out[6][43] , \mux_out[6][42] , \mux_out[6][41] , \mux_out[6][40] , 
        \mux_out[6][39] , \mux_out[6][38] , \mux_out[6][37] , \mux_out[6][36] , 
        \mux_out[6][35] , \mux_out[6][34] , \mux_out[6][33] , \mux_out[6][32] , 
        \mux_out[6][31] , \mux_out[6][30] , \mux_out[6][29] , \mux_out[6][28] , 
        \mux_out[6][27] , \mux_out[6][26] , \mux_out[6][25] , \mux_out[6][24] , 
        \mux_out[6][23] , \mux_out[6][22] , \mux_out[6][21] , \mux_out[6][20] , 
        \mux_out[6][19] , \mux_out[6][18] , \mux_out[6][17] , \mux_out[6][16] , 
        \mux_out[6][15] , \mux_out[6][14] , \mux_out[6][13] , \mux_out[6][12] , 
        \mux_out[6][11] , \mux_out[6][10] , \mux_out[6][9] , \mux_out[6][8] , 
        \mux_out[6][7] , \mux_out[6][6] , \mux_out[6][5] , \mux_out[6][4] , 
        \mux_out[6][3] , \mux_out[6][2] , \mux_out[6][1] , \mux_out[6][0] })
         );
  MUX51_GENERIC_N64_9 mux_i_7 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n556, n556, 
        n556, n556, n556, n556, n556, n555, n555, n555, n555, n555, n555, n555, 
        n554, n554, n554, n554, n554, n499, n489, n479, n469, n459, n449, n439, 
        n429, n419, n409, n399, n389, n379, n369, n359, n349, n339, n329, n319, 
        n309, n299, n289, n279, n269, n259, n249, n239, n229, n219, n209, n199, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n643, n643, n643, n643, n643, n644, n644, n644, n644, 
        n644, n644, n644, n644, n644, n644, n644, n644, n645, n645, n505, n495, 
        n485, n475, n465, n455, n445, n435, n425, n415, n405, n395, n385, n375, 
        n365, n355, n345, n335, n325, n315, n305, n295, n285, n275, n265, n255, 
        n245, n235, n225, n215, n205, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n554, n554, n553, n553, 
        n553, n553, n553, n553, n553, n552, n552, n552, n552, n552, n552, n552, 
        n551, n551, n499, n489, n479, n469, n459, n449, n439, n429, n419, n409, 
        n399, n389, n379, n369, n359, n349, n339, n329, n319, n309, n299, n289, 
        n279, n269, n259, n249, n239, n229, n219, n209, n199, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n680, n680, n668, n668, n668, n668, n668, n668, n668, n650, n663, n660, 
        n661, n660, n660, n661, n660, n660, n507, n497, n487, n477, n467, n457, 
        n447, n437, n427, n417, n407, n397, n387, n377, n367, n357, n347, n337, 
        n327, n317, n307, n297, n287, n277, n267, n257, n247, n237, n227, n217, 
        n207, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[23:21]), .Y({
        \mux_out[7][63] , \mux_out[7][62] , \mux_out[7][61] , \mux_out[7][60] , 
        \mux_out[7][59] , \mux_out[7][58] , \mux_out[7][57] , \mux_out[7][56] , 
        \mux_out[7][55] , \mux_out[7][54] , \mux_out[7][53] , \mux_out[7][52] , 
        \mux_out[7][51] , \mux_out[7][50] , \mux_out[7][49] , \mux_out[7][48] , 
        \mux_out[7][47] , \mux_out[7][46] , \mux_out[7][45] , \mux_out[7][44] , 
        \mux_out[7][43] , \mux_out[7][42] , \mux_out[7][41] , \mux_out[7][40] , 
        \mux_out[7][39] , \mux_out[7][38] , \mux_out[7][37] , \mux_out[7][36] , 
        \mux_out[7][35] , \mux_out[7][34] , \mux_out[7][33] , \mux_out[7][32] , 
        \mux_out[7][31] , \mux_out[7][30] , \mux_out[7][29] , \mux_out[7][28] , 
        \mux_out[7][27] , \mux_out[7][26] , \mux_out[7][25] , \mux_out[7][24] , 
        \mux_out[7][23] , \mux_out[7][22] , \mux_out[7][21] , \mux_out[7][20] , 
        \mux_out[7][19] , \mux_out[7][18] , \mux_out[7][17] , \mux_out[7][16] , 
        \mux_out[7][15] , \mux_out[7][14] , \mux_out[7][13] , \mux_out[7][12] , 
        \mux_out[7][11] , \mux_out[7][10] , \mux_out[7][9] , \mux_out[7][8] , 
        \mux_out[7][7] , \mux_out[7][6] , \mux_out[7][5] , \mux_out[7][4] , 
        \mux_out[7][3] , \mux_out[7][2] , \mux_out[7][1] , \mux_out[7][0] })
         );
  MUX51_GENERIC_N64_8 mux_i_8 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n561, n561, 
        n561, n561, n561, n560, n560, n560, n560, n560, n560, n560, n559, n559, 
        n559, n559, n559, n500, n490, n480, n470, n460, n450, n440, n430, n420, 
        n410, n400, n390, n380, n370, n360, n350, n340, n330, n320, n310, n300, 
        n290, n280, n270, n260, n250, n240, n230, n220, n210, n200, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n645, n645, n645, n645, n645, n645, n645, n645, n645, 
        n645, n646, n646, n646, n646, n646, n646, n646, n506, n496, n486, n476, 
        n466, n456, n446, n436, n426, n416, n406, n396, n386, n376, n366, n356, 
        n346, n336, n326, n316, n306, n296, n286, n276, n266, n256, n246, n236, 
        n226, n216, n206, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n559, n559, n558, n558, 
        n558, n558, n558, n558, n558, n557, n557, n557, n557, n557, n557, n557, 
        n500, n490, n480, n470, n460, n450, n440, n430, n420, n410, n400, n390, 
        n380, n370, n360, n350, n340, n330, n320, n310, n300, n290, n280, n270, 
        n260, n250, n240, n230, n220, n210, n200, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n660, n660, n660, n660, n660, n660, n661, n661, n661, n661, n661, n661, 
        n661, n661, n661, n662, n507, n497, n487, n477, n467, n457, n447, n437, 
        n427, n417, n407, n397, n387, n377, n367, n357, n347, n337, n327, n317, 
        n307, n297, n287, n277, n267, n257, n247, n237, n227, n217, n207, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[26:24]), .Y({
        \mux_out[8][63] , \mux_out[8][62] , \mux_out[8][61] , \mux_out[8][60] , 
        \mux_out[8][59] , \mux_out[8][58] , \mux_out[8][57] , \mux_out[8][56] , 
        \mux_out[8][55] , \mux_out[8][54] , \mux_out[8][53] , \mux_out[8][52] , 
        \mux_out[8][51] , \mux_out[8][50] , \mux_out[8][49] , \mux_out[8][48] , 
        \mux_out[8][47] , \mux_out[8][46] , \mux_out[8][45] , \mux_out[8][44] , 
        \mux_out[8][43] , \mux_out[8][42] , \mux_out[8][41] , \mux_out[8][40] , 
        \mux_out[8][39] , \mux_out[8][38] , \mux_out[8][37] , \mux_out[8][36] , 
        \mux_out[8][35] , \mux_out[8][34] , \mux_out[8][33] , \mux_out[8][32] , 
        \mux_out[8][31] , \mux_out[8][30] , \mux_out[8][29] , \mux_out[8][28] , 
        \mux_out[8][27] , \mux_out[8][26] , \mux_out[8][25] , \mux_out[8][24] , 
        \mux_out[8][23] , \mux_out[8][22] , \mux_out[8][21] , \mux_out[8][20] , 
        \mux_out[8][19] , \mux_out[8][18] , \mux_out[8][17] , \mux_out[8][16] , 
        \mux_out[8][15] , \mux_out[8][14] , \mux_out[8][13] , \mux_out[8][12] , 
        \mux_out[8][11] , \mux_out[8][10] , \mux_out[8][9] , \mux_out[8][8] , 
        \mux_out[8][7] , \mux_out[8][6] , \mux_out[8][5] , \mux_out[8][4] , 
        \mux_out[8][3] , \mux_out[8][2] , \mux_out[8][1] , \mux_out[8][0] })
         );
  MUX51_GENERIC_N64_7 mux_i_9 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n565, n565, 
        n565, n565, n565, n565, n564, n564, n564, n564, n564, n564, n564, n563, 
        n563, n500, n490, n480, n470, n460, n450, n440, n430, n420, n410, n400, 
        n390, n380, n370, n360, n350, n340, n330, n320, n310, n300, n290, n280, 
        n270, n260, n250, n240, n230, n220, n210, n200, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n646, n646, n646, n646, n646, n647, n647, n647, n647, 
        n647, n647, n647, n647, n647, n647, n506, n496, n486, n476, n466, n456, 
        n446, n436, n426, n416, n406, n396, n386, n376, n366, n356, n346, n336, 
        n326, n316, n306, n296, n286, n276, n266, n256, n246, n236, n226, n216, 
        n206, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n563, n563, n563, n563, 
        n563, n562, n562, n562, n562, n562, n562, n562, n561, n561, n500, n490, 
        n480, n470, n460, n450, n440, n430, n420, n410, n400, n390, n380, n370, 
        n360, n350, n340, n330, n320, n310, n300, n290, n280, n270, n260, n250, 
        n240, n230, n220, n210, n200, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n663, n663, n663, n663, n663, n663, n663, n664, n664, n664, n664, n664, 
        n664, n664, n506, n496, n486, n476, n466, n456, n446, n436, n426, n416, 
        n406, n396, n386, n376, n366, n356, n346, n336, n326, n316, n306, n296, 
        n286, n276, n266, n256, n246, n236, n226, n216, n206, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[29:27]), .Y({
        \mux_out[9][63] , \mux_out[9][62] , \mux_out[9][61] , \mux_out[9][60] , 
        \mux_out[9][59] , \mux_out[9][58] , \mux_out[9][57] , \mux_out[9][56] , 
        \mux_out[9][55] , \mux_out[9][54] , \mux_out[9][53] , \mux_out[9][52] , 
        \mux_out[9][51] , \mux_out[9][50] , \mux_out[9][49] , \mux_out[9][48] , 
        \mux_out[9][47] , \mux_out[9][46] , \mux_out[9][45] , \mux_out[9][44] , 
        \mux_out[9][43] , \mux_out[9][42] , \mux_out[9][41] , \mux_out[9][40] , 
        \mux_out[9][39] , \mux_out[9][38] , \mux_out[9][37] , \mux_out[9][36] , 
        \mux_out[9][35] , \mux_out[9][34] , \mux_out[9][33] , \mux_out[9][32] , 
        \mux_out[9][31] , \mux_out[9][30] , \mux_out[9][29] , \mux_out[9][28] , 
        \mux_out[9][27] , \mux_out[9][26] , \mux_out[9][25] , \mux_out[9][24] , 
        \mux_out[9][23] , \mux_out[9][22] , \mux_out[9][21] , \mux_out[9][20] , 
        \mux_out[9][19] , \mux_out[9][18] , \mux_out[9][17] , \mux_out[9][16] , 
        \mux_out[9][15] , \mux_out[9][14] , \mux_out[9][13] , \mux_out[9][12] , 
        \mux_out[9][11] , \mux_out[9][10] , \mux_out[9][9] , \mux_out[9][8] , 
        \mux_out[9][7] , \mux_out[9][6] , \mux_out[9][5] , \mux_out[9][4] , 
        \mux_out[9][3] , \mux_out[9][2] , \mux_out[9][1] , \mux_out[9][0] })
         );
  MUX51_GENERIC_N64_6 mux_i_10 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n569, n569, 
        n569, n568, n568, n568, n568, n568, n568, n568, n567, n567, n567, n500, 
        n490, n480, n470, n460, n450, n440, n430, n420, n410, n400, n390, n380, 
        n370, n360, n350, n340, n330, n320, n310, n300, n290, n280, n270, n260, 
        n250, n240, n230, n220, n210, n200, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n647, n647, n648, n648, n648, n648, n648, n648, n648, 
        n648, n648, n648, n648, n506, n496, n486, n476, n466, n456, n446, n436, 
        n426, n416, n406, n396, n386, n376, n366, n356, n346, n336, n326, n316, 
        n306, n296, n286, n276, n266, n256, n246, n236, n226, n216, n206, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n567, n567, n567, n567, 
        n566, n566, n566, n566, n566, n566, n566, n565, n500, n490, n480, n470, 
        n460, n450, n440, n430, n420, n410, n400, n390, n380, n370, n360, n350, 
        n340, n330, n320, n310, n300, n290, n280, n270, n260, n250, n240, n230, 
        n220, n210, n200, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n665, n665, n665, n665, n666, n666, n666, n666, n666, n666, n666, n666, 
        n506, n496, n486, n476, n466, n456, n446, n436, n426, n416, n406, n396, 
        n386, n376, n366, n356, n346, n336, n326, n316, n306, n296, n286, n276, 
        n266, n256, n246, n236, n226, n216, n206, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[32:30]), .Y({
        \mux_out[10][63] , \mux_out[10][62] , \mux_out[10][61] , 
        \mux_out[10][60] , \mux_out[10][59] , \mux_out[10][58] , 
        \mux_out[10][57] , \mux_out[10][56] , \mux_out[10][55] , 
        \mux_out[10][54] , \mux_out[10][53] , \mux_out[10][52] , 
        \mux_out[10][51] , \mux_out[10][50] , \mux_out[10][49] , 
        \mux_out[10][48] , \mux_out[10][47] , \mux_out[10][46] , 
        \mux_out[10][45] , \mux_out[10][44] , \mux_out[10][43] , 
        \mux_out[10][42] , \mux_out[10][41] , \mux_out[10][40] , 
        \mux_out[10][39] , \mux_out[10][38] , \mux_out[10][37] , 
        \mux_out[10][36] , \mux_out[10][35] , \mux_out[10][34] , 
        \mux_out[10][33] , \mux_out[10][32] , \mux_out[10][31] , 
        \mux_out[10][30] , \mux_out[10][29] , \mux_out[10][28] , 
        \mux_out[10][27] , \mux_out[10][26] , \mux_out[10][25] , 
        \mux_out[10][24] , \mux_out[10][23] , \mux_out[10][22] , 
        \mux_out[10][21] , \mux_out[10][20] , \mux_out[10][19] , 
        \mux_out[10][18] , \mux_out[10][17] , \mux_out[10][16] , 
        \mux_out[10][15] , \mux_out[10][14] , \mux_out[10][13] , 
        \mux_out[10][12] , \mux_out[10][11] , \mux_out[10][10] , 
        \mux_out[10][9] , \mux_out[10][8] , \mux_out[10][7] , \mux_out[10][6] , 
        \mux_out[10][5] , \mux_out[10][4] , \mux_out[10][3] , \mux_out[10][2] , 
        \mux_out[10][1] , \mux_out[10][0] }) );
  MUX51_GENERIC_N64_5 mux_i_11 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n572, n572, 
        n572, n571, n571, n571, n571, n571, n571, n571, n570, n501, n491, n481, 
        n471, n461, n451, n441, n431, n421, n411, n401, n391, n381, n371, n361, 
        n351, n341, n331, n321, n311, n301, n291, n281, n271, n261, n251, n241, 
        n231, n221, n211, n201, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n648, n649, n649, n649, n649, n649, n649, n649, n649, 
        n649, n649, n506, n496, n486, n476, n466, n456, n446, n436, n426, n416, 
        n406, n396, n386, n376, n366, n356, n346, n336, n326, n316, n306, n296, 
        n286, n276, n266, n256, n246, n236, n226, n216, n206, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n570, n570, n570, n570, 
        n570, n570, n569, n569, n569, n569, n500, n490, n480, n470, n460, n450, 
        n440, n430, n420, n410, n400, n390, n380, n370, n360, n350, n340, n330, 
        n320, n310, n300, n290, n280, n270, n260, n250, n240, n230, n220, n210, 
        n200, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n666, n667, n667, n667, n667, n667, n667, n667, n667, n667, n506, n496, 
        n486, n476, n466, n456, n446, n436, n426, n416, n406, n396, n386, n376, 
        n366, n356, n346, n336, n326, n316, n306, n296, n286, n276, n266, n256, 
        n246, n236, n226, n216, n206, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[35:33]), .Y({
        \mux_out[11][63] , \mux_out[11][62] , \mux_out[11][61] , 
        \mux_out[11][60] , \mux_out[11][59] , \mux_out[11][58] , 
        \mux_out[11][57] , \mux_out[11][56] , \mux_out[11][55] , 
        \mux_out[11][54] , \mux_out[11][53] , \mux_out[11][52] , 
        \mux_out[11][51] , \mux_out[11][50] , \mux_out[11][49] , 
        \mux_out[11][48] , \mux_out[11][47] , \mux_out[11][46] , 
        \mux_out[11][45] , \mux_out[11][44] , \mux_out[11][43] , 
        \mux_out[11][42] , \mux_out[11][41] , \mux_out[11][40] , 
        \mux_out[11][39] , \mux_out[11][38] , \mux_out[11][37] , 
        \mux_out[11][36] , \mux_out[11][35] , \mux_out[11][34] , 
        \mux_out[11][33] , \mux_out[11][32] , \mux_out[11][31] , 
        \mux_out[11][30] , \mux_out[11][29] , \mux_out[11][28] , 
        \mux_out[11][27] , \mux_out[11][26] , \mux_out[11][25] , 
        \mux_out[11][24] , \mux_out[11][23] , \mux_out[11][22] , 
        \mux_out[11][21] , \mux_out[11][20] , \mux_out[11][19] , 
        \mux_out[11][18] , \mux_out[11][17] , \mux_out[11][16] , 
        \mux_out[11][15] , \mux_out[11][14] , \mux_out[11][13] , 
        \mux_out[11][12] , \mux_out[11][11] , \mux_out[11][10] , 
        \mux_out[11][9] , \mux_out[11][8] , \mux_out[11][7] , \mux_out[11][6] , 
        \mux_out[11][5] , \mux_out[11][4] , \mux_out[11][3] , \mux_out[11][2] , 
        \mux_out[11][1] , \mux_out[11][0] }) );
  MUX51_GENERIC_N64_4 mux_i_12 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n574, n574, 
        n574, n574, n574, n574, n573, n573, n573, n501, n491, n481, n471, n461, 
        n451, n441, n431, n421, n411, n401, n391, n381, n371, n361, n351, n341, 
        n331, n321, n311, n301, n291, n281, n271, n261, n251, n241, n231, n221, 
        n211, n201, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n649, n649, n650, n650, n650, n650, n650, n650, n650, 
        n505, n495, n485, n475, n465, n455, n445, n435, n425, n415, n405, n395, 
        n385, n375, n365, n355, n345, n335, n325, n315, n305, n295, n285, n275, 
        n265, n255, n245, n235, n225, n215, n205, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n573, n573, n573, n573, 
        n572, n572, n572, n572, n501, n491, n481, n471, n461, n451, n441, n431, 
        n421, n411, n401, n391, n381, n371, n361, n351, n341, n331, n321, n311, 
        n301, n291, n281, n271, n261, n251, n241, n231, n221, n211, n201, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n667, n667, n667, n668, n668, n668, n668, n668, n506, n496, n486, n476, 
        n466, n456, n446, n436, n426, n416, n406, n396, n386, n376, n366, n356, 
        n346, n336, n326, n316, n306, n296, n286, n276, n266, n256, n246, n236, 
        n226, n216, n206, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[38:36]), .Y({
        \mux_out[12][63] , \mux_out[12][62] , \mux_out[12][61] , 
        \mux_out[12][60] , \mux_out[12][59] , \mux_out[12][58] , 
        \mux_out[12][57] , \mux_out[12][56] , \mux_out[12][55] , 
        \mux_out[12][54] , \mux_out[12][53] , \mux_out[12][52] , 
        \mux_out[12][51] , \mux_out[12][50] , \mux_out[12][49] , 
        \mux_out[12][48] , \mux_out[12][47] , \mux_out[12][46] , 
        \mux_out[12][45] , \mux_out[12][44] , \mux_out[12][43] , 
        \mux_out[12][42] , \mux_out[12][41] , \mux_out[12][40] , 
        \mux_out[12][39] , \mux_out[12][38] , \mux_out[12][37] , 
        \mux_out[12][36] , \mux_out[12][35] , \mux_out[12][34] , 
        \mux_out[12][33] , \mux_out[12][32] , \mux_out[12][31] , 
        \mux_out[12][30] , \mux_out[12][29] , \mux_out[12][28] , 
        \mux_out[12][27] , \mux_out[12][26] , \mux_out[12][25] , 
        \mux_out[12][24] , \mux_out[12][23] , \mux_out[12][22] , 
        \mux_out[12][21] , \mux_out[12][20] , \mux_out[12][19] , 
        \mux_out[12][18] , \mux_out[12][17] , \mux_out[12][16] , 
        \mux_out[12][15] , \mux_out[12][14] , \mux_out[12][13] , 
        \mux_out[12][12] , \mux_out[12][11] , \mux_out[12][10] , 
        \mux_out[12][9] , \mux_out[12][8] , \mux_out[12][7] , \mux_out[12][6] , 
        \mux_out[12][5] , \mux_out[12][4] , \mux_out[12][3] , \mux_out[12][2] , 
        \mux_out[12][1] , \mux_out[12][0] }) );
  MUX51_GENERIC_N64_3 mux_i_13 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n576, n576, 
        n576, n576, n576, n575, n575, n501, n491, n481, n471, n461, n451, n441, 
        n431, n421, n411, n401, n391, n381, n371, n361, n351, n341, n331, n321, 
        n311, n301, n291, n281, n271, n261, n251, n241, n231, n221, n211, n201, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n650, n650, n650, n650, n650, n651, n651, n505, n495, 
        n485, n475, n465, n455, n445, n435, n425, n415, n405, n395, n385, n375, 
        n365, n355, n345, n335, n325, n315, n305, n295, n285, n275, n265, n255, 
        n245, n235, n225, n215, n205, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n575, n575, n575, n575, 
        n575, n574, n501, n491, n481, n471, n461, n451, n441, n431, n421, n411, 
        n401, n391, n381, n371, n361, n351, n341, n331, n321, n311, n301, n291, 
        n281, n271, n261, n251, n241, n231, n221, n211, n201, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n668, n668, n668, n668, n668, n668, n506, n496, n486, n476, n466, n456, 
        n446, n436, n426, n416, n406, n396, n386, n376, n366, n356, n346, n336, 
        n326, n316, n306, n296, n286, n276, n266, n256, n246, n236, n226, n216, 
        n206, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[41:39]), .Y({
        \mux_out[13][63] , \mux_out[13][62] , \mux_out[13][61] , 
        \mux_out[13][60] , \mux_out[13][59] , \mux_out[13][58] , 
        \mux_out[13][57] , \mux_out[13][56] , \mux_out[13][55] , 
        \mux_out[13][54] , \mux_out[13][53] , \mux_out[13][52] , 
        \mux_out[13][51] , \mux_out[13][50] , \mux_out[13][49] , 
        \mux_out[13][48] , \mux_out[13][47] , \mux_out[13][46] , 
        \mux_out[13][45] , \mux_out[13][44] , \mux_out[13][43] , 
        \mux_out[13][42] , \mux_out[13][41] , \mux_out[13][40] , 
        \mux_out[13][39] , \mux_out[13][38] , \mux_out[13][37] , 
        \mux_out[13][36] , \mux_out[13][35] , \mux_out[13][34] , 
        \mux_out[13][33] , \mux_out[13][32] , \mux_out[13][31] , 
        \mux_out[13][30] , \mux_out[13][29] , \mux_out[13][28] , 
        \mux_out[13][27] , \mux_out[13][26] , \mux_out[13][25] , 
        \mux_out[13][24] , \mux_out[13][23] , \mux_out[13][22] , 
        \mux_out[13][21] , \mux_out[13][20] , \mux_out[13][19] , 
        \mux_out[13][18] , \mux_out[13][17] , \mux_out[13][16] , 
        \mux_out[13][15] , \mux_out[13][14] , \mux_out[13][13] , 
        \mux_out[13][12] , \mux_out[13][11] , \mux_out[13][10] , 
        \mux_out[13][9] , \mux_out[13][8] , \mux_out[13][7] , \mux_out[13][6] , 
        \mux_out[13][5] , \mux_out[13][4] , \mux_out[13][3] , \mux_out[13][2] , 
        \mux_out[13][1] , \mux_out[13][0] }) );
  MUX51_GENERIC_N64_2 mux_i_14 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n577, n577, 
        n577, n577, n577, n501, n491, n481, n471, n461, n451, n441, n431, n421, 
        n411, n401, n391, n381, n371, n361, n351, n341, n331, n321, n311, n301, 
        n291, n281, n271, n261, n251, n241, n231, n221, n211, n201, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n651, n651, n651, n651, n651, n505, n495, n485, n475, 
        n465, n455, n445, n435, n425, n415, n405, n395, n385, n375, n365, n355, 
        n345, n335, n325, n315, n305, n295, n285, n275, n265, n255, n245, n235, 
        n225, n215, n205, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n577, n577, n576, n576, 
        n501, n491, n481, n471, n461, n451, n441, n431, n421, n411, n401, n391, 
        n381, n371, n361, n351, n341, n331, n321, n311, n301, n291, n281, n271, 
        n261, n251, n241, n231, n221, n211, n201, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n668, n669, n669, n669, n506, n496, n486, n476, n466, n456, n446, n436, 
        n426, n416, n406, n396, n386, n376, n366, n356, n346, n336, n326, n316, 
        n306, n296, n286, n276, n266, n256, n246, n236, n226, n216, n206, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[44:42]), .Y({
        \mux_out[14][63] , \mux_out[14][62] , \mux_out[14][61] , 
        \mux_out[14][60] , \mux_out[14][59] , \mux_out[14][58] , 
        \mux_out[14][57] , \mux_out[14][56] , \mux_out[14][55] , 
        \mux_out[14][54] , \mux_out[14][53] , \mux_out[14][52] , 
        \mux_out[14][51] , \mux_out[14][50] , \mux_out[14][49] , 
        \mux_out[14][48] , \mux_out[14][47] , \mux_out[14][46] , 
        \mux_out[14][45] , \mux_out[14][44] , \mux_out[14][43] , 
        \mux_out[14][42] , \mux_out[14][41] , \mux_out[14][40] , 
        \mux_out[14][39] , \mux_out[14][38] , \mux_out[14][37] , 
        \mux_out[14][36] , \mux_out[14][35] , \mux_out[14][34] , 
        \mux_out[14][33] , \mux_out[14][32] , \mux_out[14][31] , 
        \mux_out[14][30] , \mux_out[14][29] , \mux_out[14][28] , 
        \mux_out[14][27] , \mux_out[14][26] , \mux_out[14][25] , 
        \mux_out[14][24] , \mux_out[14][23] , \mux_out[14][22] , 
        \mux_out[14][21] , \mux_out[14][20] , \mux_out[14][19] , 
        \mux_out[14][18] , \mux_out[14][17] , \mux_out[14][16] , 
        \mux_out[14][15] , \mux_out[14][14] , \mux_out[14][13] , 
        \mux_out[14][12] , \mux_out[14][11] , \mux_out[14][10] , 
        \mux_out[14][9] , \mux_out[14][8] , \mux_out[14][7] , \mux_out[14][6] , 
        \mux_out[14][5] , \mux_out[14][4] , \mux_out[14][3] , \mux_out[14][2] , 
        \mux_out[14][1] , \mux_out[14][0] }) );
  MUX51_GENERIC_N64_1 mux_i_15 ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({n578, n578, 
        n578, n502, n492, n482, n472, n462, n452, n442, n432, n422, n412, n402, 
        n392, n382, n372, n362, n352, n342, n332, n322, n312, n302, n292, n282, 
        n272, n262, n252, n242, n232, n222, n212, n202, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .C({n651, n651, n636, n505, n495, n485, n475, n465, n455, 
        n445, n435, n425, n415, n405, n395, n385, n375, n365, n355, n345, n335, 
        n325, n315, n305, n295, n285, n275, n265, n255, n245, n235, n225, n215, 
        n205, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .D({n578, n578, n502, n492, 
        n482, n472, n462, n452, n442, n432, n422, n412, n402, n392, n382, n372, 
        n362, n352, n342, n332, n322, n312, n302, n292, n282, n272, n262, n252, 
        n242, n232, n222, n212, n202, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .E({n669, n669, n506, n496, n486, n476, n466, n456, n446, n436, n426, n416, 
        n406, n396, n386, n376, n366, n356, n346, n336, n326, n316, n306, n296, 
        n286, n276, n266, n256, n246, n236, n226, n216, n206, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .SEL(encoder_out[47:45]), .Y({
        \mux_out[15][63] , \mux_out[15][62] , \mux_out[15][61] , 
        \mux_out[15][60] , \mux_out[15][59] , \mux_out[15][58] , 
        \mux_out[15][57] , \mux_out[15][56] , \mux_out[15][55] , 
        \mux_out[15][54] , \mux_out[15][53] , \mux_out[15][52] , 
        \mux_out[15][51] , \mux_out[15][50] , \mux_out[15][49] , 
        \mux_out[15][48] , \mux_out[15][47] , \mux_out[15][46] , 
        \mux_out[15][45] , \mux_out[15][44] , \mux_out[15][43] , 
        \mux_out[15][42] , \mux_out[15][41] , \mux_out[15][40] , 
        \mux_out[15][39] , \mux_out[15][38] , \mux_out[15][37] , 
        \mux_out[15][36] , \mux_out[15][35] , \mux_out[15][34] , 
        \mux_out[15][33] , \mux_out[15][32] , \mux_out[15][31] , 
        \mux_out[15][30] , \mux_out[15][29] , \mux_out[15][28] , 
        \mux_out[15][27] , \mux_out[15][26] , \mux_out[15][25] , 
        \mux_out[15][24] , \mux_out[15][23] , \mux_out[15][22] , 
        \mux_out[15][21] , \mux_out[15][20] , \mux_out[15][19] , 
        \mux_out[15][18] , \mux_out[15][17] , \mux_out[15][16] , 
        \mux_out[15][15] , \mux_out[15][14] , \mux_out[15][13] , 
        \mux_out[15][12] , \mux_out[15][11] , \mux_out[15][10] , 
        \mux_out[15][9] , \mux_out[15][8] , \mux_out[15][7] , \mux_out[15][6] , 
        \mux_out[15][5] , \mux_out[15][4] , \mux_out[15][3] , \mux_out[15][2] , 
        \mux_out[15][1] , \mux_out[15][0] }) );
  RCA_generic_N64_0 add_i_0 ( .A({\mux_out[1][63] , \mux_out[1][62] , 
        \mux_out[1][61] , \mux_out[1][60] , \mux_out[1][59] , \mux_out[1][58] , 
        \mux_out[1][57] , \mux_out[1][56] , \mux_out[1][55] , \mux_out[1][54] , 
        \mux_out[1][53] , \mux_out[1][52] , \mux_out[1][51] , \mux_out[1][50] , 
        \mux_out[1][49] , \mux_out[1][48] , \mux_out[1][47] , \mux_out[1][46] , 
        \mux_out[1][45] , \mux_out[1][44] , \mux_out[1][43] , \mux_out[1][42] , 
        \mux_out[1][41] , \mux_out[1][40] , \mux_out[1][39] , \mux_out[1][38] , 
        \mux_out[1][37] , \mux_out[1][36] , \mux_out[1][35] , \mux_out[1][34] , 
        \mux_out[1][33] , \mux_out[1][32] , \mux_out[1][31] , \mux_out[1][30] , 
        \mux_out[1][29] , \mux_out[1][28] , \mux_out[1][27] , \mux_out[1][26] , 
        \mux_out[1][25] , \mux_out[1][24] , \mux_out[1][23] , \mux_out[1][22] , 
        \mux_out[1][21] , \mux_out[1][20] , \mux_out[1][19] , \mux_out[1][18] , 
        \mux_out[1][17] , \mux_out[1][16] , \mux_out[1][15] , \mux_out[1][14] , 
        \mux_out[1][13] , \mux_out[1][12] , \mux_out[1][11] , \mux_out[1][10] , 
        \mux_out[1][9] , \mux_out[1][8] , \mux_out[1][7] , \mux_out[1][6] , 
        \mux_out[1][5] , \mux_out[1][4] , \mux_out[1][3] , \mux_out[1][2] , 
        \mux_out[1][1] , \mux_out[1][0] }), .B({\add_in[0][63] , 
        \add_in[0][62] , \add_in[0][61] , \add_in[0][60] , \add_in[0][59] , 
        \add_in[0][58] , \add_in[0][57] , \add_in[0][56] , \add_in[0][55] , 
        \add_in[0][54] , \add_in[0][53] , \add_in[0][52] , \add_in[0][51] , 
        \add_in[0][50] , \add_in[0][49] , \add_in[0][48] , \add_in[0][47] , 
        \add_in[0][46] , \add_in[0][45] , \add_in[0][44] , \add_in[0][43] , 
        \add_in[0][42] , \add_in[0][41] , \add_in[0][40] , \add_in[0][39] , 
        \add_in[0][38] , \add_in[0][37] , \add_in[0][36] , \add_in[0][35] , 
        \add_in[0][34] , \add_in[0][33] , \add_in[0][32] , \add_in[0][31] , 
        \add_in[0][30] , \add_in[0][29] , \add_in[0][28] , \add_in[0][27] , 
        \add_in[0][26] , \add_in[0][25] , \add_in[0][24] , \add_in[0][23] , 
        \add_in[0][22] , \add_in[0][21] , \add_in[0][20] , \add_in[0][19] , 
        \add_in[0][18] , \add_in[0][17] , \add_in[0][16] , \add_in[0][15] , 
        \add_in[0][14] , \add_in[0][13] , \add_in[0][12] , \add_in[0][11] , 
        \add_in[0][10] , \add_in[0][9] , \add_in[0][8] , \add_in[0][7] , 
        \add_in[0][6] , \add_in[0][5] , \add_in[0][4] , \add_in[0][3] , 
        \add_in[0][2] , \add_in[0][1] , \add_in[0][0] }), .Ci(mode[0]), .S({
        \add_in[1][63] , \add_in[1][62] , \add_in[1][61] , \add_in[1][60] , 
        \add_in[1][59] , \add_in[1][58] , \add_in[1][57] , \add_in[1][56] , 
        \add_in[1][55] , \add_in[1][54] , \add_in[1][53] , \add_in[1][52] , 
        \add_in[1][51] , \add_in[1][50] , \add_in[1][49] , \add_in[1][48] , 
        \add_in[1][47] , \add_in[1][46] , \add_in[1][45] , \add_in[1][44] , 
        \add_in[1][43] , \add_in[1][42] , \add_in[1][41] , \add_in[1][40] , 
        \add_in[1][39] , \add_in[1][38] , \add_in[1][37] , \add_in[1][36] , 
        \add_in[1][35] , \add_in[1][34] , \add_in[1][33] , \add_in[1][32] , 
        \add_in[1][31] , \add_in[1][30] , \add_in[1][29] , \add_in[1][28] , 
        \add_in[1][27] , \add_in[1][26] , \add_in[1][25] , \add_in[1][24] , 
        \add_in[1][23] , \add_in[1][22] , \add_in[1][21] , \add_in[1][20] , 
        \add_in[1][19] , \add_in[1][18] , \add_in[1][17] , \add_in[1][16] , 
        \add_in[1][15] , \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , 
        \add_in[1][11] , \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , 
        \add_in[1][7] , \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , 
        \add_in[1][3] , \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }) );
  RCA_generic_N64_14 add_i_1 ( .A({\mux_out[2][63] , \mux_out[2][62] , 
        \mux_out[2][61] , \mux_out[2][60] , \mux_out[2][59] , \mux_out[2][58] , 
        \mux_out[2][57] , \mux_out[2][56] , \mux_out[2][55] , \mux_out[2][54] , 
        \mux_out[2][53] , \mux_out[2][52] , \mux_out[2][51] , \mux_out[2][50] , 
        \mux_out[2][49] , \mux_out[2][48] , \mux_out[2][47] , \mux_out[2][46] , 
        \mux_out[2][45] , \mux_out[2][44] , \mux_out[2][43] , \mux_out[2][42] , 
        \mux_out[2][41] , \mux_out[2][40] , \mux_out[2][39] , \mux_out[2][38] , 
        \mux_out[2][37] , \mux_out[2][36] , \mux_out[2][35] , \mux_out[2][34] , 
        \mux_out[2][33] , \mux_out[2][32] , \mux_out[2][31] , \mux_out[2][30] , 
        \mux_out[2][29] , \mux_out[2][28] , \mux_out[2][27] , \mux_out[2][26] , 
        \mux_out[2][25] , \mux_out[2][24] , \mux_out[2][23] , \mux_out[2][22] , 
        \mux_out[2][21] , \mux_out[2][20] , \mux_out[2][19] , \mux_out[2][18] , 
        \mux_out[2][17] , \mux_out[2][16] , \mux_out[2][15] , \mux_out[2][14] , 
        \mux_out[2][13] , \mux_out[2][12] , \mux_out[2][11] , \mux_out[2][10] , 
        \mux_out[2][9] , \mux_out[2][8] , \mux_out[2][7] , \mux_out[2][6] , 
        \mux_out[2][5] , \mux_out[2][4] , \mux_out[2][3] , \mux_out[2][2] , 
        \mux_out[2][1] , \mux_out[2][0] }), .B({\add_in[1][63] , 
        \add_in[1][62] , \add_in[1][61] , \add_in[1][60] , \add_in[1][59] , 
        \add_in[1][58] , \add_in[1][57] , \add_in[1][56] , \add_in[1][55] , 
        \add_in[1][54] , \add_in[1][53] , \add_in[1][52] , \add_in[1][51] , 
        \add_in[1][50] , \add_in[1][49] , \add_in[1][48] , \add_in[1][47] , 
        \add_in[1][46] , \add_in[1][45] , \add_in[1][44] , \add_in[1][43] , 
        \add_in[1][42] , \add_in[1][41] , \add_in[1][40] , \add_in[1][39] , 
        \add_in[1][38] , \add_in[1][37] , \add_in[1][36] , \add_in[1][35] , 
        \add_in[1][34] , \add_in[1][33] , \add_in[1][32] , \add_in[1][31] , 
        \add_in[1][30] , \add_in[1][29] , \add_in[1][28] , \add_in[1][27] , 
        \add_in[1][26] , \add_in[1][25] , \add_in[1][24] , \add_in[1][23] , 
        \add_in[1][22] , \add_in[1][21] , \add_in[1][20] , \add_in[1][19] , 
        \add_in[1][18] , \add_in[1][17] , \add_in[1][16] , \add_in[1][15] , 
        \add_in[1][14] , \add_in[1][13] , \add_in[1][12] , \add_in[1][11] , 
        \add_in[1][10] , \add_in[1][9] , \add_in[1][8] , \add_in[1][7] , 
        \add_in[1][6] , \add_in[1][5] , \add_in[1][4] , \add_in[1][3] , 
        \add_in[1][2] , \add_in[1][1] , \add_in[1][0] }), .Ci(mode[1]), .S({
        \add_in[2][63] , \add_in[2][62] , \add_in[2][61] , \add_in[2][60] , 
        \add_in[2][59] , \add_in[2][58] , \add_in[2][57] , \add_in[2][56] , 
        \add_in[2][55] , \add_in[2][54] , \add_in[2][53] , \add_in[2][52] , 
        \add_in[2][51] , \add_in[2][50] , \add_in[2][49] , \add_in[2][48] , 
        \add_in[2][47] , \add_in[2][46] , \add_in[2][45] , \add_in[2][44] , 
        \add_in[2][43] , \add_in[2][42] , \add_in[2][41] , \add_in[2][40] , 
        \add_in[2][39] , \add_in[2][38] , \add_in[2][37] , \add_in[2][36] , 
        \add_in[2][35] , \add_in[2][34] , \add_in[2][33] , \add_in[2][32] , 
        \add_in[2][31] , \add_in[2][30] , \add_in[2][29] , \add_in[2][28] , 
        \add_in[2][27] , \add_in[2][26] , \add_in[2][25] , \add_in[2][24] , 
        \add_in[2][23] , \add_in[2][22] , \add_in[2][21] , \add_in[2][20] , 
        \add_in[2][19] , \add_in[2][18] , \add_in[2][17] , \add_in[2][16] , 
        \add_in[2][15] , \add_in[2][14] , \add_in[2][13] , \add_in[2][12] , 
        \add_in[2][11] , \add_in[2][10] , \add_in[2][9] , \add_in[2][8] , 
        \add_in[2][7] , \add_in[2][6] , \add_in[2][5] , \add_in[2][4] , 
        \add_in[2][3] , \add_in[2][2] , \add_in[2][1] , \add_in[2][0] }) );
  RCA_generic_N64_13 add_i_2 ( .A({\mux_out[3][63] , \mux_out[3][62] , 
        \mux_out[3][61] , \mux_out[3][60] , \mux_out[3][59] , \mux_out[3][58] , 
        \mux_out[3][57] , \mux_out[3][56] , \mux_out[3][55] , \mux_out[3][54] , 
        \mux_out[3][53] , \mux_out[3][52] , \mux_out[3][51] , \mux_out[3][50] , 
        \mux_out[3][49] , \mux_out[3][48] , \mux_out[3][47] , \mux_out[3][46] , 
        \mux_out[3][45] , \mux_out[3][44] , \mux_out[3][43] , \mux_out[3][42] , 
        \mux_out[3][41] , \mux_out[3][40] , \mux_out[3][39] , \mux_out[3][38] , 
        \mux_out[3][37] , \mux_out[3][36] , \mux_out[3][35] , \mux_out[3][34] , 
        \mux_out[3][33] , \mux_out[3][32] , \mux_out[3][31] , \mux_out[3][30] , 
        \mux_out[3][29] , \mux_out[3][28] , \mux_out[3][27] , \mux_out[3][26] , 
        \mux_out[3][25] , \mux_out[3][24] , \mux_out[3][23] , \mux_out[3][22] , 
        \mux_out[3][21] , \mux_out[3][20] , \mux_out[3][19] , \mux_out[3][18] , 
        \mux_out[3][17] , \mux_out[3][16] , \mux_out[3][15] , \mux_out[3][14] , 
        \mux_out[3][13] , \mux_out[3][12] , \mux_out[3][11] , \mux_out[3][10] , 
        \mux_out[3][9] , \mux_out[3][8] , \mux_out[3][7] , \mux_out[3][6] , 
        \mux_out[3][5] , \mux_out[3][4] , \mux_out[3][3] , \mux_out[3][2] , 
        \mux_out[3][1] , \mux_out[3][0] }), .B({\add_in[2][63] , 
        \add_in[2][62] , \add_in[2][61] , \add_in[2][60] , \add_in[2][59] , 
        \add_in[2][58] , \add_in[2][57] , \add_in[2][56] , \add_in[2][55] , 
        \add_in[2][54] , \add_in[2][53] , \add_in[2][52] , \add_in[2][51] , 
        \add_in[2][50] , \add_in[2][49] , \add_in[2][48] , \add_in[2][47] , 
        \add_in[2][46] , \add_in[2][45] , \add_in[2][44] , \add_in[2][43] , 
        \add_in[2][42] , \add_in[2][41] , \add_in[2][40] , \add_in[2][39] , 
        \add_in[2][38] , \add_in[2][37] , \add_in[2][36] , \add_in[2][35] , 
        \add_in[2][34] , \add_in[2][33] , \add_in[2][32] , \add_in[2][31] , 
        \add_in[2][30] , \add_in[2][29] , \add_in[2][28] , \add_in[2][27] , 
        \add_in[2][26] , \add_in[2][25] , \add_in[2][24] , \add_in[2][23] , 
        \add_in[2][22] , \add_in[2][21] , \add_in[2][20] , \add_in[2][19] , 
        \add_in[2][18] , \add_in[2][17] , \add_in[2][16] , \add_in[2][15] , 
        \add_in[2][14] , \add_in[2][13] , \add_in[2][12] , \add_in[2][11] , 
        \add_in[2][10] , \add_in[2][9] , \add_in[2][8] , \add_in[2][7] , 
        \add_in[2][6] , \add_in[2][5] , \add_in[2][4] , \add_in[2][3] , 
        \add_in[2][2] , \add_in[2][1] , \add_in[2][0] }), .Ci(mode[2]), .S({
        \add_in[3][63] , \add_in[3][62] , \add_in[3][61] , \add_in[3][60] , 
        \add_in[3][59] , \add_in[3][58] , \add_in[3][57] , \add_in[3][56] , 
        \add_in[3][55] , \add_in[3][54] , \add_in[3][53] , \add_in[3][52] , 
        \add_in[3][51] , \add_in[3][50] , \add_in[3][49] , \add_in[3][48] , 
        \add_in[3][47] , \add_in[3][46] , \add_in[3][45] , \add_in[3][44] , 
        \add_in[3][43] , \add_in[3][42] , \add_in[3][41] , \add_in[3][40] , 
        \add_in[3][39] , \add_in[3][38] , \add_in[3][37] , \add_in[3][36] , 
        \add_in[3][35] , \add_in[3][34] , \add_in[3][33] , \add_in[3][32] , 
        \add_in[3][31] , \add_in[3][30] , \add_in[3][29] , \add_in[3][28] , 
        \add_in[3][27] , \add_in[3][26] , \add_in[3][25] , \add_in[3][24] , 
        \add_in[3][23] , \add_in[3][22] , \add_in[3][21] , \add_in[3][20] , 
        \add_in[3][19] , \add_in[3][18] , \add_in[3][17] , \add_in[3][16] , 
        \add_in[3][15] , \add_in[3][14] , \add_in[3][13] , \add_in[3][12] , 
        \add_in[3][11] , \add_in[3][10] , \add_in[3][9] , \add_in[3][8] , 
        \add_in[3][7] , \add_in[3][6] , \add_in[3][5] , \add_in[3][4] , 
        \add_in[3][3] , \add_in[3][2] , \add_in[3][1] , \add_in[3][0] }) );
  RCA_generic_N64_12 add_i_3 ( .A({\mux_out[4][63] , \mux_out[4][62] , 
        \mux_out[4][61] , \mux_out[4][60] , \mux_out[4][59] , \mux_out[4][58] , 
        \mux_out[4][57] , \mux_out[4][56] , \mux_out[4][55] , \mux_out[4][54] , 
        \mux_out[4][53] , \mux_out[4][52] , \mux_out[4][51] , \mux_out[4][50] , 
        \mux_out[4][49] , \mux_out[4][48] , \mux_out[4][47] , \mux_out[4][46] , 
        \mux_out[4][45] , \mux_out[4][44] , \mux_out[4][43] , \mux_out[4][42] , 
        \mux_out[4][41] , \mux_out[4][40] , \mux_out[4][39] , \mux_out[4][38] , 
        \mux_out[4][37] , \mux_out[4][36] , \mux_out[4][35] , \mux_out[4][34] , 
        \mux_out[4][33] , \mux_out[4][32] , \mux_out[4][31] , \mux_out[4][30] , 
        \mux_out[4][29] , \mux_out[4][28] , \mux_out[4][27] , \mux_out[4][26] , 
        \mux_out[4][25] , \mux_out[4][24] , \mux_out[4][23] , \mux_out[4][22] , 
        \mux_out[4][21] , \mux_out[4][20] , \mux_out[4][19] , \mux_out[4][18] , 
        \mux_out[4][17] , \mux_out[4][16] , \mux_out[4][15] , \mux_out[4][14] , 
        \mux_out[4][13] , \mux_out[4][12] , \mux_out[4][11] , \mux_out[4][10] , 
        \mux_out[4][9] , \mux_out[4][8] , \mux_out[4][7] , \mux_out[4][6] , 
        \mux_out[4][5] , \mux_out[4][4] , \mux_out[4][3] , \mux_out[4][2] , 
        \mux_out[4][1] , \mux_out[4][0] }), .B({\add_in[3][63] , 
        \add_in[3][62] , \add_in[3][61] , \add_in[3][60] , \add_in[3][59] , 
        \add_in[3][58] , \add_in[3][57] , \add_in[3][56] , \add_in[3][55] , 
        \add_in[3][54] , \add_in[3][53] , \add_in[3][52] , \add_in[3][51] , 
        \add_in[3][50] , \add_in[3][49] , \add_in[3][48] , \add_in[3][47] , 
        \add_in[3][46] , \add_in[3][45] , \add_in[3][44] , \add_in[3][43] , 
        \add_in[3][42] , \add_in[3][41] , \add_in[3][40] , \add_in[3][39] , 
        \add_in[3][38] , \add_in[3][37] , \add_in[3][36] , \add_in[3][35] , 
        \add_in[3][34] , \add_in[3][33] , \add_in[3][32] , \add_in[3][31] , 
        \add_in[3][30] , \add_in[3][29] , \add_in[3][28] , \add_in[3][27] , 
        \add_in[3][26] , \add_in[3][25] , \add_in[3][24] , \add_in[3][23] , 
        \add_in[3][22] , \add_in[3][21] , \add_in[3][20] , \add_in[3][19] , 
        \add_in[3][18] , \add_in[3][17] , \add_in[3][16] , \add_in[3][15] , 
        \add_in[3][14] , \add_in[3][13] , \add_in[3][12] , \add_in[3][11] , 
        \add_in[3][10] , \add_in[3][9] , \add_in[3][8] , \add_in[3][7] , 
        \add_in[3][6] , \add_in[3][5] , \add_in[3][4] , \add_in[3][3] , 
        \add_in[3][2] , \add_in[3][1] , \add_in[3][0] }), .Ci(mode[3]), .S({
        \add_in[4][63] , \add_in[4][62] , \add_in[4][61] , \add_in[4][60] , 
        \add_in[4][59] , \add_in[4][58] , \add_in[4][57] , \add_in[4][56] , 
        \add_in[4][55] , \add_in[4][54] , \add_in[4][53] , \add_in[4][52] , 
        \add_in[4][51] , \add_in[4][50] , \add_in[4][49] , \add_in[4][48] , 
        \add_in[4][47] , \add_in[4][46] , \add_in[4][45] , \add_in[4][44] , 
        \add_in[4][43] , \add_in[4][42] , \add_in[4][41] , \add_in[4][40] , 
        \add_in[4][39] , \add_in[4][38] , \add_in[4][37] , \add_in[4][36] , 
        \add_in[4][35] , \add_in[4][34] , \add_in[4][33] , \add_in[4][32] , 
        \add_in[4][31] , \add_in[4][30] , \add_in[4][29] , \add_in[4][28] , 
        \add_in[4][27] , \add_in[4][26] , \add_in[4][25] , \add_in[4][24] , 
        \add_in[4][23] , \add_in[4][22] , \add_in[4][21] , \add_in[4][20] , 
        \add_in[4][19] , \add_in[4][18] , \add_in[4][17] , \add_in[4][16] , 
        \add_in[4][15] , \add_in[4][14] , \add_in[4][13] , \add_in[4][12] , 
        \add_in[4][11] , \add_in[4][10] , \add_in[4][9] , \add_in[4][8] , 
        \add_in[4][7] , \add_in[4][6] , \add_in[4][5] , \add_in[4][4] , 
        \add_in[4][3] , \add_in[4][2] , \add_in[4][1] , \add_in[4][0] }) );
  RCA_generic_N64_11 add_i_4 ( .A({\mux_out[5][63] , \mux_out[5][62] , 
        \mux_out[5][61] , \mux_out[5][60] , \mux_out[5][59] , \mux_out[5][58] , 
        \mux_out[5][57] , \mux_out[5][56] , \mux_out[5][55] , \mux_out[5][54] , 
        \mux_out[5][53] , \mux_out[5][52] , \mux_out[5][51] , \mux_out[5][50] , 
        \mux_out[5][49] , \mux_out[5][48] , \mux_out[5][47] , \mux_out[5][46] , 
        \mux_out[5][45] , \mux_out[5][44] , \mux_out[5][43] , \mux_out[5][42] , 
        \mux_out[5][41] , \mux_out[5][40] , \mux_out[5][39] , \mux_out[5][38] , 
        \mux_out[5][37] , \mux_out[5][36] , \mux_out[5][35] , \mux_out[5][34] , 
        \mux_out[5][33] , \mux_out[5][32] , \mux_out[5][31] , \mux_out[5][30] , 
        \mux_out[5][29] , \mux_out[5][28] , \mux_out[5][27] , \mux_out[5][26] , 
        \mux_out[5][25] , \mux_out[5][24] , \mux_out[5][23] , \mux_out[5][22] , 
        \mux_out[5][21] , \mux_out[5][20] , \mux_out[5][19] , \mux_out[5][18] , 
        \mux_out[5][17] , \mux_out[5][16] , \mux_out[5][15] , \mux_out[5][14] , 
        \mux_out[5][13] , \mux_out[5][12] , \mux_out[5][11] , \mux_out[5][10] , 
        \mux_out[5][9] , \mux_out[5][8] , \mux_out[5][7] , \mux_out[5][6] , 
        \mux_out[5][5] , \mux_out[5][4] , \mux_out[5][3] , \mux_out[5][2] , 
        \mux_out[5][1] , \mux_out[5][0] }), .B({\add_in[4][63] , 
        \add_in[4][62] , \add_in[4][61] , \add_in[4][60] , \add_in[4][59] , 
        \add_in[4][58] , \add_in[4][57] , \add_in[4][56] , \add_in[4][55] , 
        \add_in[4][54] , \add_in[4][53] , \add_in[4][52] , \add_in[4][51] , 
        \add_in[4][50] , \add_in[4][49] , \add_in[4][48] , \add_in[4][47] , 
        \add_in[4][46] , \add_in[4][45] , \add_in[4][44] , \add_in[4][43] , 
        \add_in[4][42] , \add_in[4][41] , \add_in[4][40] , \add_in[4][39] , 
        \add_in[4][38] , \add_in[4][37] , \add_in[4][36] , \add_in[4][35] , 
        \add_in[4][34] , \add_in[4][33] , \add_in[4][32] , \add_in[4][31] , 
        \add_in[4][30] , \add_in[4][29] , \add_in[4][28] , \add_in[4][27] , 
        \add_in[4][26] , \add_in[4][25] , \add_in[4][24] , \add_in[4][23] , 
        \add_in[4][22] , \add_in[4][21] , \add_in[4][20] , \add_in[4][19] , 
        \add_in[4][18] , \add_in[4][17] , \add_in[4][16] , \add_in[4][15] , 
        \add_in[4][14] , \add_in[4][13] , \add_in[4][12] , \add_in[4][11] , 
        \add_in[4][10] , \add_in[4][9] , \add_in[4][8] , \add_in[4][7] , 
        \add_in[4][6] , \add_in[4][5] , \add_in[4][4] , \add_in[4][3] , 
        \add_in[4][2] , \add_in[4][1] , \add_in[4][0] }), .Ci(mode[4]), .S({
        \add_in[5][63] , \add_in[5][62] , \add_in[5][61] , \add_in[5][60] , 
        \add_in[5][59] , \add_in[5][58] , \add_in[5][57] , \add_in[5][56] , 
        \add_in[5][55] , \add_in[5][54] , \add_in[5][53] , \add_in[5][52] , 
        \add_in[5][51] , \add_in[5][50] , \add_in[5][49] , \add_in[5][48] , 
        \add_in[5][47] , \add_in[5][46] , \add_in[5][45] , \add_in[5][44] , 
        \add_in[5][43] , \add_in[5][42] , \add_in[5][41] , \add_in[5][40] , 
        \add_in[5][39] , \add_in[5][38] , \add_in[5][37] , \add_in[5][36] , 
        \add_in[5][35] , \add_in[5][34] , \add_in[5][33] , \add_in[5][32] , 
        \add_in[5][31] , \add_in[5][30] , \add_in[5][29] , \add_in[5][28] , 
        \add_in[5][27] , \add_in[5][26] , \add_in[5][25] , \add_in[5][24] , 
        \add_in[5][23] , \add_in[5][22] , \add_in[5][21] , \add_in[5][20] , 
        \add_in[5][19] , \add_in[5][18] , \add_in[5][17] , \add_in[5][16] , 
        \add_in[5][15] , \add_in[5][14] , \add_in[5][13] , \add_in[5][12] , 
        \add_in[5][11] , \add_in[5][10] , \add_in[5][9] , \add_in[5][8] , 
        \add_in[5][7] , \add_in[5][6] , \add_in[5][5] , \add_in[5][4] , 
        \add_in[5][3] , \add_in[5][2] , \add_in[5][1] , \add_in[5][0] }) );
  RCA_generic_N64_10 add_i_5 ( .A({\mux_out[6][63] , \mux_out[6][62] , 
        \mux_out[6][61] , \mux_out[6][60] , \mux_out[6][59] , \mux_out[6][58] , 
        \mux_out[6][57] , \mux_out[6][56] , \mux_out[6][55] , \mux_out[6][54] , 
        \mux_out[6][53] , \mux_out[6][52] , \mux_out[6][51] , \mux_out[6][50] , 
        \mux_out[6][49] , \mux_out[6][48] , \mux_out[6][47] , \mux_out[6][46] , 
        \mux_out[6][45] , \mux_out[6][44] , \mux_out[6][43] , \mux_out[6][42] , 
        \mux_out[6][41] , \mux_out[6][40] , \mux_out[6][39] , \mux_out[6][38] , 
        \mux_out[6][37] , \mux_out[6][36] , \mux_out[6][35] , \mux_out[6][34] , 
        \mux_out[6][33] , \mux_out[6][32] , \mux_out[6][31] , \mux_out[6][30] , 
        \mux_out[6][29] , \mux_out[6][28] , \mux_out[6][27] , \mux_out[6][26] , 
        \mux_out[6][25] , \mux_out[6][24] , \mux_out[6][23] , \mux_out[6][22] , 
        \mux_out[6][21] , \mux_out[6][20] , \mux_out[6][19] , \mux_out[6][18] , 
        \mux_out[6][17] , \mux_out[6][16] , \mux_out[6][15] , \mux_out[6][14] , 
        \mux_out[6][13] , \mux_out[6][12] , \mux_out[6][11] , \mux_out[6][10] , 
        \mux_out[6][9] , \mux_out[6][8] , \mux_out[6][7] , \mux_out[6][6] , 
        \mux_out[6][5] , \mux_out[6][4] , \mux_out[6][3] , \mux_out[6][2] , 
        \mux_out[6][1] , \mux_out[6][0] }), .B({\add_in[5][63] , 
        \add_in[5][62] , \add_in[5][61] , \add_in[5][60] , \add_in[5][59] , 
        \add_in[5][58] , \add_in[5][57] , \add_in[5][56] , \add_in[5][55] , 
        \add_in[5][54] , \add_in[5][53] , \add_in[5][52] , \add_in[5][51] , 
        \add_in[5][50] , \add_in[5][49] , \add_in[5][48] , \add_in[5][47] , 
        \add_in[5][46] , \add_in[5][45] , \add_in[5][44] , \add_in[5][43] , 
        \add_in[5][42] , \add_in[5][41] , \add_in[5][40] , \add_in[5][39] , 
        \add_in[5][38] , \add_in[5][37] , \add_in[5][36] , \add_in[5][35] , 
        \add_in[5][34] , \add_in[5][33] , \add_in[5][32] , \add_in[5][31] , 
        \add_in[5][30] , \add_in[5][29] , \add_in[5][28] , \add_in[5][27] , 
        \add_in[5][26] , \add_in[5][25] , \add_in[5][24] , \add_in[5][23] , 
        \add_in[5][22] , \add_in[5][21] , \add_in[5][20] , \add_in[5][19] , 
        \add_in[5][18] , \add_in[5][17] , \add_in[5][16] , \add_in[5][15] , 
        \add_in[5][14] , \add_in[5][13] , \add_in[5][12] , \add_in[5][11] , 
        \add_in[5][10] , \add_in[5][9] , \add_in[5][8] , \add_in[5][7] , 
        \add_in[5][6] , \add_in[5][5] , \add_in[5][4] , \add_in[5][3] , 
        \add_in[5][2] , \add_in[5][1] , \add_in[5][0] }), .Ci(mode[5]), .S({
        \add_in[6][63] , \add_in[6][62] , \add_in[6][61] , \add_in[6][60] , 
        \add_in[6][59] , \add_in[6][58] , \add_in[6][57] , \add_in[6][56] , 
        \add_in[6][55] , \add_in[6][54] , \add_in[6][53] , \add_in[6][52] , 
        \add_in[6][51] , \add_in[6][50] , \add_in[6][49] , \add_in[6][48] , 
        \add_in[6][47] , \add_in[6][46] , \add_in[6][45] , \add_in[6][44] , 
        \add_in[6][43] , \add_in[6][42] , \add_in[6][41] , \add_in[6][40] , 
        \add_in[6][39] , \add_in[6][38] , \add_in[6][37] , \add_in[6][36] , 
        \add_in[6][35] , \add_in[6][34] , \add_in[6][33] , \add_in[6][32] , 
        \add_in[6][31] , \add_in[6][30] , \add_in[6][29] , \add_in[6][28] , 
        \add_in[6][27] , \add_in[6][26] , \add_in[6][25] , \add_in[6][24] , 
        \add_in[6][23] , \add_in[6][22] , \add_in[6][21] , \add_in[6][20] , 
        \add_in[6][19] , \add_in[6][18] , \add_in[6][17] , \add_in[6][16] , 
        \add_in[6][15] , \add_in[6][14] , \add_in[6][13] , \add_in[6][12] , 
        \add_in[6][11] , \add_in[6][10] , \add_in[6][9] , \add_in[6][8] , 
        \add_in[6][7] , \add_in[6][6] , \add_in[6][5] , \add_in[6][4] , 
        \add_in[6][3] , \add_in[6][2] , \add_in[6][1] , \add_in[6][0] }) );
  RCA_generic_N64_9 add_i_6 ( .A({\mux_out[7][63] , \mux_out[7][62] , 
        \mux_out[7][61] , \mux_out[7][60] , \mux_out[7][59] , \mux_out[7][58] , 
        \mux_out[7][57] , \mux_out[7][56] , \mux_out[7][55] , \mux_out[7][54] , 
        \mux_out[7][53] , \mux_out[7][52] , \mux_out[7][51] , \mux_out[7][50] , 
        \mux_out[7][49] , \mux_out[7][48] , \mux_out[7][47] , \mux_out[7][46] , 
        \mux_out[7][45] , \mux_out[7][44] , \mux_out[7][43] , \mux_out[7][42] , 
        \mux_out[7][41] , \mux_out[7][40] , \mux_out[7][39] , \mux_out[7][38] , 
        \mux_out[7][37] , \mux_out[7][36] , \mux_out[7][35] , \mux_out[7][34] , 
        \mux_out[7][33] , \mux_out[7][32] , \mux_out[7][31] , \mux_out[7][30] , 
        \mux_out[7][29] , \mux_out[7][28] , \mux_out[7][27] , \mux_out[7][26] , 
        \mux_out[7][25] , \mux_out[7][24] , \mux_out[7][23] , \mux_out[7][22] , 
        \mux_out[7][21] , \mux_out[7][20] , \mux_out[7][19] , \mux_out[7][18] , 
        \mux_out[7][17] , \mux_out[7][16] , \mux_out[7][15] , \mux_out[7][14] , 
        \mux_out[7][13] , \mux_out[7][12] , \mux_out[7][11] , \mux_out[7][10] , 
        \mux_out[7][9] , \mux_out[7][8] , \mux_out[7][7] , \mux_out[7][6] , 
        \mux_out[7][5] , \mux_out[7][4] , \mux_out[7][3] , \mux_out[7][2] , 
        \mux_out[7][1] , \mux_out[7][0] }), .B({\add_in[6][63] , 
        \add_in[6][62] , \add_in[6][61] , \add_in[6][60] , \add_in[6][59] , 
        \add_in[6][58] , \add_in[6][57] , \add_in[6][56] , \add_in[6][55] , 
        \add_in[6][54] , \add_in[6][53] , \add_in[6][52] , \add_in[6][51] , 
        \add_in[6][50] , \add_in[6][49] , \add_in[6][48] , \add_in[6][47] , 
        \add_in[6][46] , \add_in[6][45] , \add_in[6][44] , \add_in[6][43] , 
        \add_in[6][42] , \add_in[6][41] , \add_in[6][40] , \add_in[6][39] , 
        \add_in[6][38] , \add_in[6][37] , \add_in[6][36] , \add_in[6][35] , 
        \add_in[6][34] , \add_in[6][33] , \add_in[6][32] , \add_in[6][31] , 
        \add_in[6][30] , \add_in[6][29] , \add_in[6][28] , \add_in[6][27] , 
        \add_in[6][26] , \add_in[6][25] , \add_in[6][24] , \add_in[6][23] , 
        \add_in[6][22] , \add_in[6][21] , \add_in[6][20] , \add_in[6][19] , 
        \add_in[6][18] , \add_in[6][17] , \add_in[6][16] , \add_in[6][15] , 
        \add_in[6][14] , \add_in[6][13] , \add_in[6][12] , \add_in[6][11] , 
        \add_in[6][10] , \add_in[6][9] , \add_in[6][8] , \add_in[6][7] , 
        \add_in[6][6] , \add_in[6][5] , \add_in[6][4] , \add_in[6][3] , 
        \add_in[6][2] , \add_in[6][1] , \add_in[6][0] }), .Ci(mode[6]), .S({
        \add_in[7][63] , \add_in[7][62] , \add_in[7][61] , \add_in[7][60] , 
        \add_in[7][59] , \add_in[7][58] , \add_in[7][57] , \add_in[7][56] , 
        \add_in[7][55] , \add_in[7][54] , \add_in[7][53] , \add_in[7][52] , 
        \add_in[7][51] , \add_in[7][50] , \add_in[7][49] , \add_in[7][48] , 
        \add_in[7][47] , \add_in[7][46] , \add_in[7][45] , \add_in[7][44] , 
        \add_in[7][43] , \add_in[7][42] , \add_in[7][41] , \add_in[7][40] , 
        \add_in[7][39] , \add_in[7][38] , \add_in[7][37] , \add_in[7][36] , 
        \add_in[7][35] , \add_in[7][34] , \add_in[7][33] , \add_in[7][32] , 
        \add_in[7][31] , \add_in[7][30] , \add_in[7][29] , \add_in[7][28] , 
        \add_in[7][27] , \add_in[7][26] , \add_in[7][25] , \add_in[7][24] , 
        \add_in[7][23] , \add_in[7][22] , \add_in[7][21] , \add_in[7][20] , 
        \add_in[7][19] , \add_in[7][18] , \add_in[7][17] , \add_in[7][16] , 
        \add_in[7][15] , \add_in[7][14] , \add_in[7][13] , \add_in[7][12] , 
        \add_in[7][11] , \add_in[7][10] , \add_in[7][9] , \add_in[7][8] , 
        \add_in[7][7] , \add_in[7][6] , \add_in[7][5] , \add_in[7][4] , 
        \add_in[7][3] , \add_in[7][2] , \add_in[7][1] , \add_in[7][0] }) );
  RCA_generic_N64_8 add_i_7 ( .A({\mux_out[8][63] , \mux_out[8][62] , 
        \mux_out[8][61] , \mux_out[8][60] , \mux_out[8][59] , \mux_out[8][58] , 
        \mux_out[8][57] , \mux_out[8][56] , \mux_out[8][55] , \mux_out[8][54] , 
        \mux_out[8][53] , \mux_out[8][52] , \mux_out[8][51] , \mux_out[8][50] , 
        \mux_out[8][49] , \mux_out[8][48] , \mux_out[8][47] , \mux_out[8][46] , 
        \mux_out[8][45] , \mux_out[8][44] , \mux_out[8][43] , \mux_out[8][42] , 
        \mux_out[8][41] , \mux_out[8][40] , \mux_out[8][39] , \mux_out[8][38] , 
        \mux_out[8][37] , \mux_out[8][36] , \mux_out[8][35] , \mux_out[8][34] , 
        \mux_out[8][33] , \mux_out[8][32] , \mux_out[8][31] , \mux_out[8][30] , 
        \mux_out[8][29] , \mux_out[8][28] , \mux_out[8][27] , \mux_out[8][26] , 
        \mux_out[8][25] , \mux_out[8][24] , \mux_out[8][23] , \mux_out[8][22] , 
        \mux_out[8][21] , \mux_out[8][20] , \mux_out[8][19] , \mux_out[8][18] , 
        \mux_out[8][17] , \mux_out[8][16] , \mux_out[8][15] , \mux_out[8][14] , 
        \mux_out[8][13] , \mux_out[8][12] , \mux_out[8][11] , \mux_out[8][10] , 
        \mux_out[8][9] , \mux_out[8][8] , \mux_out[8][7] , \mux_out[8][6] , 
        \mux_out[8][5] , \mux_out[8][4] , \mux_out[8][3] , \mux_out[8][2] , 
        \mux_out[8][1] , \mux_out[8][0] }), .B({\add_in[7][63] , 
        \add_in[7][62] , \add_in[7][61] , \add_in[7][60] , \add_in[7][59] , 
        \add_in[7][58] , \add_in[7][57] , \add_in[7][56] , \add_in[7][55] , 
        \add_in[7][54] , \add_in[7][53] , \add_in[7][52] , \add_in[7][51] , 
        \add_in[7][50] , \add_in[7][49] , \add_in[7][48] , \add_in[7][47] , 
        \add_in[7][46] , \add_in[7][45] , \add_in[7][44] , \add_in[7][43] , 
        \add_in[7][42] , \add_in[7][41] , \add_in[7][40] , \add_in[7][39] , 
        \add_in[7][38] , \add_in[7][37] , \add_in[7][36] , \add_in[7][35] , 
        \add_in[7][34] , \add_in[7][33] , \add_in[7][32] , \add_in[7][31] , 
        \add_in[7][30] , \add_in[7][29] , \add_in[7][28] , \add_in[7][27] , 
        \add_in[7][26] , \add_in[7][25] , \add_in[7][24] , \add_in[7][23] , 
        \add_in[7][22] , \add_in[7][21] , \add_in[7][20] , \add_in[7][19] , 
        \add_in[7][18] , \add_in[7][17] , \add_in[7][16] , \add_in[7][15] , 
        \add_in[7][14] , \add_in[7][13] , \add_in[7][12] , \add_in[7][11] , 
        \add_in[7][10] , \add_in[7][9] , \add_in[7][8] , \add_in[7][7] , 
        \add_in[7][6] , \add_in[7][5] , \add_in[7][4] , \add_in[7][3] , 
        \add_in[7][2] , \add_in[7][1] , \add_in[7][0] }), .Ci(mode[7]), .S({
        \add_in[8][63] , \add_in[8][62] , \add_in[8][61] , \add_in[8][60] , 
        \add_in[8][59] , \add_in[8][58] , \add_in[8][57] , \add_in[8][56] , 
        \add_in[8][55] , \add_in[8][54] , \add_in[8][53] , \add_in[8][52] , 
        \add_in[8][51] , \add_in[8][50] , \add_in[8][49] , \add_in[8][48] , 
        \add_in[8][47] , \add_in[8][46] , \add_in[8][45] , \add_in[8][44] , 
        \add_in[8][43] , \add_in[8][42] , \add_in[8][41] , \add_in[8][40] , 
        \add_in[8][39] , \add_in[8][38] , \add_in[8][37] , \add_in[8][36] , 
        \add_in[8][35] , \add_in[8][34] , \add_in[8][33] , \add_in[8][32] , 
        \add_in[8][31] , \add_in[8][30] , \add_in[8][29] , \add_in[8][28] , 
        \add_in[8][27] , \add_in[8][26] , \add_in[8][25] , \add_in[8][24] , 
        \add_in[8][23] , \add_in[8][22] , \add_in[8][21] , \add_in[8][20] , 
        \add_in[8][19] , \add_in[8][18] , \add_in[8][17] , \add_in[8][16] , 
        \add_in[8][15] , \add_in[8][14] , \add_in[8][13] , \add_in[8][12] , 
        \add_in[8][11] , \add_in[8][10] , \add_in[8][9] , \add_in[8][8] , 
        \add_in[8][7] , \add_in[8][6] , \add_in[8][5] , \add_in[8][4] , 
        \add_in[8][3] , \add_in[8][2] , \add_in[8][1] , \add_in[8][0] }) );
  RCA_generic_N64_7 add_i_8 ( .A({\mux_out[9][63] , \mux_out[9][62] , 
        \mux_out[9][61] , \mux_out[9][60] , \mux_out[9][59] , \mux_out[9][58] , 
        \mux_out[9][57] , \mux_out[9][56] , \mux_out[9][55] , \mux_out[9][54] , 
        \mux_out[9][53] , \mux_out[9][52] , \mux_out[9][51] , \mux_out[9][50] , 
        \mux_out[9][49] , \mux_out[9][48] , \mux_out[9][47] , \mux_out[9][46] , 
        \mux_out[9][45] , \mux_out[9][44] , \mux_out[9][43] , \mux_out[9][42] , 
        \mux_out[9][41] , \mux_out[9][40] , \mux_out[9][39] , \mux_out[9][38] , 
        \mux_out[9][37] , \mux_out[9][36] , \mux_out[9][35] , \mux_out[9][34] , 
        \mux_out[9][33] , \mux_out[9][32] , \mux_out[9][31] , \mux_out[9][30] , 
        \mux_out[9][29] , \mux_out[9][28] , \mux_out[9][27] , \mux_out[9][26] , 
        \mux_out[9][25] , \mux_out[9][24] , \mux_out[9][23] , \mux_out[9][22] , 
        \mux_out[9][21] , \mux_out[9][20] , \mux_out[9][19] , \mux_out[9][18] , 
        \mux_out[9][17] , \mux_out[9][16] , \mux_out[9][15] , \mux_out[9][14] , 
        \mux_out[9][13] , \mux_out[9][12] , \mux_out[9][11] , \mux_out[9][10] , 
        \mux_out[9][9] , \mux_out[9][8] , \mux_out[9][7] , \mux_out[9][6] , 
        \mux_out[9][5] , \mux_out[9][4] , \mux_out[9][3] , \mux_out[9][2] , 
        \mux_out[9][1] , \mux_out[9][0] }), .B({\add_in[8][63] , 
        \add_in[8][62] , \add_in[8][61] , \add_in[8][60] , \add_in[8][59] , 
        \add_in[8][58] , \add_in[8][57] , \add_in[8][56] , \add_in[8][55] , 
        \add_in[8][54] , \add_in[8][53] , \add_in[8][52] , \add_in[8][51] , 
        \add_in[8][50] , \add_in[8][49] , \add_in[8][48] , \add_in[8][47] , 
        \add_in[8][46] , \add_in[8][45] , \add_in[8][44] , \add_in[8][43] , 
        \add_in[8][42] , \add_in[8][41] , \add_in[8][40] , \add_in[8][39] , 
        \add_in[8][38] , \add_in[8][37] , \add_in[8][36] , \add_in[8][35] , 
        \add_in[8][34] , \add_in[8][33] , \add_in[8][32] , \add_in[8][31] , 
        \add_in[8][30] , \add_in[8][29] , \add_in[8][28] , \add_in[8][27] , 
        \add_in[8][26] , \add_in[8][25] , \add_in[8][24] , \add_in[8][23] , 
        \add_in[8][22] , \add_in[8][21] , \add_in[8][20] , \add_in[8][19] , 
        \add_in[8][18] , \add_in[8][17] , \add_in[8][16] , \add_in[8][15] , 
        \add_in[8][14] , \add_in[8][13] , \add_in[8][12] , \add_in[8][11] , 
        \add_in[8][10] , \add_in[8][9] , \add_in[8][8] , \add_in[8][7] , 
        \add_in[8][6] , \add_in[8][5] , \add_in[8][4] , \add_in[8][3] , 
        \add_in[8][2] , \add_in[8][1] , \add_in[8][0] }), .Ci(mode[8]), .S({
        \add_in[9][63] , \add_in[9][62] , \add_in[9][61] , \add_in[9][60] , 
        \add_in[9][59] , \add_in[9][58] , \add_in[9][57] , \add_in[9][56] , 
        \add_in[9][55] , \add_in[9][54] , \add_in[9][53] , \add_in[9][52] , 
        \add_in[9][51] , \add_in[9][50] , \add_in[9][49] , \add_in[9][48] , 
        \add_in[9][47] , \add_in[9][46] , \add_in[9][45] , \add_in[9][44] , 
        \add_in[9][43] , \add_in[9][42] , \add_in[9][41] , \add_in[9][40] , 
        \add_in[9][39] , \add_in[9][38] , \add_in[9][37] , \add_in[9][36] , 
        \add_in[9][35] , \add_in[9][34] , \add_in[9][33] , \add_in[9][32] , 
        \add_in[9][31] , \add_in[9][30] , \add_in[9][29] , \add_in[9][28] , 
        \add_in[9][27] , \add_in[9][26] , \add_in[9][25] , \add_in[9][24] , 
        \add_in[9][23] , \add_in[9][22] , \add_in[9][21] , \add_in[9][20] , 
        \add_in[9][19] , \add_in[9][18] , \add_in[9][17] , \add_in[9][16] , 
        \add_in[9][15] , \add_in[9][14] , \add_in[9][13] , \add_in[9][12] , 
        \add_in[9][11] , \add_in[9][10] , \add_in[9][9] , \add_in[9][8] , 
        \add_in[9][7] , \add_in[9][6] , \add_in[9][5] , \add_in[9][4] , 
        \add_in[9][3] , \add_in[9][2] , \add_in[9][1] , \add_in[9][0] }) );
  RCA_generic_N64_6 add_i_9 ( .A({\mux_out[10][63] , \mux_out[10][62] , 
        \mux_out[10][61] , \mux_out[10][60] , \mux_out[10][59] , 
        \mux_out[10][58] , \mux_out[10][57] , \mux_out[10][56] , 
        \mux_out[10][55] , \mux_out[10][54] , \mux_out[10][53] , 
        \mux_out[10][52] , \mux_out[10][51] , \mux_out[10][50] , 
        \mux_out[10][49] , \mux_out[10][48] , \mux_out[10][47] , 
        \mux_out[10][46] , \mux_out[10][45] , \mux_out[10][44] , 
        \mux_out[10][43] , \mux_out[10][42] , \mux_out[10][41] , 
        \mux_out[10][40] , \mux_out[10][39] , \mux_out[10][38] , 
        \mux_out[10][37] , \mux_out[10][36] , \mux_out[10][35] , 
        \mux_out[10][34] , \mux_out[10][33] , \mux_out[10][32] , 
        \mux_out[10][31] , \mux_out[10][30] , \mux_out[10][29] , 
        \mux_out[10][28] , \mux_out[10][27] , \mux_out[10][26] , 
        \mux_out[10][25] , \mux_out[10][24] , \mux_out[10][23] , 
        \mux_out[10][22] , \mux_out[10][21] , \mux_out[10][20] , 
        \mux_out[10][19] , \mux_out[10][18] , \mux_out[10][17] , 
        \mux_out[10][16] , \mux_out[10][15] , \mux_out[10][14] , 
        \mux_out[10][13] , \mux_out[10][12] , \mux_out[10][11] , 
        \mux_out[10][10] , \mux_out[10][9] , \mux_out[10][8] , 
        \mux_out[10][7] , \mux_out[10][6] , \mux_out[10][5] , \mux_out[10][4] , 
        \mux_out[10][3] , \mux_out[10][2] , \mux_out[10][1] , \mux_out[10][0] }), .B({\add_in[9][63] , \add_in[9][62] , \add_in[9][61] , \add_in[9][60] , 
        \add_in[9][59] , \add_in[9][58] , \add_in[9][57] , \add_in[9][56] , 
        \add_in[9][55] , \add_in[9][54] , \add_in[9][53] , \add_in[9][52] , 
        \add_in[9][51] , \add_in[9][50] , \add_in[9][49] , \add_in[9][48] , 
        \add_in[9][47] , \add_in[9][46] , \add_in[9][45] , \add_in[9][44] , 
        \add_in[9][43] , \add_in[9][42] , \add_in[9][41] , \add_in[9][40] , 
        \add_in[9][39] , \add_in[9][38] , \add_in[9][37] , \add_in[9][36] , 
        \add_in[9][35] , \add_in[9][34] , \add_in[9][33] , \add_in[9][32] , 
        \add_in[9][31] , \add_in[9][30] , \add_in[9][29] , \add_in[9][28] , 
        \add_in[9][27] , \add_in[9][26] , \add_in[9][25] , \add_in[9][24] , 
        \add_in[9][23] , \add_in[9][22] , \add_in[9][21] , \add_in[9][20] , 
        \add_in[9][19] , \add_in[9][18] , \add_in[9][17] , \add_in[9][16] , 
        \add_in[9][15] , \add_in[9][14] , \add_in[9][13] , \add_in[9][12] , 
        \add_in[9][11] , \add_in[9][10] , \add_in[9][9] , \add_in[9][8] , 
        \add_in[9][7] , \add_in[9][6] , \add_in[9][5] , \add_in[9][4] , 
        \add_in[9][3] , \add_in[9][2] , \add_in[9][1] , \add_in[9][0] }), .Ci(
        mode[9]), .S({\add_in[10][63] , \add_in[10][62] , \add_in[10][61] , 
        \add_in[10][60] , \add_in[10][59] , \add_in[10][58] , \add_in[10][57] , 
        \add_in[10][56] , \add_in[10][55] , \add_in[10][54] , \add_in[10][53] , 
        \add_in[10][52] , \add_in[10][51] , \add_in[10][50] , \add_in[10][49] , 
        \add_in[10][48] , \add_in[10][47] , \add_in[10][46] , \add_in[10][45] , 
        \add_in[10][44] , \add_in[10][43] , \add_in[10][42] , \add_in[10][41] , 
        \add_in[10][40] , \add_in[10][39] , \add_in[10][38] , \add_in[10][37] , 
        \add_in[10][36] , \add_in[10][35] , \add_in[10][34] , \add_in[10][33] , 
        \add_in[10][32] , \add_in[10][31] , \add_in[10][30] , \add_in[10][29] , 
        \add_in[10][28] , \add_in[10][27] , \add_in[10][26] , \add_in[10][25] , 
        \add_in[10][24] , \add_in[10][23] , \add_in[10][22] , \add_in[10][21] , 
        \add_in[10][20] , \add_in[10][19] , \add_in[10][18] , \add_in[10][17] , 
        \add_in[10][16] , \add_in[10][15] , \add_in[10][14] , \add_in[10][13] , 
        \add_in[10][12] , \add_in[10][11] , \add_in[10][10] , \add_in[10][9] , 
        \add_in[10][8] , \add_in[10][7] , \add_in[10][6] , \add_in[10][5] , 
        \add_in[10][4] , \add_in[10][3] , \add_in[10][2] , \add_in[10][1] , 
        \add_in[10][0] }) );
  RCA_generic_N64_5 add_i_10 ( .A({\mux_out[11][63] , \mux_out[11][62] , 
        \mux_out[11][61] , \mux_out[11][60] , \mux_out[11][59] , 
        \mux_out[11][58] , \mux_out[11][57] , \mux_out[11][56] , 
        \mux_out[11][55] , \mux_out[11][54] , \mux_out[11][53] , 
        \mux_out[11][52] , \mux_out[11][51] , \mux_out[11][50] , 
        \mux_out[11][49] , \mux_out[11][48] , \mux_out[11][47] , 
        \mux_out[11][46] , \mux_out[11][45] , \mux_out[11][44] , 
        \mux_out[11][43] , \mux_out[11][42] , \mux_out[11][41] , 
        \mux_out[11][40] , \mux_out[11][39] , \mux_out[11][38] , 
        \mux_out[11][37] , \mux_out[11][36] , \mux_out[11][35] , 
        \mux_out[11][34] , \mux_out[11][33] , \mux_out[11][32] , 
        \mux_out[11][31] , \mux_out[11][30] , \mux_out[11][29] , 
        \mux_out[11][28] , \mux_out[11][27] , \mux_out[11][26] , 
        \mux_out[11][25] , \mux_out[11][24] , \mux_out[11][23] , 
        \mux_out[11][22] , \mux_out[11][21] , \mux_out[11][20] , 
        \mux_out[11][19] , \mux_out[11][18] , \mux_out[11][17] , 
        \mux_out[11][16] , \mux_out[11][15] , \mux_out[11][14] , 
        \mux_out[11][13] , \mux_out[11][12] , \mux_out[11][11] , 
        \mux_out[11][10] , \mux_out[11][9] , \mux_out[11][8] , 
        \mux_out[11][7] , \mux_out[11][6] , \mux_out[11][5] , \mux_out[11][4] , 
        \mux_out[11][3] , \mux_out[11][2] , \mux_out[11][1] , \mux_out[11][0] }), .B({\add_in[10][63] , \add_in[10][62] , \add_in[10][61] , \add_in[10][60] , 
        \add_in[10][59] , \add_in[10][58] , \add_in[10][57] , \add_in[10][56] , 
        \add_in[10][55] , \add_in[10][54] , \add_in[10][53] , \add_in[10][52] , 
        \add_in[10][51] , \add_in[10][50] , \add_in[10][49] , \add_in[10][48] , 
        \add_in[10][47] , \add_in[10][46] , \add_in[10][45] , \add_in[10][44] , 
        \add_in[10][43] , \add_in[10][42] , \add_in[10][41] , \add_in[10][40] , 
        \add_in[10][39] , \add_in[10][38] , \add_in[10][37] , \add_in[10][36] , 
        \add_in[10][35] , \add_in[10][34] , \add_in[10][33] , \add_in[10][32] , 
        \add_in[10][31] , \add_in[10][30] , \add_in[10][29] , \add_in[10][28] , 
        \add_in[10][27] , \add_in[10][26] , \add_in[10][25] , \add_in[10][24] , 
        \add_in[10][23] , \add_in[10][22] , \add_in[10][21] , \add_in[10][20] , 
        \add_in[10][19] , \add_in[10][18] , \add_in[10][17] , \add_in[10][16] , 
        \add_in[10][15] , \add_in[10][14] , \add_in[10][13] , \add_in[10][12] , 
        \add_in[10][11] , \add_in[10][10] , \add_in[10][9] , \add_in[10][8] , 
        \add_in[10][7] , \add_in[10][6] , \add_in[10][5] , \add_in[10][4] , 
        \add_in[10][3] , \add_in[10][2] , \add_in[10][1] , \add_in[10][0] }), 
        .Ci(mode[10]), .S({\add_in[11][63] , \add_in[11][62] , 
        \add_in[11][61] , \add_in[11][60] , \add_in[11][59] , \add_in[11][58] , 
        \add_in[11][57] , \add_in[11][56] , \add_in[11][55] , \add_in[11][54] , 
        \add_in[11][53] , \add_in[11][52] , \add_in[11][51] , \add_in[11][50] , 
        \add_in[11][49] , \add_in[11][48] , \add_in[11][47] , \add_in[11][46] , 
        \add_in[11][45] , \add_in[11][44] , \add_in[11][43] , \add_in[11][42] , 
        \add_in[11][41] , \add_in[11][40] , \add_in[11][39] , \add_in[11][38] , 
        \add_in[11][37] , \add_in[11][36] , \add_in[11][35] , \add_in[11][34] , 
        \add_in[11][33] , \add_in[11][32] , \add_in[11][31] , \add_in[11][30] , 
        \add_in[11][29] , \add_in[11][28] , \add_in[11][27] , \add_in[11][26] , 
        \add_in[11][25] , \add_in[11][24] , \add_in[11][23] , \add_in[11][22] , 
        \add_in[11][21] , \add_in[11][20] , \add_in[11][19] , \add_in[11][18] , 
        \add_in[11][17] , \add_in[11][16] , \add_in[11][15] , \add_in[11][14] , 
        \add_in[11][13] , \add_in[11][12] , \add_in[11][11] , \add_in[11][10] , 
        \add_in[11][9] , \add_in[11][8] , \add_in[11][7] , \add_in[11][6] , 
        \add_in[11][5] , \add_in[11][4] , \add_in[11][3] , \add_in[11][2] , 
        \add_in[11][1] , \add_in[11][0] }) );
  RCA_generic_N64_4 add_i_11 ( .A({\mux_out[12][63] , \mux_out[12][62] , 
        \mux_out[12][61] , \mux_out[12][60] , \mux_out[12][59] , 
        \mux_out[12][58] , \mux_out[12][57] , \mux_out[12][56] , 
        \mux_out[12][55] , \mux_out[12][54] , \mux_out[12][53] , 
        \mux_out[12][52] , \mux_out[12][51] , \mux_out[12][50] , 
        \mux_out[12][49] , \mux_out[12][48] , \mux_out[12][47] , 
        \mux_out[12][46] , \mux_out[12][45] , \mux_out[12][44] , 
        \mux_out[12][43] , \mux_out[12][42] , \mux_out[12][41] , 
        \mux_out[12][40] , \mux_out[12][39] , \mux_out[12][38] , 
        \mux_out[12][37] , \mux_out[12][36] , \mux_out[12][35] , 
        \mux_out[12][34] , \mux_out[12][33] , \mux_out[12][32] , 
        \mux_out[12][31] , \mux_out[12][30] , \mux_out[12][29] , 
        \mux_out[12][28] , \mux_out[12][27] , \mux_out[12][26] , 
        \mux_out[12][25] , \mux_out[12][24] , \mux_out[12][23] , 
        \mux_out[12][22] , \mux_out[12][21] , \mux_out[12][20] , 
        \mux_out[12][19] , \mux_out[12][18] , \mux_out[12][17] , 
        \mux_out[12][16] , \mux_out[12][15] , \mux_out[12][14] , 
        \mux_out[12][13] , \mux_out[12][12] , \mux_out[12][11] , 
        \mux_out[12][10] , \mux_out[12][9] , \mux_out[12][8] , 
        \mux_out[12][7] , \mux_out[12][6] , \mux_out[12][5] , \mux_out[12][4] , 
        \mux_out[12][3] , \mux_out[12][2] , \mux_out[12][1] , \mux_out[12][0] }), .B({\add_in[11][63] , \add_in[11][62] , \add_in[11][61] , \add_in[11][60] , 
        \add_in[11][59] , \add_in[11][58] , \add_in[11][57] , \add_in[11][56] , 
        \add_in[11][55] , \add_in[11][54] , \add_in[11][53] , \add_in[11][52] , 
        \add_in[11][51] , \add_in[11][50] , \add_in[11][49] , \add_in[11][48] , 
        \add_in[11][47] , \add_in[11][46] , \add_in[11][45] , \add_in[11][44] , 
        \add_in[11][43] , \add_in[11][42] , \add_in[11][41] , \add_in[11][40] , 
        \add_in[11][39] , \add_in[11][38] , \add_in[11][37] , \add_in[11][36] , 
        \add_in[11][35] , \add_in[11][34] , \add_in[11][33] , \add_in[11][32] , 
        \add_in[11][31] , \add_in[11][30] , \add_in[11][29] , \add_in[11][28] , 
        \add_in[11][27] , \add_in[11][26] , \add_in[11][25] , \add_in[11][24] , 
        \add_in[11][23] , \add_in[11][22] , \add_in[11][21] , \add_in[11][20] , 
        \add_in[11][19] , \add_in[11][18] , \add_in[11][17] , \add_in[11][16] , 
        \add_in[11][15] , \add_in[11][14] , \add_in[11][13] , \add_in[11][12] , 
        \add_in[11][11] , \add_in[11][10] , \add_in[11][9] , \add_in[11][8] , 
        \add_in[11][7] , \add_in[11][6] , \add_in[11][5] , \add_in[11][4] , 
        \add_in[11][3] , \add_in[11][2] , \add_in[11][1] , \add_in[11][0] }), 
        .Ci(mode[11]), .S({\add_in[12][63] , \add_in[12][62] , 
        \add_in[12][61] , \add_in[12][60] , \add_in[12][59] , \add_in[12][58] , 
        \add_in[12][57] , \add_in[12][56] , \add_in[12][55] , \add_in[12][54] , 
        \add_in[12][53] , \add_in[12][52] , \add_in[12][51] , \add_in[12][50] , 
        \add_in[12][49] , \add_in[12][48] , \add_in[12][47] , \add_in[12][46] , 
        \add_in[12][45] , \add_in[12][44] , \add_in[12][43] , \add_in[12][42] , 
        \add_in[12][41] , \add_in[12][40] , \add_in[12][39] , \add_in[12][38] , 
        \add_in[12][37] , \add_in[12][36] , \add_in[12][35] , \add_in[12][34] , 
        \add_in[12][33] , \add_in[12][32] , \add_in[12][31] , \add_in[12][30] , 
        \add_in[12][29] , \add_in[12][28] , \add_in[12][27] , \add_in[12][26] , 
        \add_in[12][25] , \add_in[12][24] , \add_in[12][23] , \add_in[12][22] , 
        \add_in[12][21] , \add_in[12][20] , \add_in[12][19] , \add_in[12][18] , 
        \add_in[12][17] , \add_in[12][16] , \add_in[12][15] , \add_in[12][14] , 
        \add_in[12][13] , \add_in[12][12] , \add_in[12][11] , \add_in[12][10] , 
        \add_in[12][9] , \add_in[12][8] , \add_in[12][7] , \add_in[12][6] , 
        \add_in[12][5] , \add_in[12][4] , \add_in[12][3] , \add_in[12][2] , 
        \add_in[12][1] , \add_in[12][0] }) );
  RCA_generic_N64_3 add_i_12 ( .A({\mux_out[13][63] , \mux_out[13][62] , 
        \mux_out[13][61] , \mux_out[13][60] , \mux_out[13][59] , 
        \mux_out[13][58] , \mux_out[13][57] , \mux_out[13][56] , 
        \mux_out[13][55] , \mux_out[13][54] , \mux_out[13][53] , 
        \mux_out[13][52] , \mux_out[13][51] , \mux_out[13][50] , 
        \mux_out[13][49] , \mux_out[13][48] , \mux_out[13][47] , 
        \mux_out[13][46] , \mux_out[13][45] , \mux_out[13][44] , 
        \mux_out[13][43] , \mux_out[13][42] , \mux_out[13][41] , 
        \mux_out[13][40] , \mux_out[13][39] , \mux_out[13][38] , 
        \mux_out[13][37] , \mux_out[13][36] , \mux_out[13][35] , 
        \mux_out[13][34] , \mux_out[13][33] , \mux_out[13][32] , 
        \mux_out[13][31] , \mux_out[13][30] , \mux_out[13][29] , 
        \mux_out[13][28] , \mux_out[13][27] , \mux_out[13][26] , 
        \mux_out[13][25] , \mux_out[13][24] , \mux_out[13][23] , 
        \mux_out[13][22] , \mux_out[13][21] , \mux_out[13][20] , 
        \mux_out[13][19] , \mux_out[13][18] , \mux_out[13][17] , 
        \mux_out[13][16] , \mux_out[13][15] , \mux_out[13][14] , 
        \mux_out[13][13] , \mux_out[13][12] , \mux_out[13][11] , 
        \mux_out[13][10] , \mux_out[13][9] , \mux_out[13][8] , 
        \mux_out[13][7] , \mux_out[13][6] , \mux_out[13][5] , \mux_out[13][4] , 
        \mux_out[13][3] , \mux_out[13][2] , \mux_out[13][1] , \mux_out[13][0] }), .B({\add_in[12][63] , \add_in[12][62] , \add_in[12][61] , \add_in[12][60] , 
        \add_in[12][59] , \add_in[12][58] , \add_in[12][57] , \add_in[12][56] , 
        \add_in[12][55] , \add_in[12][54] , \add_in[12][53] , \add_in[12][52] , 
        \add_in[12][51] , \add_in[12][50] , \add_in[12][49] , \add_in[12][48] , 
        \add_in[12][47] , \add_in[12][46] , \add_in[12][45] , \add_in[12][44] , 
        \add_in[12][43] , \add_in[12][42] , \add_in[12][41] , \add_in[12][40] , 
        \add_in[12][39] , \add_in[12][38] , \add_in[12][37] , \add_in[12][36] , 
        \add_in[12][35] , \add_in[12][34] , \add_in[12][33] , \add_in[12][32] , 
        \add_in[12][31] , \add_in[12][30] , \add_in[12][29] , \add_in[12][28] , 
        \add_in[12][27] , \add_in[12][26] , \add_in[12][25] , \add_in[12][24] , 
        \add_in[12][23] , \add_in[12][22] , \add_in[12][21] , \add_in[12][20] , 
        \add_in[12][19] , \add_in[12][18] , \add_in[12][17] , \add_in[12][16] , 
        \add_in[12][15] , \add_in[12][14] , \add_in[12][13] , \add_in[12][12] , 
        \add_in[12][11] , \add_in[12][10] , \add_in[12][9] , \add_in[12][8] , 
        \add_in[12][7] , \add_in[12][6] , \add_in[12][5] , \add_in[12][4] , 
        \add_in[12][3] , \add_in[12][2] , \add_in[12][1] , \add_in[12][0] }), 
        .Ci(mode[12]), .S({\add_in[13][63] , \add_in[13][62] , 
        \add_in[13][61] , \add_in[13][60] , \add_in[13][59] , \add_in[13][58] , 
        \add_in[13][57] , \add_in[13][56] , \add_in[13][55] , \add_in[13][54] , 
        \add_in[13][53] , \add_in[13][52] , \add_in[13][51] , \add_in[13][50] , 
        \add_in[13][49] , \add_in[13][48] , \add_in[13][47] , \add_in[13][46] , 
        \add_in[13][45] , \add_in[13][44] , \add_in[13][43] , \add_in[13][42] , 
        \add_in[13][41] , \add_in[13][40] , \add_in[13][39] , \add_in[13][38] , 
        \add_in[13][37] , \add_in[13][36] , \add_in[13][35] , \add_in[13][34] , 
        \add_in[13][33] , \add_in[13][32] , \add_in[13][31] , \add_in[13][30] , 
        \add_in[13][29] , \add_in[13][28] , \add_in[13][27] , \add_in[13][26] , 
        \add_in[13][25] , \add_in[13][24] , \add_in[13][23] , \add_in[13][22] , 
        \add_in[13][21] , \add_in[13][20] , \add_in[13][19] , \add_in[13][18] , 
        \add_in[13][17] , \add_in[13][16] , \add_in[13][15] , \add_in[13][14] , 
        \add_in[13][13] , \add_in[13][12] , \add_in[13][11] , \add_in[13][10] , 
        \add_in[13][9] , \add_in[13][8] , \add_in[13][7] , \add_in[13][6] , 
        \add_in[13][5] , \add_in[13][4] , \add_in[13][3] , \add_in[13][2] , 
        \add_in[13][1] , \add_in[13][0] }) );
  RCA_generic_N64_2 add_i_13 ( .A({\mux_out[14][63] , \mux_out[14][62] , 
        \mux_out[14][61] , \mux_out[14][60] , \mux_out[14][59] , 
        \mux_out[14][58] , \mux_out[14][57] , \mux_out[14][56] , 
        \mux_out[14][55] , \mux_out[14][54] , \mux_out[14][53] , 
        \mux_out[14][52] , \mux_out[14][51] , \mux_out[14][50] , 
        \mux_out[14][49] , \mux_out[14][48] , \mux_out[14][47] , 
        \mux_out[14][46] , \mux_out[14][45] , \mux_out[14][44] , 
        \mux_out[14][43] , \mux_out[14][42] , \mux_out[14][41] , 
        \mux_out[14][40] , \mux_out[14][39] , \mux_out[14][38] , 
        \mux_out[14][37] , \mux_out[14][36] , \mux_out[14][35] , 
        \mux_out[14][34] , \mux_out[14][33] , \mux_out[14][32] , 
        \mux_out[14][31] , \mux_out[14][30] , \mux_out[14][29] , 
        \mux_out[14][28] , \mux_out[14][27] , \mux_out[14][26] , 
        \mux_out[14][25] , \mux_out[14][24] , \mux_out[14][23] , 
        \mux_out[14][22] , \mux_out[14][21] , \mux_out[14][20] , 
        \mux_out[14][19] , \mux_out[14][18] , \mux_out[14][17] , 
        \mux_out[14][16] , \mux_out[14][15] , \mux_out[14][14] , 
        \mux_out[14][13] , \mux_out[14][12] , \mux_out[14][11] , 
        \mux_out[14][10] , \mux_out[14][9] , \mux_out[14][8] , 
        \mux_out[14][7] , \mux_out[14][6] , \mux_out[14][5] , \mux_out[14][4] , 
        \mux_out[14][3] , \mux_out[14][2] , \mux_out[14][1] , \mux_out[14][0] }), .B({\add_in[13][63] , \add_in[13][62] , \add_in[13][61] , \add_in[13][60] , 
        \add_in[13][59] , \add_in[13][58] , \add_in[13][57] , \add_in[13][56] , 
        \add_in[13][55] , \add_in[13][54] , \add_in[13][53] , \add_in[13][52] , 
        \add_in[13][51] , \add_in[13][50] , \add_in[13][49] , \add_in[13][48] , 
        \add_in[13][47] , \add_in[13][46] , \add_in[13][45] , \add_in[13][44] , 
        \add_in[13][43] , \add_in[13][42] , \add_in[13][41] , \add_in[13][40] , 
        \add_in[13][39] , \add_in[13][38] , \add_in[13][37] , \add_in[13][36] , 
        \add_in[13][35] , \add_in[13][34] , \add_in[13][33] , \add_in[13][32] , 
        \add_in[13][31] , \add_in[13][30] , \add_in[13][29] , \add_in[13][28] , 
        \add_in[13][27] , \add_in[13][26] , \add_in[13][25] , \add_in[13][24] , 
        \add_in[13][23] , \add_in[13][22] , \add_in[13][21] , \add_in[13][20] , 
        \add_in[13][19] , \add_in[13][18] , \add_in[13][17] , \add_in[13][16] , 
        \add_in[13][15] , \add_in[13][14] , \add_in[13][13] , \add_in[13][12] , 
        \add_in[13][11] , \add_in[13][10] , \add_in[13][9] , \add_in[13][8] , 
        \add_in[13][7] , \add_in[13][6] , \add_in[13][5] , \add_in[13][4] , 
        \add_in[13][3] , \add_in[13][2] , \add_in[13][1] , \add_in[13][0] }), 
        .Ci(mode[13]), .S({\add_in[14][63] , \add_in[14][62] , 
        \add_in[14][61] , \add_in[14][60] , \add_in[14][59] , \add_in[14][58] , 
        \add_in[14][57] , \add_in[14][56] , \add_in[14][55] , \add_in[14][54] , 
        \add_in[14][53] , \add_in[14][52] , \add_in[14][51] , \add_in[14][50] , 
        \add_in[14][49] , \add_in[14][48] , \add_in[14][47] , \add_in[14][46] , 
        \add_in[14][45] , \add_in[14][44] , \add_in[14][43] , \add_in[14][42] , 
        \add_in[14][41] , \add_in[14][40] , \add_in[14][39] , \add_in[14][38] , 
        \add_in[14][37] , \add_in[14][36] , \add_in[14][35] , \add_in[14][34] , 
        \add_in[14][33] , \add_in[14][32] , \add_in[14][31] , \add_in[14][30] , 
        \add_in[14][29] , \add_in[14][28] , \add_in[14][27] , \add_in[14][26] , 
        \add_in[14][25] , \add_in[14][24] , \add_in[14][23] , \add_in[14][22] , 
        \add_in[14][21] , \add_in[14][20] , \add_in[14][19] , \add_in[14][18] , 
        \add_in[14][17] , \add_in[14][16] , \add_in[14][15] , \add_in[14][14] , 
        \add_in[14][13] , \add_in[14][12] , \add_in[14][11] , \add_in[14][10] , 
        \add_in[14][9] , \add_in[14][8] , \add_in[14][7] , \add_in[14][6] , 
        \add_in[14][5] , \add_in[14][4] , \add_in[14][3] , \add_in[14][2] , 
        \add_in[14][1] , \add_in[14][0] }) );
  RCA_generic_N64_1 add_i_14 ( .A({\mux_out[15][63] , \mux_out[15][62] , 
        \mux_out[15][61] , \mux_out[15][60] , \mux_out[15][59] , 
        \mux_out[15][58] , \mux_out[15][57] , \mux_out[15][56] , 
        \mux_out[15][55] , \mux_out[15][54] , \mux_out[15][53] , 
        \mux_out[15][52] , \mux_out[15][51] , \mux_out[15][50] , 
        \mux_out[15][49] , \mux_out[15][48] , \mux_out[15][47] , 
        \mux_out[15][46] , \mux_out[15][45] , \mux_out[15][44] , 
        \mux_out[15][43] , \mux_out[15][42] , \mux_out[15][41] , 
        \mux_out[15][40] , \mux_out[15][39] , \mux_out[15][38] , 
        \mux_out[15][37] , \mux_out[15][36] , \mux_out[15][35] , 
        \mux_out[15][34] , \mux_out[15][33] , \mux_out[15][32] , 
        \mux_out[15][31] , \mux_out[15][30] , \mux_out[15][29] , 
        \mux_out[15][28] , \mux_out[15][27] , \mux_out[15][26] , 
        \mux_out[15][25] , \mux_out[15][24] , \mux_out[15][23] , 
        \mux_out[15][22] , \mux_out[15][21] , \mux_out[15][20] , 
        \mux_out[15][19] , \mux_out[15][18] , \mux_out[15][17] , 
        \mux_out[15][16] , \mux_out[15][15] , \mux_out[15][14] , 
        \mux_out[15][13] , \mux_out[15][12] , \mux_out[15][11] , 
        \mux_out[15][10] , \mux_out[15][9] , \mux_out[15][8] , 
        \mux_out[15][7] , \mux_out[15][6] , \mux_out[15][5] , \mux_out[15][4] , 
        \mux_out[15][3] , \mux_out[15][2] , \mux_out[15][1] , \mux_out[15][0] }), .B({\add_in[14][63] , \add_in[14][62] , \add_in[14][61] , \add_in[14][60] , 
        \add_in[14][59] , \add_in[14][58] , \add_in[14][57] , \add_in[14][56] , 
        \add_in[14][55] , \add_in[14][54] , \add_in[14][53] , \add_in[14][52] , 
        \add_in[14][51] , \add_in[14][50] , \add_in[14][49] , \add_in[14][48] , 
        \add_in[14][47] , \add_in[14][46] , \add_in[14][45] , \add_in[14][44] , 
        \add_in[14][43] , \add_in[14][42] , \add_in[14][41] , \add_in[14][40] , 
        \add_in[14][39] , \add_in[14][38] , \add_in[14][37] , \add_in[14][36] , 
        \add_in[14][35] , \add_in[14][34] , \add_in[14][33] , \add_in[14][32] , 
        \add_in[14][31] , \add_in[14][30] , \add_in[14][29] , \add_in[14][28] , 
        \add_in[14][27] , \add_in[14][26] , \add_in[14][25] , \add_in[14][24] , 
        \add_in[14][23] , \add_in[14][22] , \add_in[14][21] , \add_in[14][20] , 
        \add_in[14][19] , \add_in[14][18] , \add_in[14][17] , \add_in[14][16] , 
        \add_in[14][15] , \add_in[14][14] , \add_in[14][13] , \add_in[14][12] , 
        \add_in[14][11] , \add_in[14][10] , \add_in[14][9] , \add_in[14][8] , 
        \add_in[14][7] , \add_in[14][6] , \add_in[14][5] , \add_in[14][4] , 
        \add_in[14][3] , \add_in[14][2] , \add_in[14][1] , \add_in[14][0] }), 
        .Ci(mode[14]), .S({\add_in[15][63] , \add_in[15][62] , 
        \add_in[15][61] , \add_in[15][60] , \add_in[15][59] , \add_in[15][58] , 
        \add_in[15][57] , \add_in[15][56] , \add_in[15][55] , \add_in[15][54] , 
        \add_in[15][53] , \add_in[15][52] , \add_in[15][51] , \add_in[15][50] , 
        \add_in[15][49] , \add_in[15][48] , \add_in[15][47] , \add_in[15][46] , 
        \add_in[15][45] , \add_in[15][44] , \add_in[15][43] , \add_in[15][42] , 
        \add_in[15][41] , \add_in[15][40] , \add_in[15][39] , \add_in[15][38] , 
        \add_in[15][37] , \add_in[15][36] , \add_in[15][35] , \add_in[15][34] , 
        \add_in[15][33] , \add_in[15][32] , \add_in[15][31] , \add_in[15][30] , 
        \add_in[15][29] , \add_in[15][28] , \add_in[15][27] , \add_in[15][26] , 
        \add_in[15][25] , \add_in[15][24] , \add_in[15][23] , \add_in[15][22] , 
        \add_in[15][21] , \add_in[15][20] , \add_in[15][19] , \add_in[15][18] , 
        \add_in[15][17] , \add_in[15][16] , \add_in[15][15] , \add_in[15][14] , 
        \add_in[15][13] , \add_in[15][12] , \add_in[15][11] , \add_in[15][10] , 
        \add_in[15][9] , \add_in[15][8] , \add_in[15][7] , \add_in[15][6] , 
        \add_in[15][5] , \add_in[15][4] , \add_in[15][3] , \add_in[15][2] , 
        \add_in[15][1] , \add_in[15][0] }) );
  BOOTHMUL_N32_DW01_add_0 add_128 ( .A({\add_in[15][63] , \add_in[15][62] , 
        \add_in[15][61] , \add_in[15][60] , \add_in[15][59] , \add_in[15][58] , 
        \add_in[15][57] , \add_in[15][56] , \add_in[15][55] , \add_in[15][54] , 
        \add_in[15][53] , \add_in[15][52] , \add_in[15][51] , \add_in[15][50] , 
        \add_in[15][49] , \add_in[15][48] , \add_in[15][47] , \add_in[15][46] , 
        \add_in[15][45] , \add_in[15][44] , \add_in[15][43] , \add_in[15][42] , 
        \add_in[15][41] , \add_in[15][40] , \add_in[15][39] , \add_in[15][38] , 
        \add_in[15][37] , \add_in[15][36] , \add_in[15][35] , \add_in[15][34] , 
        \add_in[15][33] , \add_in[15][32] , \add_in[15][31] , \add_in[15][30] , 
        \add_in[15][29] , \add_in[15][28] , \add_in[15][27] , \add_in[15][26] , 
        \add_in[15][25] , \add_in[15][24] , \add_in[15][23] , \add_in[15][22] , 
        \add_in[15][21] , \add_in[15][20] , \add_in[15][19] , \add_in[15][18] , 
        \add_in[15][17] , \add_in[15][16] , \add_in[15][15] , \add_in[15][14] , 
        \add_in[15][13] , \add_in[15][12] , \add_in[15][11] , \add_in[15][10] , 
        \add_in[15][9] , \add_in[15][8] , \add_in[15][7] , \add_in[15][6] , 
        \add_in[15][5] , \add_in[15][4] , \add_in[15][3] , \add_in[15][2] , 
        \add_in[15][1] , \add_in[15][0] }), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, mode[15]}), 
        .CI(1'b0), .SUM(P) );
  BUF_X1 U130 ( .A(n596), .Z(n589) );
  CLKBUF_X1 U131 ( .A(n619), .Z(n521) );
  CLKBUF_X1 U132 ( .A(n622), .Z(n513) );
  CLKBUF_X1 U133 ( .A(n623), .Z(n509) );
  CLKBUF_X1 U134 ( .A(n598), .Z(n585) );
  BUF_X1 U135 ( .A(n596), .Z(n591) );
  BUF_X1 U136 ( .A(n596), .Z(n590) );
  CLKBUF_X1 U137 ( .A(n595), .Z(n594) );
  CLKBUF_X1 U138 ( .A(n610), .Z(n549) );
  CLKBUF_X1 U139 ( .A(n613), .Z(n540) );
  CLKBUF_X1 U140 ( .A(n612), .Z(n543) );
  CLKBUF_X1 U141 ( .A(n615), .Z(n533) );
  CLKBUF_X1 U142 ( .A(n614), .Z(n537) );
  CLKBUF_X1 U143 ( .A(n616), .Z(n530) );
  CLKBUF_X1 U144 ( .A(n609), .Z(n552) );
  CLKBUF_X1 U145 ( .A(n605), .Z(n564) );
  CLKBUF_X1 U146 ( .A(n624), .Z(n623) );
  CLKBUF_X1 U147 ( .A(n632), .Z(n597) );
  CLKBUF_X1 U148 ( .A(n625), .Z(n620) );
  CLKBUF_X1 U149 ( .A(n627), .Z(n612) );
  CLKBUF_X1 U150 ( .A(n629), .Z(n606) );
  BUF_X1 U151 ( .A(n403), .Z(n402) );
  CLKBUF_X1 U152 ( .A(n635), .Z(n625) );
  CLKBUF_X1 U153 ( .A(n634), .Z(n632) );
  CLKBUF_X1 U154 ( .A(n635), .Z(n626) );
  INV_X1 U155 ( .A(n592), .ZN(n654) );
  INV_X1 U156 ( .A(n594), .ZN(n637) );
  INV_X1 U157 ( .A(n591), .ZN(n661) );
  INV_X1 U158 ( .A(n589), .ZN(n674) );
  INV_X1 U159 ( .A(n594), .ZN(n640) );
  INV_X1 U160 ( .A(n594), .ZN(n639) );
  INV_X1 U161 ( .A(n594), .ZN(n638) );
  INV_X1 U162 ( .A(n588), .ZN(n680) );
  INV_X1 U163 ( .A(n593), .ZN(n647) );
  INV_X1 U164 ( .A(n590), .ZN(n668) );
  BUF_X2 U165 ( .A(n595), .Z(n592) );
  BUF_X1 U166 ( .A(n597), .Z(n588) );
  BUF_X1 U167 ( .A(n600), .Z(n578) );
  BUF_X1 U168 ( .A(n618), .Z(n525) );
  BUF_X1 U169 ( .A(n599), .Z(n580) );
  BUF_X1 U170 ( .A(n620), .Z(n517) );
  BUF_X1 U171 ( .A(n598), .Z(n583) );
  BUF_X1 U172 ( .A(n622), .Z(n512) );
  CLKBUF_X1 U173 ( .A(n600), .Z(n579) );
  BUF_X1 U174 ( .A(n623), .Z(n508) );
  CLKBUF_X1 U175 ( .A(n598), .Z(n584) );
  BUF_X1 U176 ( .A(n619), .Z(n520) );
  BUF_X1 U177 ( .A(n621), .Z(n516) );
  BUF_X1 U178 ( .A(n617), .Z(n528) );
  BUF_X1 U179 ( .A(n618), .Z(n524) );
  CLKBUF_X1 U180 ( .A(n595), .Z(n593) );
  BUF_X1 U181 ( .A(n611), .Z(n546) );
  CLKBUF_X1 U182 ( .A(n617), .Z(n526) );
  BUF_X1 U183 ( .A(n614), .Z(n536) );
  CLKBUF_X1 U184 ( .A(n615), .Z(n534) );
  BUF_X1 U185 ( .A(n613), .Z(n539) );
  BUF_X1 U186 ( .A(n616), .Z(n529) );
  CLKBUF_X1 U187 ( .A(n619), .Z(n522) );
  CLKBUF_X1 U188 ( .A(n620), .Z(n518) );
  BUF_X1 U189 ( .A(n610), .Z(n548) );
  CLKBUF_X1 U190 ( .A(n621), .Z(n514) );
  BUF_X1 U191 ( .A(n611), .Z(n545) );
  CLKBUF_X1 U192 ( .A(n599), .Z(n581) );
  CLKBUF_X1 U193 ( .A(n623), .Z(n510) );
  BUF_X1 U194 ( .A(n612), .Z(n542) );
  BUF_X1 U195 ( .A(n615), .Z(n532) );
  CLKBUF_X1 U196 ( .A(n617), .Z(n527) );
  CLKBUF_X1 U197 ( .A(n618), .Z(n523) );
  CLKBUF_X1 U198 ( .A(n597), .Z(n586) );
  CLKBUF_X1 U199 ( .A(n616), .Z(n531) );
  CLKBUF_X1 U200 ( .A(n620), .Z(n519) );
  BUF_X1 U201 ( .A(n614), .Z(n535) );
  CLKBUF_X1 U202 ( .A(n621), .Z(n515) );
  CLKBUF_X1 U203 ( .A(n599), .Z(n582) );
  CLKBUF_X1 U204 ( .A(n622), .Z(n511) );
  CLKBUF_X1 U205 ( .A(n597), .Z(n587) );
  BUF_X1 U206 ( .A(n607), .Z(n557) );
  BUF_X1 U207 ( .A(n606), .Z(n559) );
  BUF_X1 U208 ( .A(n604), .Z(n567) );
  BUF_X1 U209 ( .A(n605), .Z(n563) );
  CLKBUF_X1 U210 ( .A(n605), .Z(n562) );
  BUF_X1 U211 ( .A(n608), .Z(n554) );
  CLKBUF_X1 U212 ( .A(n608), .Z(n555) );
  CLKBUF_X1 U213 ( .A(n606), .Z(n561) );
  CLKBUF_X1 U214 ( .A(n606), .Z(n560) );
  BUF_X1 U215 ( .A(n604), .Z(n565) );
  CLKBUF_X1 U216 ( .A(n610), .Z(n547) );
  CLKBUF_X1 U217 ( .A(n609), .Z(n550) );
  CLKBUF_X1 U218 ( .A(n611), .Z(n544) );
  CLKBUF_X1 U219 ( .A(n607), .Z(n558) );
  CLKBUF_X1 U220 ( .A(n608), .Z(n553) );
  BUF_X1 U221 ( .A(n609), .Z(n551) );
  CLKBUF_X1 U222 ( .A(n612), .Z(n541) );
  CLKBUF_X1 U223 ( .A(n607), .Z(n556) );
  CLKBUF_X1 U224 ( .A(n613), .Z(n538) );
  CLKBUF_X1 U225 ( .A(n604), .Z(n566) );
  BUF_X1 U226 ( .A(n603), .Z(n570) );
  BUF_X1 U227 ( .A(n602), .Z(n571) );
  BUF_X1 U228 ( .A(n603), .Z(n568) );
  CLKBUF_X1 U229 ( .A(n602), .Z(n573) );
  CLKBUF_X1 U230 ( .A(n603), .Z(n569) );
  BUF_X1 U231 ( .A(n601), .Z(n574) );
  CLKBUF_X1 U232 ( .A(n602), .Z(n572) );
  BUF_X1 U233 ( .A(n601), .Z(n575) );
  CLKBUF_X1 U234 ( .A(n601), .Z(n576) );
  CLKBUF_X1 U235 ( .A(n600), .Z(n577) );
  INV_X1 U236 ( .A(n202), .ZN(n205) );
  INV_X1 U237 ( .A(n212), .ZN(n215) );
  INV_X1 U238 ( .A(n222), .ZN(n225) );
  INV_X1 U239 ( .A(n232), .ZN(n235) );
  INV_X1 U240 ( .A(n242), .ZN(n245) );
  INV_X1 U241 ( .A(n252), .ZN(n255) );
  INV_X1 U242 ( .A(n262), .ZN(n265) );
  INV_X1 U243 ( .A(n272), .ZN(n275) );
  INV_X1 U244 ( .A(n282), .ZN(n285) );
  INV_X1 U245 ( .A(n292), .ZN(n295) );
  INV_X1 U246 ( .A(n302), .ZN(n305) );
  INV_X1 U247 ( .A(n312), .ZN(n315) );
  INV_X1 U248 ( .A(n322), .ZN(n325) );
  INV_X1 U249 ( .A(n332), .ZN(n335) );
  INV_X1 U250 ( .A(n202), .ZN(n206) );
  INV_X1 U251 ( .A(n212), .ZN(n216) );
  INV_X1 U252 ( .A(n222), .ZN(n226) );
  INV_X1 U253 ( .A(n232), .ZN(n236) );
  INV_X1 U254 ( .A(n242), .ZN(n246) );
  INV_X1 U255 ( .A(n252), .ZN(n256) );
  INV_X1 U256 ( .A(n262), .ZN(n266) );
  INV_X1 U257 ( .A(n272), .ZN(n276) );
  INV_X1 U258 ( .A(n282), .ZN(n286) );
  INV_X1 U259 ( .A(n292), .ZN(n296) );
  INV_X1 U260 ( .A(n302), .ZN(n306) );
  INV_X1 U261 ( .A(n312), .ZN(n316) );
  INV_X1 U262 ( .A(n322), .ZN(n326) );
  INV_X1 U263 ( .A(n452), .ZN(n455) );
  INV_X1 U264 ( .A(n472), .ZN(n475) );
  INV_X1 U265 ( .A(n462), .ZN(n465) );
  INV_X1 U266 ( .A(n432), .ZN(n435) );
  INV_X1 U267 ( .A(n492), .ZN(n495) );
  INV_X1 U268 ( .A(n482), .ZN(n485) );
  INV_X1 U269 ( .A(n442), .ZN(n445) );
  INV_X1 U270 ( .A(n412), .ZN(n415) );
  INV_X1 U271 ( .A(n422), .ZN(n425) );
  INV_X1 U272 ( .A(n402), .ZN(n405) );
  INV_X1 U273 ( .A(n342), .ZN(n345) );
  INV_X1 U274 ( .A(n352), .ZN(n355) );
  INV_X1 U275 ( .A(n362), .ZN(n365) );
  INV_X1 U276 ( .A(n372), .ZN(n375) );
  INV_X1 U277 ( .A(n382), .ZN(n385) );
  INV_X1 U278 ( .A(n392), .ZN(n395) );
  INV_X1 U279 ( .A(n472), .ZN(n476) );
  INV_X1 U280 ( .A(n462), .ZN(n466) );
  INV_X1 U281 ( .A(n452), .ZN(n456) );
  INV_X1 U282 ( .A(n442), .ZN(n446) );
  INV_X1 U283 ( .A(n432), .ZN(n436) );
  INV_X1 U284 ( .A(n422), .ZN(n426) );
  INV_X1 U285 ( .A(n412), .ZN(n416) );
  INV_X1 U286 ( .A(n402), .ZN(n406) );
  INV_X1 U287 ( .A(n332), .ZN(n336) );
  INV_X1 U288 ( .A(n342), .ZN(n346) );
  INV_X1 U289 ( .A(n352), .ZN(n356) );
  INV_X1 U290 ( .A(n362), .ZN(n366) );
  INV_X1 U291 ( .A(n372), .ZN(n376) );
  INV_X1 U292 ( .A(n382), .ZN(n386) );
  INV_X1 U293 ( .A(n392), .ZN(n396) );
  INV_X1 U294 ( .A(n502), .ZN(n505) );
  INV_X1 U295 ( .A(n502), .ZN(n506) );
  INV_X1 U296 ( .A(n482), .ZN(n486) );
  INV_X1 U297 ( .A(n492), .ZN(n496) );
  BUF_X1 U298 ( .A(n631), .Z(n600) );
  BUF_X1 U299 ( .A(n626), .Z(n617) );
  BUF_X1 U300 ( .A(n625), .Z(n619) );
  BUF_X1 U301 ( .A(n632), .Z(n598) );
  CLKBUF_X1 U302 ( .A(n625), .Z(n618) );
  CLKBUF_X1 U303 ( .A(n632), .Z(n599) );
  CLKBUF_X1 U304 ( .A(n624), .Z(n621) );
  BUF_X1 U305 ( .A(n624), .Z(n622) );
  BUF_X1 U306 ( .A(n633), .Z(n595) );
  CLKBUF_X1 U307 ( .A(n633), .Z(n596) );
  BUF_X1 U308 ( .A(n628), .Z(n610) );
  CLKBUF_X1 U309 ( .A(n628), .Z(n611) );
  CLKBUF_X1 U310 ( .A(n627), .Z(n613) );
  CLKBUF_X1 U311 ( .A(n626), .Z(n615) );
  BUF_X1 U312 ( .A(n627), .Z(n614) );
  CLKBUF_X1 U313 ( .A(n626), .Z(n616) );
  BUF_X1 U314 ( .A(n630), .Z(n605) );
  CLKBUF_X1 U315 ( .A(n630), .Z(n604) );
  CLKBUF_X1 U316 ( .A(n629), .Z(n607) );
  BUF_X1 U317 ( .A(n629), .Z(n608) );
  CLKBUF_X1 U318 ( .A(n628), .Z(n609) );
  CLKBUF_X1 U319 ( .A(n630), .Z(n603) );
  CLKBUF_X1 U320 ( .A(n631), .Z(n602) );
  CLKBUF_X1 U321 ( .A(n631), .Z(n601) );
  BUF_X2 U322 ( .A(n203), .Z(n202) );
  BUF_X2 U323 ( .A(n213), .Z(n212) );
  BUF_X1 U324 ( .A(n223), .Z(n222) );
  BUF_X1 U325 ( .A(n233), .Z(n232) );
  BUF_X1 U326 ( .A(n243), .Z(n242) );
  BUF_X1 U327 ( .A(n253), .Z(n252) );
  BUF_X1 U328 ( .A(n263), .Z(n262) );
  BUF_X1 U329 ( .A(n273), .Z(n272) );
  BUF_X1 U330 ( .A(n283), .Z(n282) );
  BUF_X1 U331 ( .A(n293), .Z(n292) );
  BUF_X1 U332 ( .A(n303), .Z(n302) );
  BUF_X1 U333 ( .A(n313), .Z(n312) );
  BUF_X1 U334 ( .A(n323), .Z(n322) );
  BUF_X1 U335 ( .A(n333), .Z(n332) );
  BUF_X1 U336 ( .A(n204), .Z(n198) );
  BUF_X1 U337 ( .A(n214), .Z(n208) );
  BUF_X1 U338 ( .A(n224), .Z(n218) );
  BUF_X1 U339 ( .A(n234), .Z(n228) );
  BUF_X1 U340 ( .A(n244), .Z(n238) );
  BUF_X1 U341 ( .A(n254), .Z(n248) );
  BUF_X1 U342 ( .A(n264), .Z(n258) );
  BUF_X1 U343 ( .A(n274), .Z(n268) );
  BUF_X1 U344 ( .A(n284), .Z(n278) );
  BUF_X1 U345 ( .A(n294), .Z(n288) );
  BUF_X2 U346 ( .A(n453), .Z(n452) );
  BUF_X2 U347 ( .A(n493), .Z(n492) );
  BUF_X2 U348 ( .A(n473), .Z(n472) );
  BUF_X2 U349 ( .A(n463), .Z(n462) );
  BUF_X2 U350 ( .A(n483), .Z(n482) );
  BUF_X2 U351 ( .A(n433), .Z(n432) );
  BUF_X2 U352 ( .A(n443), .Z(n442) );
  BUF_X2 U353 ( .A(n413), .Z(n412) );
  BUF_X2 U354 ( .A(n423), .Z(n422) );
  BUF_X1 U355 ( .A(n343), .Z(n342) );
  BUF_X1 U356 ( .A(n353), .Z(n352) );
  BUF_X1 U357 ( .A(n363), .Z(n362) );
  BUF_X1 U358 ( .A(n373), .Z(n372) );
  BUF_X1 U359 ( .A(n383), .Z(n382) );
  BUF_X1 U360 ( .A(n393), .Z(n392) );
  BUF_X1 U361 ( .A(n304), .Z(n298) );
  BUF_X1 U362 ( .A(n314), .Z(n308) );
  BUF_X1 U363 ( .A(n324), .Z(n318) );
  CLKBUF_X1 U364 ( .A(n204), .Z(n199) );
  BUF_X1 U365 ( .A(n334), .Z(n328) );
  BUF_X1 U366 ( .A(n344), .Z(n338) );
  CLKBUF_X1 U367 ( .A(n214), .Z(n209) );
  BUF_X1 U368 ( .A(n354), .Z(n348) );
  CLKBUF_X1 U369 ( .A(n224), .Z(n219) );
  BUF_X1 U370 ( .A(n364), .Z(n358) );
  CLKBUF_X1 U371 ( .A(n234), .Z(n229) );
  BUF_X1 U372 ( .A(n374), .Z(n368) );
  CLKBUF_X1 U373 ( .A(n244), .Z(n239) );
  BUF_X1 U374 ( .A(n384), .Z(n378) );
  CLKBUF_X1 U375 ( .A(n254), .Z(n249) );
  BUF_X1 U376 ( .A(n394), .Z(n388) );
  CLKBUF_X1 U377 ( .A(n264), .Z(n259) );
  BUF_X1 U378 ( .A(n404), .Z(n398) );
  CLKBUF_X1 U379 ( .A(n274), .Z(n269) );
  BUF_X1 U380 ( .A(n414), .Z(n408) );
  CLKBUF_X1 U381 ( .A(n284), .Z(n279) );
  BUF_X1 U382 ( .A(n424), .Z(n418) );
  CLKBUF_X1 U383 ( .A(n294), .Z(n289) );
  BUF_X1 U384 ( .A(n434), .Z(n428) );
  CLKBUF_X1 U385 ( .A(n304), .Z(n299) );
  BUF_X1 U386 ( .A(n444), .Z(n438) );
  CLKBUF_X1 U387 ( .A(n314), .Z(n309) );
  BUF_X1 U388 ( .A(n454), .Z(n448) );
  BUF_X2 U389 ( .A(n503), .Z(n502) );
  CLKBUF_X1 U390 ( .A(n203), .Z(n200) );
  CLKBUF_X1 U391 ( .A(n213), .Z(n210) );
  CLKBUF_X1 U392 ( .A(n223), .Z(n220) );
  CLKBUF_X1 U393 ( .A(n233), .Z(n230) );
  CLKBUF_X1 U394 ( .A(n243), .Z(n240) );
  CLKBUF_X1 U395 ( .A(n253), .Z(n250) );
  CLKBUF_X1 U396 ( .A(n263), .Z(n260) );
  CLKBUF_X1 U397 ( .A(n273), .Z(n270) );
  CLKBUF_X1 U398 ( .A(n283), .Z(n280) );
  CLKBUF_X1 U399 ( .A(n293), .Z(n290) );
  CLKBUF_X1 U400 ( .A(n324), .Z(n319) );
  BUF_X1 U401 ( .A(n464), .Z(n458) );
  CLKBUF_X1 U402 ( .A(n334), .Z(n329) );
  BUF_X1 U403 ( .A(n474), .Z(n468) );
  BUF_X1 U404 ( .A(n484), .Z(n478) );
  CLKBUF_X1 U405 ( .A(n344), .Z(n339) );
  BUF_X1 U406 ( .A(n494), .Z(n488) );
  CLKBUF_X1 U407 ( .A(n354), .Z(n349) );
  CLKBUF_X1 U408 ( .A(n364), .Z(n359) );
  BUF_X1 U409 ( .A(n504), .Z(n498) );
  CLKBUF_X1 U410 ( .A(n374), .Z(n369) );
  CLKBUF_X1 U411 ( .A(n384), .Z(n379) );
  CLKBUF_X1 U412 ( .A(n474), .Z(n469) );
  CLKBUF_X1 U413 ( .A(n394), .Z(n389) );
  CLKBUF_X1 U414 ( .A(n404), .Z(n399) );
  CLKBUF_X1 U415 ( .A(n414), .Z(n409) );
  CLKBUF_X1 U416 ( .A(n424), .Z(n419) );
  CLKBUF_X1 U417 ( .A(n434), .Z(n429) );
  CLKBUF_X1 U418 ( .A(n464), .Z(n459) );
  CLKBUF_X1 U419 ( .A(n444), .Z(n439) );
  CLKBUF_X1 U420 ( .A(n454), .Z(n449) );
  CLKBUF_X1 U421 ( .A(n634), .Z(n631) );
  BUF_X1 U422 ( .A(n635), .Z(n624) );
  BUF_X1 U423 ( .A(n634), .Z(n633) );
  CLKBUF_X1 U424 ( .A(n443), .Z(n440) );
  CLKBUF_X1 U425 ( .A(n433), .Z(n430) );
  CLKBUF_X1 U426 ( .A(n423), .Z(n420) );
  CLKBUF_X1 U427 ( .A(n303), .Z(n300) );
  CLKBUF_X1 U428 ( .A(n313), .Z(n310) );
  CLKBUF_X1 U429 ( .A(n323), .Z(n320) );
  CLKBUF_X1 U430 ( .A(n333), .Z(n330) );
  CLKBUF_X1 U431 ( .A(n203), .Z(n201) );
  CLKBUF_X1 U432 ( .A(n343), .Z(n340) );
  CLKBUF_X1 U433 ( .A(n213), .Z(n211) );
  CLKBUF_X1 U434 ( .A(n353), .Z(n350) );
  CLKBUF_X1 U435 ( .A(n223), .Z(n221) );
  CLKBUF_X1 U436 ( .A(n363), .Z(n360) );
  CLKBUF_X1 U437 ( .A(n233), .Z(n231) );
  CLKBUF_X1 U438 ( .A(n373), .Z(n370) );
  CLKBUF_X1 U439 ( .A(n413), .Z(n410) );
  CLKBUF_X1 U440 ( .A(n243), .Z(n241) );
  CLKBUF_X1 U441 ( .A(n383), .Z(n380) );
  CLKBUF_X1 U442 ( .A(n253), .Z(n251) );
  CLKBUF_X1 U443 ( .A(n393), .Z(n390) );
  CLKBUF_X1 U444 ( .A(n263), .Z(n261) );
  CLKBUF_X1 U445 ( .A(n403), .Z(n400) );
  CLKBUF_X1 U446 ( .A(n273), .Z(n271) );
  CLKBUF_X1 U447 ( .A(n283), .Z(n281) );
  CLKBUF_X1 U448 ( .A(n293), .Z(n291) );
  CLKBUF_X1 U449 ( .A(n303), .Z(n301) );
  CLKBUF_X1 U450 ( .A(n504), .Z(n499) );
  CLKBUF_X1 U451 ( .A(n494), .Z(n489) );
  CLKBUF_X1 U452 ( .A(n484), .Z(n479) );
  CLKBUF_X1 U453 ( .A(n635), .Z(n628) );
  CLKBUF_X1 U454 ( .A(n635), .Z(n627) );
  CLKBUF_X1 U455 ( .A(n503), .Z(n500) );
  CLKBUF_X1 U456 ( .A(n463), .Z(n461) );
  CLKBUF_X1 U457 ( .A(n453), .Z(n451) );
  CLKBUF_X1 U458 ( .A(n493), .Z(n490) );
  CLKBUF_X1 U459 ( .A(n443), .Z(n441) );
  CLKBUF_X1 U460 ( .A(n483), .Z(n480) );
  CLKBUF_X1 U461 ( .A(n433), .Z(n431) );
  CLKBUF_X1 U462 ( .A(n473), .Z(n470) );
  CLKBUF_X1 U463 ( .A(n423), .Z(n421) );
  CLKBUF_X1 U464 ( .A(n463), .Z(n460) );
  CLKBUF_X1 U465 ( .A(n453), .Z(n450) );
  CLKBUF_X1 U466 ( .A(n413), .Z(n411) );
  CLKBUF_X1 U467 ( .A(n403), .Z(n401) );
  CLKBUF_X1 U468 ( .A(n393), .Z(n391) );
  CLKBUF_X1 U469 ( .A(n313), .Z(n311) );
  CLKBUF_X1 U470 ( .A(n323), .Z(n321) );
  CLKBUF_X1 U471 ( .A(n333), .Z(n331) );
  CLKBUF_X1 U472 ( .A(n343), .Z(n341) );
  CLKBUF_X1 U473 ( .A(n353), .Z(n351) );
  CLKBUF_X1 U474 ( .A(n363), .Z(n361) );
  CLKBUF_X1 U475 ( .A(n373), .Z(n371) );
  CLKBUF_X1 U476 ( .A(n383), .Z(n381) );
  CLKBUF_X1 U477 ( .A(n634), .Z(n630) );
  CLKBUF_X1 U478 ( .A(n634), .Z(n629) );
  CLKBUF_X1 U479 ( .A(n473), .Z(n471) );
  CLKBUF_X1 U480 ( .A(n483), .Z(n481) );
  CLKBUF_X1 U481 ( .A(n493), .Z(n491) );
  CLKBUF_X1 U482 ( .A(n503), .Z(n501) );
  BUF_X1 U483 ( .A(A[0]), .Z(n203) );
  BUF_X1 U484 ( .A(A[1]), .Z(n213) );
  BUF_X1 U485 ( .A(A[2]), .Z(n223) );
  BUF_X1 U486 ( .A(A[3]), .Z(n233) );
  BUF_X1 U487 ( .A(A[4]), .Z(n243) );
  BUF_X1 U488 ( .A(A[5]), .Z(n253) );
  BUF_X1 U489 ( .A(A[6]), .Z(n263) );
  BUF_X1 U490 ( .A(A[7]), .Z(n273) );
  BUF_X1 U491 ( .A(A[8]), .Z(n283) );
  BUF_X1 U492 ( .A(A[9]), .Z(n293) );
  BUF_X1 U493 ( .A(A[10]), .Z(n303) );
  BUF_X1 U494 ( .A(A[11]), .Z(n313) );
  BUF_X1 U495 ( .A(A[12]), .Z(n323) );
  BUF_X1 U496 ( .A(A[13]), .Z(n333) );
  BUF_X1 U497 ( .A(A[0]), .Z(n204) );
  BUF_X1 U498 ( .A(A[1]), .Z(n214) );
  BUF_X1 U499 ( .A(A[2]), .Z(n224) );
  BUF_X1 U500 ( .A(A[3]), .Z(n234) );
  BUF_X1 U501 ( .A(A[4]), .Z(n244) );
  BUF_X1 U502 ( .A(A[5]), .Z(n254) );
  BUF_X1 U503 ( .A(A[6]), .Z(n264) );
  BUF_X1 U504 ( .A(A[7]), .Z(n274) );
  BUF_X1 U505 ( .A(A[8]), .Z(n284) );
  BUF_X1 U506 ( .A(A[9]), .Z(n294) );
  BUF_X1 U507 ( .A(A[29]), .Z(n493) );
  BUF_X1 U508 ( .A(A[27]), .Z(n473) );
  BUF_X1 U509 ( .A(A[28]), .Z(n483) );
  BUF_X1 U510 ( .A(A[25]), .Z(n453) );
  BUF_X1 U511 ( .A(A[26]), .Z(n463) );
  BUF_X1 U512 ( .A(A[23]), .Z(n433) );
  BUF_X1 U513 ( .A(A[24]), .Z(n443) );
  BUF_X1 U514 ( .A(A[22]), .Z(n423) );
  BUF_X1 U515 ( .A(A[21]), .Z(n413) );
  BUF_X1 U516 ( .A(A[20]), .Z(n403) );
  BUF_X1 U517 ( .A(A[14]), .Z(n343) );
  BUF_X1 U518 ( .A(A[15]), .Z(n353) );
  BUF_X1 U519 ( .A(A[16]), .Z(n363) );
  BUF_X1 U520 ( .A(A[17]), .Z(n373) );
  BUF_X1 U521 ( .A(A[19]), .Z(n393) );
  BUF_X1 U522 ( .A(A[18]), .Z(n383) );
  BUF_X1 U523 ( .A(A[10]), .Z(n304) );
  BUF_X1 U524 ( .A(A[11]), .Z(n314) );
  BUF_X1 U525 ( .A(A[12]), .Z(n324) );
  BUF_X1 U526 ( .A(A[13]), .Z(n334) );
  BUF_X1 U527 ( .A(A[14]), .Z(n344) );
  BUF_X1 U528 ( .A(A[15]), .Z(n354) );
  BUF_X1 U529 ( .A(A[16]), .Z(n364) );
  BUF_X1 U530 ( .A(A[17]), .Z(n374) );
  BUF_X1 U531 ( .A(A[18]), .Z(n384) );
  BUF_X1 U532 ( .A(A[19]), .Z(n394) );
  BUF_X1 U533 ( .A(A[20]), .Z(n404) );
  BUF_X1 U534 ( .A(A[21]), .Z(n414) );
  BUF_X1 U535 ( .A(A[22]), .Z(n424) );
  BUF_X1 U536 ( .A(A[23]), .Z(n434) );
  BUF_X1 U537 ( .A(A[24]), .Z(n444) );
  BUF_X1 U538 ( .A(A[25]), .Z(n454) );
  BUF_X1 U539 ( .A(A[30]), .Z(n503) );
  BUF_X2 U540 ( .A(A[31]), .Z(n634) );
  BUF_X1 U541 ( .A(A[31]), .Z(n635) );
  BUF_X1 U542 ( .A(A[30]), .Z(n504) );
  BUF_X1 U543 ( .A(A[29]), .Z(n494) );
  BUF_X1 U544 ( .A(A[28]), .Z(n484) );
  BUF_X1 U545 ( .A(A[27]), .Z(n474) );
  BUF_X1 U546 ( .A(A[26]), .Z(n464) );
  INV_X1 U547 ( .A(n202), .ZN(n207) );
  INV_X1 U548 ( .A(n212), .ZN(n217) );
  INV_X1 U549 ( .A(n222), .ZN(n227) );
  INV_X1 U550 ( .A(n232), .ZN(n237) );
  INV_X1 U551 ( .A(n242), .ZN(n247) );
  INV_X1 U552 ( .A(n252), .ZN(n257) );
  INV_X1 U553 ( .A(n262), .ZN(n267) );
  INV_X1 U554 ( .A(n272), .ZN(n277) );
  INV_X1 U555 ( .A(n282), .ZN(n287) );
  INV_X1 U556 ( .A(n292), .ZN(n297) );
  INV_X1 U557 ( .A(n302), .ZN(n307) );
  INV_X1 U558 ( .A(n312), .ZN(n317) );
  INV_X1 U559 ( .A(n322), .ZN(n327) );
  INV_X1 U560 ( .A(n332), .ZN(n337) );
  INV_X1 U561 ( .A(n342), .ZN(n347) );
  INV_X1 U562 ( .A(n352), .ZN(n357) );
  INV_X1 U563 ( .A(n362), .ZN(n367) );
  INV_X1 U564 ( .A(n372), .ZN(n377) );
  INV_X1 U565 ( .A(n382), .ZN(n387) );
  INV_X1 U566 ( .A(n392), .ZN(n397) );
  INV_X1 U567 ( .A(n402), .ZN(n407) );
  INV_X1 U568 ( .A(n412), .ZN(n417) );
  INV_X1 U569 ( .A(n422), .ZN(n427) );
  INV_X1 U570 ( .A(n432), .ZN(n437) );
  INV_X1 U571 ( .A(n442), .ZN(n447) );
  INV_X1 U572 ( .A(n452), .ZN(n457) );
  INV_X1 U573 ( .A(n462), .ZN(n467) );
  INV_X1 U574 ( .A(n472), .ZN(n477) );
  INV_X1 U575 ( .A(n482), .ZN(n487) );
  INV_X1 U576 ( .A(n492), .ZN(n497) );
  INV_X1 U577 ( .A(n502), .ZN(n507) );
  INV_X1 U578 ( .A(n594), .ZN(n636) );
  INV_X1 U579 ( .A(n593), .ZN(n641) );
  INV_X1 U580 ( .A(n593), .ZN(n642) );
  INV_X1 U581 ( .A(n593), .ZN(n643) );
  INV_X1 U582 ( .A(n593), .ZN(n644) );
  INV_X1 U583 ( .A(n593), .ZN(n645) );
  INV_X1 U584 ( .A(n593), .ZN(n646) );
  INV_X1 U585 ( .A(n592), .ZN(n648) );
  INV_X1 U586 ( .A(n592), .ZN(n649) );
  INV_X1 U587 ( .A(n592), .ZN(n650) );
  INV_X1 U588 ( .A(n592), .ZN(n651) );
  INV_X1 U589 ( .A(n592), .ZN(n652) );
  INV_X1 U590 ( .A(n592), .ZN(n653) );
  INV_X1 U591 ( .A(n591), .ZN(n655) );
  INV_X1 U592 ( .A(n591), .ZN(n656) );
  INV_X1 U593 ( .A(n591), .ZN(n657) );
  INV_X1 U594 ( .A(n591), .ZN(n658) );
  INV_X1 U595 ( .A(n591), .ZN(n659) );
  INV_X1 U596 ( .A(n591), .ZN(n660) );
  INV_X1 U597 ( .A(n590), .ZN(n662) );
  INV_X1 U598 ( .A(n590), .ZN(n663) );
  INV_X1 U599 ( .A(n590), .ZN(n664) );
  INV_X1 U600 ( .A(n590), .ZN(n665) );
  INV_X1 U601 ( .A(n590), .ZN(n666) );
  INV_X1 U602 ( .A(n590), .ZN(n667) );
  INV_X1 U603 ( .A(n589), .ZN(n669) );
  INV_X1 U604 ( .A(n589), .ZN(n670) );
  INV_X1 U605 ( .A(n589), .ZN(n671) );
  INV_X1 U606 ( .A(n589), .ZN(n672) );
  INV_X1 U607 ( .A(n589), .ZN(n673) );
  INV_X1 U608 ( .A(n588), .ZN(n675) );
  INV_X1 U609 ( .A(n588), .ZN(n676) );
  INV_X1 U610 ( .A(n588), .ZN(n677) );
  INV_X1 U611 ( .A(n588), .ZN(n678) );
  INV_X1 U612 ( .A(n588), .ZN(n679) );
  INV_X1 U613 ( .A(B[29]), .ZN(n681) );
  AOI21_X1 U614 ( .B1(B[28]), .B2(B[27]), .A(n681), .ZN(mode[14]) );
  INV_X1 U615 ( .A(B[27]), .ZN(n682) );
  AOI21_X1 U616 ( .B1(B[26]), .B2(B[25]), .A(n682), .ZN(mode[13]) );
  INV_X1 U617 ( .A(B[25]), .ZN(n683) );
  AOI21_X1 U618 ( .B1(B[24]), .B2(B[23]), .A(n683), .ZN(mode[12]) );
  INV_X1 U619 ( .A(B[23]), .ZN(n684) );
  AOI21_X1 U620 ( .B1(B[22]), .B2(B[21]), .A(n684), .ZN(mode[11]) );
  INV_X1 U621 ( .A(B[21]), .ZN(n685) );
  AOI21_X1 U622 ( .B1(B[20]), .B2(B[19]), .A(n685), .ZN(mode[10]) );
  INV_X1 U623 ( .A(B[19]), .ZN(n686) );
  AOI21_X1 U624 ( .B1(B[18]), .B2(B[17]), .A(n686), .ZN(mode[9]) );
  INV_X1 U625 ( .A(B[17]), .ZN(n687) );
  AOI21_X1 U626 ( .B1(B[16]), .B2(B[15]), .A(n687), .ZN(mode[8]) );
  INV_X1 U627 ( .A(B[15]), .ZN(n688) );
  AOI21_X1 U628 ( .B1(B[14]), .B2(B[13]), .A(n688), .ZN(mode[7]) );
  INV_X1 U629 ( .A(B[13]), .ZN(n689) );
  AOI21_X1 U630 ( .B1(B[12]), .B2(B[11]), .A(n689), .ZN(mode[6]) );
  INV_X1 U631 ( .A(B[11]), .ZN(n690) );
  AOI21_X1 U632 ( .B1(B[10]), .B2(B[9]), .A(n690), .ZN(mode[5]) );
  INV_X1 U633 ( .A(B[9]), .ZN(n691) );
  AOI21_X1 U634 ( .B1(B[8]), .B2(B[7]), .A(n691), .ZN(mode[4]) );
  INV_X1 U635 ( .A(B[7]), .ZN(n692) );
  AOI21_X1 U636 ( .B1(B[6]), .B2(B[5]), .A(n692), .ZN(mode[3]) );
  INV_X1 U637 ( .A(B[5]), .ZN(n693) );
  AOI21_X1 U638 ( .B1(B[4]), .B2(B[3]), .A(n693), .ZN(mode[2]) );
  INV_X1 U639 ( .A(B[3]), .ZN(n694) );
  AOI21_X1 U640 ( .B1(B[2]), .B2(mode[0]), .A(n694), .ZN(mode[1]) );
  INV_X1 U641 ( .A(B[31]), .ZN(n695) );
  AOI21_X1 U642 ( .B1(B[30]), .B2(B[29]), .A(n695), .ZN(mode[15]) );
endmodule

