
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file_reg_size32_file_size64 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file_reg_size32_file_size64;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file_reg_size32_file_size64.all;

entity register_file_reg_size32_file_size64 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (5 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_reg_size32_file_size64;

architecture SYN_BEHAVIORAL of register_file_reg_size32_file_size64 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
      n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, 
      n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, 
      n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, 
      n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, 
      n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, 
      n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, 
      n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, 
      n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, 
      n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, 
      n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, 
      n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, 
      n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, 
      n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, 
      n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, 
      n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, 
      n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, 
      n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, 
      n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, 
      n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, 
      n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, 
      n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, 
      n4538, n4539, n4540, n4541, n4670, n4671, n4672, n4673, n4674, n4675, 
      n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, 
      n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, 
      n4696, n4697, n4698, n4699, n4700, n4701, n4798, n4799, n4800, n4801, 
      n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, 
      n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, 
      n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n5022, n5023, 
      n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, 
      n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, 
      n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, 
      n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, 
      n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, 
      n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, 
      n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, 
      n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, 
      n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, 
      n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, 
      n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, 
      n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, 
      n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, 
      n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, 
      n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, 
      n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, 
      n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, 
      n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, 
      n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, 
      n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, 
      n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, 
      n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, 
      n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, 
      n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, 
      n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, 
      n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, 
      n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, 
      n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, 
      n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, 
      n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, 
      n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, 
      n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, 
      n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, 
      n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, 
      n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, 
      n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, 
      n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, 
      n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, 
      n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, 
      n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, 
      n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, 
      n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, 
      n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, 
      n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, 
      n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, 
      n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, 
      n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, 
      n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, 
      n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, 
      n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, 
      n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, 
      n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, 
      n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, 
      n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, 
      n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, 
      n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, 
      n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, 
      n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, 
      n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, 
      n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, 
      n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, 
      n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, 
      n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, 
      n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, 
      n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, 
      n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, 
      n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, 
      n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, 
      n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, 
      n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, 
      n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, 
      n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, 
      n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, 
      n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, 
      n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, 
      n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, 
      n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, 
      n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, 
      n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, 
      n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, 
      n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, 
      n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, 
      n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, 
      n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, 
      n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, 
      n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, 
      n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, 
      n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, 
      n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, 
      n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, 
      n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, 
      n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, 
      n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, 
      n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, 
      n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, 
      n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, 
      n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, 
      n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, 
      n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, 
      n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, 
      n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, 
      n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, 
      n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, 
      n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, 
      n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, 
      n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, 
      n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, 
      n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, 
      n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, 
      n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, 
      n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, 
      n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, 
      n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, 
      n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, 
      n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, 
      n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, 
      n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, 
      n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, 
      n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, 
      n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, 
      n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, 
      n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, 
      n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, 
      n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, 
      n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, 
      n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, 
      n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, 
      n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, 
      n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, 
      n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, 
      n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, 
      n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, 
      n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, 
      n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, 
      n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, 
      n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, 
      n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, 
      n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, 
      n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, 
      n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, 
      n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, 
      n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, 
      n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, 
      n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, 
      n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, 
      n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, 
      n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, 
      n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, 
      n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, 
      n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, 
      n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, 
      n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, 
      n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, 
      n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, 
      n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, 
      n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, 
      n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, 
      n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, 
      n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, 
      n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, 
      n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, 
      n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, 
      n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, 
      n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, 
      n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, 
      n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, 
      n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, 
      n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, 
      n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, 
      n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, 
      n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, 
      n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, 
      n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, 
      n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, 
      n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, 
      n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, 
      n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, 
      n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, 
      n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, 
      n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, 
      n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, 
      n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, 
      n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, 
      n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, 
      n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, 
      n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, 
      n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, 
      n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, 
      n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, 
      n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, 
      n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, 
      n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, 
      n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, 
      n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, 
      n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, 
      n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, 
      n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, 
      n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, 
      n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, 
      n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, 
      n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, 
      n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, 
      n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, 
      n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, 
      n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, 
      n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, 
      n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, 
      n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, 
      n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, 
      n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, 
      n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, 
      n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, 
      n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, 
      n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, 
      n7452, n7453, n7454, n7456, n7457, n7466, n7467, n7474, n7475, n7478, 
      n7479, n7486, n7488, n7489, n7498, n7499, n7506, n7507, n7510, n7511, 
      n7518, n7520, n7521, n7530, n7531, n7538, n7539, n7542, n7543, n7550, 
      n7552, n7553, n7562, n7563, n7570, n7571, n7574, n7575, n7582, n7584, 
      n7585, n7594, n7595, n7602, n7603, n7606, n7607, n7614, n7616, n7617, 
      n7626, n7627, n7634, n7635, n7638, n7639, n7646, n7648, n7649, n7658, 
      n7659, n7666, n7667, n7670, n7671, n7678, n7680, n7681, n7690, n7691, 
      n7698, n7699, n7702, n7703, n7710, n7712, n7713, n7722, n7723, n7730, 
      n7731, n7734, n7735, n7742, n7744, n7745, n7754, n7755, n7762, n7763, 
      n7766, n7767, n7774, n7776, n7777, n7786, n7787, n7794, n7795, n7798, 
      n7799, n7806, n7808, n7809, n7818, n7819, n7826, n7827, n7830, n7831, 
      n7838, n7840, n7841, n7850, n7851, n7858, n7859, n7862, n7863, n7870, 
      n7872, n7873, n7882, n7883, n7890, n7891, n7894, n7895, n7904, n7905, 
      n7914, n7915, n7922, n7923, n7926, n7927, n7936, n7937, n7946, n7947, 
      n7954, n7955, n7958, n7959, n7968, n7969, n7978, n7979, n7986, n7987, 
      n7990, n7991, n8000, n8001, n8010, n8011, n8018, n8019, n8022, n8023, 
      n8032, n8033, n8042, n8043, n8050, n8051, n8054, n8055, n8064, n8065, 
      n8074, n8075, n8082, n8083, n8086, n8087, n8096, n8097, n8106, n8107, 
      n8114, n8115, n8118, n8119, n8128, n8129, n8138, n8139, n8146, n8147, 
      n8150, n8151, n8160, n8161, n8170, n8171, n8178, n8179, n8182, n8183, 
      n8192, n8193, n8202, n8203, n8210, n8211, n8214, n8215, n8224, n8225, 
      n8234, n8235, n8242, n8243, n8246, n8247, n8256, n8257, n8266, n8267, 
      n8274, n8275, n8278, n8279, n8288, n8289, n8298, n8299, n8306, n8307, 
      n8310, n8311, n8320, n8321, n8330, n8331, n8338, n8339, n8342, n8343, 
      n8352, n8353, n8362, n8363, n8370, n8371, n8374, n8375, n8384, n8385, 
      n8394, n8395, n8402, n8403, n8406, n8407, n8416, n8417, n8426, n8427, 
      n8434, n8435, n8438, n8439, n8448, n8449, n8458, n8459, n8466, n8467, 
      n8470, n8471, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, 
      n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, 
      n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, 
      n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, 
      n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, 
      n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, 
      n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, 
      n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, 
      n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, 
      n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, 
      n8576, n8578, n8580, n8582, n8584, n8585, n8586, n8587, n8589, n8591, 
      n8593, n8595, n8596, n8597, n8598, n8600, n8602, n8604, n8606, n8607, 
      n8608, n8609, n8611, n8613, n8615, n8617, n8618, n8619, n8620, n8622, 
      n8624, n8626, n8628, n8629, n8630, n8631, n8633, n8635, n8637, n8639, 
      n8640, n8641, n8642, n8644, n8646, n8648, n8650, n8651, n8652, n8653, 
      n8655, n8657, n8659, n8661, n8662, n8663, n8664, n8665, n8666, n8667, 
      n8668, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, 
      n8679, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, 
      n8690, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, 
      n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, 
      n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, 
      n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, 
      n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, 
      n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, 
      n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, 
      n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, 
      n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, 
      n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, 
      n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, 
      n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, 
      n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, 
      n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, 
      n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, 
      n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, 
      n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, 
      n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, 
      n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, 
      n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, 
      n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, 
      n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, 
      n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, 
      n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, 
      n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, 
      n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, 
      n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, 
      n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, 
      n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, 
      n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, 
      n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, 
      n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, 
      n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, 
      n9021, n9026, n9030, n9037, n9041, n9048, n9052, n9059, n9063, n9070, 
      n9074, n9081, n9085, n9092, n9096, n9103, n9107, n9112, n9114, n9115, 
      n9116, n9118, n9119, n9120, n9123, n9125, n9126, n9127, n9129, n9130, 
      n9131, n9134, n9136, n9137, n9138, n9140, n9141, n9142, n9145, n9147, 
      n9148, n9149, n9151, n9152, n9153, n9156, n9158, n9159, n9160, n9162, 
      n9163, n9164, n9167, n9169, n9170, n9171, n9173, n9174, n9175, n9178, 
      n9180, n9181, n9182, n9184, n9185, n9186, n9189, n9191, n9192, n9193, 
      n9195, n9196, n9197, n9200, n9202, n9203, n9204, n9206, n9207, n9208, 
      n9211, n9213, n9214, n9215, n9217, n9218, n9219, n9222, n9224, n9225, 
      n9226, n9228, n9229, n9230, n9233, n9235, n9236, n9237, n9239, n9240, 
      n9241, n9244, n9246, n9247, n9248, n9250, n9251, n9252, n9255, n9257, 
      n9258, n9259, n9261, n9262, n9263, n9266, n9268, n9269, n9270, n9272, 
      n9273, n9274, n9277, n9279, n9280, n9281, n9283, n9284, n9285, n9288, 
      n9290, n9291, n9292, n9294, n9295, n9296, n9299, n9301, n9302, n9303, 
      n9305, n9306, n9307, n9310, n9312, n9313, n9314, n9316, n9317, n9318, 
      n9321, n9323, n9324, n9325, n9327, n9328, n9329, n9332, n9334, n9335, 
      n9336, n9338, n9339, n9340, n9343, n9345, n9346, n9347, n9349, n9350, 
      n9351, n9354, n9356, n9357, n9358, n9360, n9361, n9362, n9365, n9367, 
      n9368, n9369, n9371, n9372, n9373, n9382, n9383, n9384, n9385, n9386, 
      n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, 
      n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9414, 
      n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, 
      n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, 
      n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, 
      n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, 
      n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, 
      n9465, n9466, n9467, n9468, n9469, n9478, n9479, n9480, n9481, n9482, 
      n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, 
      n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, 
      n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, 
      n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, 
      n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, 
      n9533, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, 
      n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, 
      n9561, n9562, n9563, n9564, n9565, n9574, n9575, n9576, n9577, n9578, 
      n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, 
      n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, 
      n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, 
      n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, 
      n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, 
      n9629, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, 
      n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, 
      n9657, n9658, n9659, n9660, n9661, n9734, n9735, n9736, n9737, n9738, 
      n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, 
      n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9766, 
      n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, 
      n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, 
      n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, 
      n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, 
      n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, 
      n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, 
      n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, 
      n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, 
      n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9886, n9887, n9888, 
      n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, 
      n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, 
      n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, 
      n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, 
      n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, 
      n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, 
      n9949, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, 
      n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, 
      n9977, n9978, n9979, n9980, n9981, n9990, n9991, n9992, n9993, n9994, 
      n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004
      , n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
      n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021, n10022, 
      n10023, n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031, 
      n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040, 
      n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048, n10049, 
      n10050, n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058, 
      n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067, 
      n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076, 
      n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085, 
      n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093, n10094, 
      n10095, n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103, 
      n10104, n10105, n10106, n10107, n10108, n10109, n10398, n10399, n10400, 
      n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408, n10409, 
      n10410, n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418, 
      n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427, 
      n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435, n10436, 
      n10437, n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445, 
      n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453, n10454, 
      n10455, n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463, 
      n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472, 
      n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480, n10481, 
      n10482, n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490, 
      n10491, n10492, n10493, n15118, n15119, n15120, n15121, n15122, n15123, 
      n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131, n15132, 
      n15133, n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141, 
      n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149, n15150, 
      n15151, n15152, n15153, n15155, n15156, n15158, n15159, n15160, n15161, 
      n15162, n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, 
      n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, 
      n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, 
      n15189, n15190, n15191, n15193, n15194, n15195, n15196, n15197, n15198, 
      n15199, n15200, n15201, n15226, n15227, n15228, n15230, n15231, n15232, 
      n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240, n15241, 
      n15242, n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250, 
      n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259, 
      n15260, n15261, n15262, n15263, n15265, n15266, n15267, n15268, n15269, 
      n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, 
      n15279, n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, 
      n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, 
      n15297, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, 
      n15307, n15331, n15333, n15334, n15335, n15336, n15337, n15338, n15339, 
      n15340, n15341, n15365, n15366, n15368, n15369, n15370, n15371, n15372, 
      n15373, n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381, 
      n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389, n15390, 
      n15391, n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399, 
      n15400, n15401, n15403, n15404, n15405, n15406, n15407, n15408, n15409, 
      n15410, n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418, 
      n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427, 
      n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435, n15437, 
      n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445, n15446, 
      n15447, n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455, 
      n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464, 
      n15465, n15466, n15467, n15468, n15469, n15471, n15472, n15473, n15474, 
      n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483, 
      n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491, n15492, 
      n15493, n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501, 
      n15502, n15503, n15504, n15506, n15507, n15508, n15509, n15510, n15511, 
      n15512, n15513, n15514, n15539, n15541, n15542, n15543, n15544, n15545, 
      n15546, n15547, n15548, n15549, n15575, n15576, n15577, n15578, n15579, 
      n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587, n15588, 
      n15589, n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597, 
      n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605, n15606, 
      n15607, n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616, 
      n15617, n15641, n15642, n15643, n15644, n15645, n15647, n15648, n15649, 
      n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658, 
      n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667, 
      n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, n15676, 
      n15677, n15678, n15679, n15680, n15682, n15683, n15684, n15685, n15686, 
      n15687, n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695, 
      n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704, 
      n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712, n15713, 
      n15714, n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723, 
      n15724, n15748, n15750, n15751, n15753, n15754, n15755, n15756, n15757, 
      n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, n15766, 
      n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775, 
      n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784, 
      n15785, n15786, n15788, n15789, n15790, n15791, n15792, n15793, n15794, 
      n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803, 
      n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811, n15812, 
      n15813, n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15822, 
      n15823, n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831, 
      n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840, 
      n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848, n15849, 
      n15850, n15851, n15852, n15853, n15854, n15856, n15857, n15858, n15859, 
      n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867, n15868, 
      n15869, n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877, 
      n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885, n15886, 
      n15887, n15888, n15890, n15891, n15893, n15895, n15896, n15897, n15898, 
      n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907, 
      n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915, n15916, 
      n15917, n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925, 
      n15926, n15927, n15929, n15930, n15931, n15932, n15933, n15934, n15935, 
      n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, 
      n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, 
      n15954, n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15963, 
      n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15996, 
      n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005, n16006, 
      n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040, 
      n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048, n16049, 
      n16050, n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058, 
      n16059, n16060, n16061, n16062, n16063, n16064, n16066, n16067, n16068, 
      n16069, n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077, 
      n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085, n16086, 
      n16087, n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095, 
      n16096, n16097, n16098, n16100, n16101, n16102, n16103, n16104, n16105, 
      n16106, n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114, 
      n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123, 
      n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131, n16132, 
      n16133, n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, 
      n16143, n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, 
      n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, 
      n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16169, n16171, 
      n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, n16180, 
      n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189, 
      n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, n16198, 
      n16199, n16200, n16201, n16202, n16203, n16204, n16206, n16207, n16208, 
      n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216, n16217, 
      n16218, n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226, 
      n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235, 
      n16236, n16237, n16238, n16239, n16241, n16242, n16243, n16244, n16245, 
      n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253, n16254, 
      n16255, n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263, 
      n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272, 
      n16273, n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282, 
      n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291, 
      n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299, n16300, 
      n16301, n16302, n16303, n16304, n16305, n16306, n16307, n16309, n16310, 
      n16311, n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319, 
      n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328, 
      n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336, n16337, 
      n16338, n16339, n16340, n16341, n16343, n16344, n16346, n16348, n16350, 
      n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, 
      n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, 
      n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, 
      n16378, n16379, n16380, n16381, n16382, n16384, n16385, n16386, n16387, 
      n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, n16396, 
      n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405, 
      n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, n16414, 
      n16415, n16416, n16417, n16419, n16420, n16421, n16422, n16423, n16424, 
      n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432, n16433, 
      n16434, n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442, 
      n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451, 
      n16453, n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461, 
      n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469, n16470, 
      n16471, n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479, 
      n16480, n16481, n16482, n16483, n16484, n16485, n16487, n16488, n16489, 
      n16490, n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498, 
      n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507, 
      n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515, n16516, 
      n16517, n16518, n16519, n16521, n16522, n16523, n16524, n16525, n16526, 
      n16527, n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535, 
      n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544, 
      n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552, n16553, 
      n16554, n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563, 
      n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571, n16572, 
      n16573, n16574, n16576, n16577, n16578, n16579, n16580, n16581, n16582, 
      n16583, n16584, n16608, n16610, n16611, n16613, n16614, n16616, n16618, 
      n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, 
      n16652, n16653, n16655, n16656, n16657, n16658, n16659, n16660, n16661, 
      n16662, n16663, n16688, n16690, n16691, n16692, n16693, n16694, n16695, 
      n16696, n16697, n16698, n16724, n16725, n16726, n16727, n16728, n16729, 
      n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738, 
      n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747, 
      n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, n16756, 
      n16758, n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767, 
      n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776, 
      n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784, n16785, 
      n16786, n16787, n16788, n16789, n16790, n16791, n16793, n16794, n16795, 
      n16797, n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805, 
      n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813, n16814, 
      n16815, n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823, 
      n16824, n16825, n16826, n16827, n16828, n16831, n16832, n16834, n16835, 
      n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, 
      n16845, n16846, n16847, n16848, n16849, n16851, n16852, n16853, n16854, 
      n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, 
      n16864, n16865, n16866, n16867, n16868, n16869, n16871, n16872, n16873, 
      n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882, 
      n16883, n16884, n16885, n16887, n16888, n16889, n16890, n16892, n16893, 
      n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901, n16903, 
      n16904, n16905, n16906, n16907, n16908, n16910, n16912, n16913, n16915, 
      n16916, n16918, n16919, n16920, n16921, n16922, n16924, n16925, n16926, 
      n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, 
      n16936, n16937, n16938, n16939, n16941, n16942, n16943, n16944, n16945, 
      n16946, n16947, n16949, n16950, n16951, n16952, n16953, n16954, n16955, 
      n16956, n16958, n16960, n16961, n16963, n16964, n16965, n16966, n16967, 
      n16969, n16971, n16972, n16975, n16977, n16978, n16979, n16980, n16981, 
      n16982, n16983, n16984, n16985, n16986, n16988, n16989, n16990, n16991, 
      n16992, n16993, n16994, n16996, n16997, n16998, n16999, n17000, n17001, 
      n17002, n17003, n17005, n17007, n17008, n17010, n17011, n17012, n17013, 
      n17014, n17016, n17018, n17019, n17022, n17024, n17025, n17026, n17027, 
      n17028, n17029, n17030, n17031, n17032, n17033, n17035, n17036, n17037, 
      n17038, n17039, n17040, n17041, n17043, n17044, n17045, n17046, n17047, 
      n17048, n17049, n17050, n17052, n17054, n17055, n17057, n17058, n17059, 
      n17060, n17061, n17063, n17065, n17066, n17069, n17071, n17072, n17073, 
      n17074, n17075, n17076, n17077, n17078, n17079, n17080, n17082, n17083, 
      n17084, n17085, n17086, n17087, n17088, n17090, n17091, n17092, n17093, 
      n17094, n17095, n17096, n17097, n17099, n17101, n17102, n17104, n17105, 
      n17106, n17107, n17108, n17110, n17112, n17113, n17116, n17118, n17119, 
      n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17129, 
      n17130, n17131, n17132, n17133, n17134, n17135, n17137, n17138, n17139, 
      n17140, n17141, n17142, n17143, n17144, n17146, n17148, n17149, n17151, 
      n17152, n17153, n17154, n17155, n17157, n17159, n17160, n17163, n17165, 
      n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173, n17174, 
      n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17184, n17185, 
      n17186, n17187, n17188, n17189, n17190, n17191, n17193, n17195, n17196, 
      n17198, n17199, n17200, n17201, n17202, n17204, n17206, n17207, n17210, 
      n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219, n17220, 
      n17221, n17223, n17224, n17225, n17226, n17227, n17228, n17229, n17231, 
      n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17240, n17242, 
      n17243, n17245, n17246, n17247, n17248, n17249, n17251, n17253, n17254, 
      n17257, n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266, 
      n17267, n17268, n17270, n17271, n17272, n17273, n17274, n17275, n17276, 
      n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17287, 
      n17289, n17290, n17292, n17293, n17294, n17295, n17296, n17298, n17300, 
      n17301, n17304, n17306, n17307, n17308, n17309, n17310, n17311, n17312, 
      n17313, n17314, n17315, n17317, n17318, n17319, n17320, n17321, n17322, 
      n17323, n17325, n17326, n17327, n17328, n17329, n17330, n17331, n17332, 
      n17334, n17336, n17337, n17339, n17340, n17341, n17342, n17343, n17345, 
      n17347, n17348, n17351, n17353, n17354, n17355, n17356, n17357, n17358, 
      n17359, n17360, n17361, n17362, n17364, n17365, n17366, n17367, n17368, 
      n17369, n17370, n17372, n17373, n17374, n17375, n17376, n17377, n17378, 
      n17379, n17381, n17383, n17384, n17386, n17387, n17388, n17389, n17390, 
      n17392, n17394, n17395, n17398, n17400, n17401, n17402, n17403, n17404, 
      n17405, n17406, n17407, n17408, n17409, n17411, n17412, n17413, n17414, 
      n17415, n17416, n17417, n17419, n17420, n17421, n17422, n17423, n17424, 
      n17425, n17426, n17428, n17430, n17431, n17433, n17434, n17435, n17436, 
      n17437, n17439, n17441, n17442, n17445, n17447, n17448, n17449, n17450, 
      n17451, n17452, n17453, n17454, n17455, n17456, n17458, n17459, n17460, 
      n17461, n17462, n17463, n17464, n17466, n17467, n17468, n17469, n17470, 
      n17471, n17472, n17473, n17475, n17477, n17478, n17480, n17481, n17482, 
      n17483, n17484, n17486, n17488, n17489, n17492, n17494, n17495, n17496, 
      n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17505, n17506, 
      n17507, n17508, n17509, n17510, n17511, n17513, n17514, n17515, n17516, 
      n17517, n17518, n17519, n17520, n17522, n17524, n17525, n17527, n17528, 
      n17529, n17530, n17531, n17533, n17535, n17536, n17539, n17541, n17542, 
      n17543, n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17552, 
      n17553, n17554, n17555, n17556, n17557, n17558, n17560, n17561, n17562, 
      n17563, n17564, n17565, n17566, n17567, n17569, n17571, n17572, n17574, 
      n17575, n17576, n17577, n17578, n17580, n17582, n17583, n17586, n17588, 
      n17589, n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597, 
      n17599, n17600, n17601, n17602, n17603, n17604, n17605, n17607, n17608, 
      n17609, n17610, n17611, n17612, n17613, n17614, n17616, n17618, n17619, 
      n17621, n17622, n17623, n17624, n17625, n17627, n17629, n17630, n17633, 
      n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643, 
      n17644, n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17654, 
      n17655, n17656, n17657, n17658, n17659, n17660, n17661, n17663, n17665, 
      n17666, n17668, n17669, n17670, n17671, n17672, n17674, n17676, n17677, 
      n17680, n17682, n17683, n17684, n17685, n17686, n17687, n17688, n17689, 
      n17690, n17691, n17693, n17694, n17695, n17696, n17697, n17698, n17699, 
      n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17710, 
      n17712, n17713, n17715, n17716, n17717, n17718, n17719, n17721, n17723, 
      n17724, n17727, n17729, n17730, n17731, n17732, n17733, n17734, n17735, 
      n17736, n17737, n17738, n17740, n17741, n17742, n17743, n17744, n17745, 
      n17746, n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755, 
      n17757, n17759, n17760, n17762, n17763, n17764, n17765, n17766, n17768, 
      n17770, n17771, n17774, n17776, n17777, n17778, n17779, n17780, n17781, 
      n17782, n17783, n17784, n17785, n17787, n17788, n17789, n17790, n17791, 
      n17792, n17793, n17795, n17796, n17797, n17798, n17799, n17800, n17801, 
      n17802, n17804, n17806, n17807, n17809, n17810, n17811, n17812, n17813, 
      n17815, n17817, n17818, n17821, n17823, n17824, n17825, n17826, n17827, 
      n17828, n17829, n17830, n17831, n17832, n17834, n17835, n17836, n17837, 
      n17838, n17839, n17840, n17842, n17843, n17844, n17845, n17846, n17847, 
      n17848, n17849, n17851, n17853, n17854, n17856, n17857, n17858, n17859, 
      n17860, n17862, n17864, n17865, n17868, n17870, n17871, n17872, n17873, 
      n17874, n17875, n17876, n17877, n17878, n17879, n17881, n17882, n17883, 
      n17884, n17885, n17886, n17887, n17889, n17890, n17891, n17892, n17893, 
      n17894, n17895, n17896, n17898, n17900, n17901, n17903, n17904, n17905, 
      n17906, n17907, n17909, n17911, n17912, n17915, n17917, n17918, n17919, 
      n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17928, n17929, 
      n17930, n17931, n17932, n17933, n17934, n17936, n17937, n17938, n17939, 
      n17940, n17941, n17942, n17943, n17945, n17947, n17948, n17950, n17951, 
      n17952, n17953, n17954, n17956, n17958, n17959, n17962, n17964, n17965, 
      n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973, n17975, 
      n17976, n17977, n17978, n17979, n17980, n17981, n17983, n17984, n17985, 
      n17986, n17987, n17988, n17989, n17990, n17992, n17994, n17995, n17997, 
      n17998, n17999, n18000, n18001, n18003, n18005, n18006, n18009, n18011, 
      n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019, n18020, 
      n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18030, n18031, 
      n18032, n18033, n18034, n18035, n18036, n18037, n18039, n18041, n18042, 
      n18044, n18045, n18046, n18047, n18048, n18050, n18052, n18053, n18056, 
      n18058, n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066, 
      n18067, n18069, n18070, n18071, n18072, n18073, n18074, n18075, n18077, 
      n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18086, n18088, 
      n18089, n18091, n18092, n18093, n18094, n18095, n18097, n18099, n18100, 
      n18103, n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112, 
      n18113, n18114, n18116, n18117, n18118, n18119, n18120, n18121, n18122, 
      n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18133, 
      n18135, n18136, n18138, n18139, n18140, n18141, n18142, n18144, n18146, 
      n18147, n18150, n18152, n18153, n18154, n18155, n18156, n18157, n18158, 
      n18159, n18160, n18161, n18163, n18164, n18165, n18166, n18167, n18168, 
      n18169, n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178, 
      n18180, n18182, n18183, n18185, n18186, n18187, n18188, n18189, n18191, 
      n18193, n18194, n18197, n18199, n18200, n18201, n18202, n18203, n18204, 
      n18205, n18206, n18207, n18208, n18210, n18211, n18212, n18213, n18214, 
      n18215, n18216, n18218, n18219, n18220, n18221, n18222, n18223, n18224, 
      n18225, n18227, n18229, n18230, n18232, n18233, n18234, n18235, n18236, 
      n18238, n18240, n18241, n18244, n18246, n18247, n18248, n18249, n18250, 
      n18251, n18252, n18253, n18254, n18255, n18257, n18258, n18259, n18260, 
      n18261, n18262, n18263, n18265, n18266, n18267, n18268, n18269, n18270, 
      n18271, n18272, n18274, n18276, n18277, n18279, n18280, n18281, n18282, 
      n18283, n18285, n18287, n18288, n18291, n18293, n18294, n18295, n18296, 
      n18297, n18298, n18299, n18300, n18301, n18302, n18304, n18305, n18306, 
      n18307, n18308, n18309, n18310, n18312, n18313, n18314, n18315, n18316, 
      n18317, n18318, n18319, n18321, n18323, n18324, n18326, n18327, n18328, 
      n18329, n18330, n18332, n18334, n18335, n18338, n18340, n18341, n18342, 
      n18343, n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351, 
      n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360, 
      n18361, n18362, n18363, n18365, n18366, n18367, n18368, n18369, n18371, 
      n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379, n18380, 
      n18382, n18384, n18385, n18387, n18388, n18389, n18390, n18391, n18393, 
      n18394, n18395, n18396, n18397, n18399, n18400, n18401, n18402, n18403, 
      n18405, n18406, n18408, n18409, n18410, n18411, n18413, n18414, n18415, 
      n18416, n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424, 
      n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432, n18433, 
      n18434, n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442, 
      n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451, 
      n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459, n18460, 
      n18461, n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469, 
      n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477, n18478, 
      n18479, n18480, n18481, n18482, n18483, n18484, n18485, n18486, n18487, 
      n18488, n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496, 
      n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504, n18505, 
      n18506, n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514, 
      n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523, 
      n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531, n18532, 
      n18533, n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541, 
      n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549, n18550, 
      n18551, n18552, n18553, n18554, n18555, n18556, n18557, n18558, n18559, 
      n18560, n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568, 
      n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576, n18577, 
      n18578, n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586, 
      n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595, 
      n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603, n18604, 
      n18605, n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613, 
      n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621, n18622, 
      n18623, n18624, n18625, n18626, n18627, n18628, n18629, n18630, n18631, 
      n18632, n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640, 
      n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648, n18649, 
      n18650, n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658, 
      n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667, 
      n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675, n18676, 
      n18677, n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685, 
      n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693, n18694, 
      n18695, n18696, n18697, n18698, n18699, n18700, n18701, n18702, n18703, 
      n18704, n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712, 
      n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720, n18721, 
      n18722, n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730, 
      n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739, 
      n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747, n18748, 
      n18749, n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757, 
      n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765, n18766, 
      n18767, n18768, n18769, n18770, n18771, n18772, n18773, n18774, n18775, 
      n18776, n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784, 
      n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792, n18793, 
      n18794, n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802, 
      n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811, 
      n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819, n18820, 
      n18821, n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829, 
      n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837, n18838, 
      n18839, n18840, n18841, n18842, n18843, n18844, n18845, n18846, n18847, 
      n18848, n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856, 
      n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864, n18865, 
      n18866, n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874, 
      n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883, 
      n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891, n18892, 
      n18893, n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901, 
      n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909, n18910, 
      n18911, n18912, n18913, n18914, n18915, n18916, n18917, n18918, n18919, 
      n18920, n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928, 
      n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936, n18937, 
      n18938, n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946, 
      n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955, 
      n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963, n18964, 
      n18965, n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973, 
      n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981, n18982, 
      n18983, n18984, n18985, n18986, n18987, n18988, n18989, n18990, n18991, 
      n18992, n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000, 
      n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008, n19009, 
      n19010, n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018, 
      n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027, 
      n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035, n19036, 
      n19037, n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045, 
      n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053, n19054, 
      n19055, n19056, n19057, n19058, n19059, n19060, n19061, n19062, n19063, 
      n19064, n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072, 
      n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080, n19081, 
      n19082, n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090, 
      n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099, 
      n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107, n19108, 
      n19109, n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117, 
      n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125, n19126, 
      n19127, n19128, n19129, n19130, n19131, n19132, n19133, n19134, n19135, 
      n19136, n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144, 
      n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152, n19153, 
      n19154, n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162, 
      n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171, 
      n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179, n19180, 
      n19181, n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189, 
      n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197, n19198, 
      n19199, n19200, n19201, n19202, n19203, n19204, n19205, n19206, n19207, 
      n19208, n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216, 
      n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224, n19225, 
      n19226, n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234, 
      n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243, 
      n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251, n19252, 
      n19253, n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261, 
      n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269, n19270, 
      n19271, n19272, n19273, n19274, n19275, n19276, n19277, n19278, n19279, 
      n19280, n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288, 
      n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296, n19297, 
      n19298, n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306, 
      n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315, 
      n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323, n19324, 
      n19325, n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333, 
      n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341, n19342, 
      n19343, n19344, n19345, n19346, n19347, n19348, n19349, n19350, n19351, 
      n19352, n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360, 
      n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368, n19369, 
      n19370, n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378, 
      n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387, 
      n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395, n19396, 
      n19397, n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405, 
      n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413, n19414, 
      n19415, n19416, n19417, n19418, n19419, n19420, n19421, n19422, n19423, 
      n19424, n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432, 
      n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440, n19441, 
      n19442, n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450, 
      n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459, 
      n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467, n19468, 
      n19469, n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477, 
      n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485, n19486, 
      n19487, n19488, n19489, n19490, n19491, n19492, n19493, n19494, n19495, 
      n19496, n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504, 
      n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512, n19513, 
      n19514, n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522, 
      n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531, 
      n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539, n19540, 
      n19541, n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549, 
      n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557, n19558, 
      n19559, n19560, n19561, n19562, n19563, n19564, n19565, n19566, n19567, 
      n19568, n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576, 
      n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584, n19585, 
      n19586, n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594, 
      n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603, 
      n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611, n19612, 
      n19613, n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621, 
      n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629, n19630, 
      n19631, n19632, n19633, n19634, n19635, n19636, n19637, n19638, n19639, 
      n19640, n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648, 
      n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656, n19657, 
      n19658, n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666, 
      n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675, 
      n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683, n19684, 
      n19685, n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693, 
      n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701, n19702, 
      n19703, n19704, n19705, n19706, n19707, n19708, n19709, n19710, n19711, 
      n19712, n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720, 
      n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728, n19729, 
      n19730, n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738, 
      n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747, 
      n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755, n19756, 
      n19757, n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765, 
      n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773, n19774, 
      n19775, n19776, n19777, n19778, n19779, n19780, n19781, n19782, n19783, 
      n19784, n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792, 
      n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800, n19801, 
      n19802, n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810, 
      n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819, 
      n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827, n19828, 
      n19829, n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837, 
      n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845, n19846, 
      n19847, n19848, n19849, n19850, n19851, n19852, n19853, n19854, n19855, 
      n19856, n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864, 
      n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872, n19873, 
      n19874, n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882, 
      n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891, 
      n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899, n19900, 
      n19901, n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909, 
      n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917, n19918, 
      n19919, n19920, n19921, n19922, n19923, n19924, n19925, n19926, n19927, 
      n19928, n19929, n19930, n19931, n19932, n19933, n19934, n19935, n19936, 
      n19937, n19938, n19939, n19940, n19941, n19942, n19943, n19944, n19945, 
      n19946, n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954, 
      n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963, 
      n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971, n19972, 
      n19973, n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981, 
      n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989, n19990, 
      n19991, n19992, n19993, n19994, n19995, n19996, n19997, n19998, n19999, 
      n20000, n20001, n20002, n20003, n20004, n20005, n20006, n20007, n20008, 
      n20009, n20010, n20011, n20012, n20013, n20014, n20015, n20016, n20017, 
      n20018, n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026, 
      n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035, 
      n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043, n20044, 
      n20045, n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053, 
      n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061, n20062, 
      n20063, n20064, n20065, n20066, n20067, n20068, n20069, n20070, n20071, 
      n20072, n20073, n20074, n20075, n20076, n20077, n20078, n20079, n20080, 
      n20081, n20082, n20083, n20084, n20085, n20086, n20087, n20088, n20089, 
      n20090, n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098, 
      n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107, 
      n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115, n20116, 
      n20117, n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125, 
      n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133, n20134, 
      n20135, n20136, n20137, n20138, n20139, n20140, n20141, n20142, n20143, 
      n20144, n20145, n20146, n20147, n20148, n20149, n20150, n20151, n20152, 
      n20153, n20154, n20155, n20156, n20157, n20158, n20159, n20160, n20161, 
      n20162, n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170, 
      n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179, 
      n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187, n20188, 
      n20189, n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197, 
      n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205, n20206, 
      n20207, n20208, n20209, n20210, n20211, n20212, n20213, n20214, n20215, 
      n20216, n20217, n20218, n20219, n20220, n20221, n20222, n20223, n20224, 
      n20225, n20226, n20227, n20228, n20229, n20230, n20231, n20232, n20233, 
      n20234, n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242, 
      n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251, 
      n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259, n20260, 
      n20261, n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269, 
      n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277, n20278, 
      n20279, n20280, n20281, n20282, n20283, n20284, n20285, n20286, n20287, 
      n20288, n20289, n20290, n20291, n20292, n20293, n20294, n20295, n20296, 
      n20297, n20298, n20299, n20300, n20301, n20302, n20303, n20304, n20305, 
      n20306, n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314, 
      n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323, 
      n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331, n20332, 
      n20333, n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341, 
      n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349, n20350, 
      n20351, n20352, n20353, n20354, n20355, n20356, n20357, n20358, n20359, 
      n20360, n20361, n20362, n20363, n20364, n20365, n20366, n20367, n20368, 
      n20369, n20370, n20371, n20372, n20373, n20374, n20375, n20376, n20377, 
      n20378, n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386, 
      n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395, 
      n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403, n20404, 
      n20405, n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413, 
      n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421, n20422, 
      n20423, n20424, n20425, n20426, n20427, n20428, n20429, n20430, n20431, 
      n20432, n20433, n20434, n20435, n20436, n20437, n20438, n20439, n20440, 
      n20441, n20442, n20443, n20444, n20445, n20446, n20447, n20448, n20449, 
      n20450, n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458, 
      n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467, 
      n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475, n20476, 
      n20477, n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485, 
      n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493, n20494, 
      n20495, n20496, n20497, n20498, n20499, n20500, n20501, n20502, n20503, 
      n20504, n20505, n20506, n20507, n20508, n20509, n20510, n20511, n20512, 
      n20513, n20514, n20515, n20516, n20517, n20518, n20519, n20520, n20521, 
      n20522, n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530, 
      n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539, 
      n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547, n20548, 
      n20549, n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557, 
      n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565, n20566, 
      n20567, n20568, n20569, n20570, n20571, n20572, n20573, n20574, n20575, 
      n20576, n20577, n20578, n20579, n20580, n20581, n20582, n20583, n20584, 
      n20585, n20586, n20587, n20588, n20589, n20590, n20591, n20592, n20593, 
      n20594, n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602, 
      n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611, 
      n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619, n20620, 
      n20621, n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629, 
      n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637, n20638, 
      n20639, n20640, n20641, n20642, n20643, n20644, n20645, n20646, n20647, 
      n20648, n20649, n20650, n20651, n20652, n20653, n20654, n20655, n20656, 
      n20657, n20658, n20659, n20660, n20661, n20662, n20663, n20664, n20665, 
      n20666, n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674, 
      n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683, 
      n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691, n20692, 
      n20693, n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701, 
      n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709, n20710, 
      n20711, n20712, n20713, n20714, n20715, n20716, n20717, n20718, n20719, 
      n20720, n20721, n20722, n20723, n20724, n20725, n20726, n20727, n20728, 
      n20729, n20730, n20731, n20732, n20733, n20734, n20735, n20736, n20737, 
      n20738, n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746, 
      n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755, 
      n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763, n20764, 
      n20765, n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773, 
      n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781, n20782, 
      n20783, n20784, n20785, n20786, n20787, n20788, n20789, n20790, n20791, 
      n20792, n20793, n20794, n20795, n20796, n20797, n20798, n20799, n20800, 
      n20801, n20802, n20803, n20804, n20805, n20806, n20807, n20808, n20809, 
      n20810, n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818, 
      n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827, 
      n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835, n20836, 
      n20837, n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845, 
      n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853, n20854, 
      n20855, n20856, n20857, n20858, n20859, n20860, n20861, n20862, n20863, 
      n20864, n20865, n20866, n20867, n20868, n20869, n20870, n20871, n20872, 
      n20873, n20874, n20875, n20876, n20877, n20878, n20879, n20880, n20881, 
      n20882, n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890, 
      n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899, 
      n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907, n20908, 
      n20909, n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917, 
      n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925, n20926, 
      n20927, n20928, n20929, n20930, n20931, n20932, n20933, n20934, n20935, 
      n20936, n20937, n20938, n20939, n20940, n20941, n20942, n20943, n20944, 
      n20945, n20946, n20947, n20948, n20949, n20950, n20951, n20952, n20953, 
      n20954, n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962, 
      n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971, 
      n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979, n20980, 
      n20981, n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989, 
      n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997, n20998, 
      n20999, n21000, n21001, n21002, n21003, n21004, n21005, n21006, n21007, 
      n21008, n21009, n21010, n21011, n21012, n21013, n21014, n21015, n21016, 
      n21017, n21018, n21019, n21020, n21021, n21022, n21023, n21024, n21025, 
      n21026, n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034, 
      n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043, 
      n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051, n21052, 
      n21053, n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061, 
      n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069, n21070, 
      n21071, n21072, n21073, n21074, n21075, n21076, n21077, n21078, n21079, 
      n21080, n21081, n21082, n21083, n21084, n21085, n21086, n21087, n21088, 
      n21089, n21090, n21091, n21092, n21093, n21094, n21095, n21096, n21097, 
      n21098, n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106, 
      n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115, 
      n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123, n21124, 
      n21125, n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133, 
      n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141, n21142, 
      n21143, n21144, n21145, n21146, n21147, n21148, n21149, n21150, n21151, 
      n21152, n21153, n21154, n21155, n21156, n21157, n21158, n21159, n21160, 
      n21161, n21162, n21163, n21164, n21165, n21166, n21167, n21168, n21169, 
      n21170, n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178, 
      n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187, 
      n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195, n21196, 
      n21197, n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205, 
      n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213, n21214, 
      n21215, n21216, n21217, n21218, n21219, n21220, n21221, n21222, n21223, 
      n21224, n21225, n21226, n21227, n21228, n21229, n21230, n21231, n21232, 
      n21233, n21234, n21235, n21236, n21237, n21238, n21239, n21240, n21241, 
      n21242, n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250, 
      n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259, 
      n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267, n21268, 
      n21269, n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277, 
      n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285, n21286, 
      n21287, n21288, n21289, n21290, n21291, n21292, n21293, n21294, n21295, 
      n21296, n21297, n21298, n21299, n21300, n21301, n21302, n21303, n21304, 
      n21305, n21306, n21307, n21308, n21309, n21310, n21311, n21312, n21313, 
      n21314, n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322, 
      n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331, 
      n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339, n21340, 
      n21341, n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349, 
      n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357, n21358, 
      n21359, n21360, n21361, n21362, n21363, n21364, n21365, n21366, n21367, 
      n21368, n21369, n21370, n21371, n21372, n21373, n21374, n21375, n21376, 
      n21377, n21378, n21379, n21380, n21381, n21382, n21383, n21384, n21385, 
      n21386, n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394, 
      n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403, 
      n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411, n21412, 
      n21413, n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421, 
      n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429, n21430, 
      n21431, n21432, n21433, n21434, n21435, n21436, n21437, n21438, n21439, 
      n21440, n21441, n21442, n21443, n21444, n21445, n21446, n21447, n21448, 
      n21449, n21450, n21451, n21452, n21453, n21454, n21455, n21456, n21457, 
      n21458, n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466, 
      n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475, 
      n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483, n21484, 
      n21485, n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493, 
      n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501, n21502, 
      n21503, n21504, n21505, n21506, n21507, n21508, n21509, n21510, n21511, 
      n21512, n21513, n21514, n21515, n21516, n21517, n21518, n21519, n21520, 
      n21521, n21522, n21523, n21524, n21525, n21526, n21527, n21528, n21529, 
      n21530, n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538, 
      n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547, 
      n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555, n21556, 
      n21557, n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565, 
      n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573, n21574, 
      n21575, n21576, n21577, n21578, n21579, n21580, n21581, n21582, n21583, 
      n21584, n21585, n21586, n21587, n21588, n21589, n21590, n21591, n21592, 
      n21593, n21594, n21595, n21596, n21597, n21598, n21599, n21600, n21601, 
      n21602, n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610, 
      n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619, 
      n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627, n21628, 
      n21629, n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637, 
      n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645, n21646, 
      n21647, n21648, n21649, n21650, n21651, n21652, n21653, n21654, n21655, 
      n21656, n21657, n21658, n21659, n21660, n21661, n21662, n21663, n21664, 
      n21665, n21666, n21667, n21668, n21669, n21670, n21671, n21672, n21673, 
      n21674, n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682, 
      n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691, 
      n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699, n21700, 
      n21701, n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709, 
      n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717, n21718, 
      n21719, n21720, n21721, n21722, n21723, n21724, n21725, n21726, n21727, 
      n21728, n21729, n21730, n21731, n21732, n21733, n21734, n21735, n21736, 
      n21737, n21738, n21739, n21740, n21741, n21742, n21743, n21744, n21745, 
      n21746, n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754, 
      n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763, 
      n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771, n21772, 
      n21773, n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781, 
      n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789, n21790, 
      n21791, n21792, n21793, n21794, n21795, n21796, n21797, n21798, n21799, 
      n21800, n21801, n21802, n21803, n21804, n21805, n21806, n21807, n21808, 
      n21809, n21810, n21811, n21812, n21813, n21814, n21815, n21816, n21817, 
      n21818, n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826, 
      n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835, 
      n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843, n21844, 
      n21845, n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853, 
      n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861, n21862, 
      n21863, n21864, n21865, n21866, n21867, n21868, n21869, n21870, n21871, 
      n21872, n21873, n21874, n21875, n21876, n21877, n21878, n21879, n21880, 
      n21881, n21882, n21883, n21884, n21885, n21886, n21887, n21888, n21889, 
      n21890, n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898, 
      n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907, 
      n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915, n21916, 
      n21917, n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925, 
      n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933, n21934, 
      n21935, n21936, n21937, n21938, n21939, n21940, n21941, n21942, n21943, 
      n21944, n21945, n21946, n21947, n21948, n21949, n21950, n21951, n21952, 
      n21953, n21954, n21955, n21956, n21957, n21958, n21959, n21960, n21961, 
      n21962, n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970, 
      n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979, 
      n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987, n21988, 
      n21989, n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997, 
      n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005, n22006, 
      n22007, n22008, n22009, n22010, n22011, n22012, n22013, n22014, n22015, 
      n22016, n22017, n22018, n22019, n22020, n22021, n22022, n22023, n22024, 
      n22025, n22026, n22027, n22028, n22029, n22030, n22031, n22032, n22033, 
      n22034, n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042, 
      n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051, 
      n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059, n22060, 
      n22061, n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069, 
      n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077, n22078, 
      n22079, n22080, n22081, n22082, n22083, n22084, n22085, n22086, n22087, 
      n22088, n22089, n22090, n22091, n22092, n22093, n22094, n22095, n22096, 
      n22097, n22098, n22099, n22100, n22101, n22102, n22103, n22104, n22105, 
      n22106, n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114, 
      n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123, 
      n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131, n22132, 
      n22133, n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141, 
      n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149, n22150, 
      n22151, n22152, n22153, n22154, n22155, n22156, n22157, n22158, n22159, 
      n22160, n22161, n22162, n22163, n22164, n22165, n22166, n22167, n22168, 
      n22169, n22170, n22171, n22172, n22173, n22174, n22175, n22176, n22177, 
      n22178, n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186, 
      n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195, 
      n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203, n22204, 
      n22205, n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213, 
      n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221, n22222, 
      n22223, n22224, n22225, n22226, n22227, n22228, n22229, n22230, n22231, 
      n22232, n22233, n22234, n22235, n22236, n22237, n22238, n22239, n22240, 
      n22241, n22242, n22243, n22244, n22245, n22246, n22247, n22248, n22249, 
      n22250, n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258, 
      n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267, 
      n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275, n22276, 
      n22277, n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285, 
      n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293, n22294, 
      n22295, n22296, n22297, n22298, n22299, n22300, n22301, n22302, n22303, 
      n22304, n22305, n22306, n22307, n22308, n22309, n22310, n22311, n22312, 
      n22313, n22314, n22315, n22316, n22317, n22318, n22319, n22320, n22321, 
      n22322, n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330, 
      n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339, 
      n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347, n22348, 
      n22349, n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357, 
      n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365, n22366, 
      n22367, n22368, n22369, n22370, n22371, n22372, n22373, n22374, n22375, 
      n22376, n22377, n22378, n22379, n22380, n22381, n22382, n22383, n22384, 
      n22385, n22386, n22387, n22388, n22389, n22390, n22391, n22392, n22393, 
      n22394, n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402, 
      n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411, 
      n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419, n22420, 
      n22421, n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429, 
      n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437, n22438, 
      n22439, n22440, n22441, n22442, n22443, n22444, n22445, n22446, n22447, 
      n22448, n22449, n22450, n22451, n22452, n22453, n22454, n22455, n22456, 
      n22457, n22458, n22459, n22460, n22461, n22462, n22463, n22464, n22465, 
      n22466, n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474, 
      n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483, 
      n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491, n22492, 
      n22493, n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501, 
      n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509, n22510, 
      n22511, n22512, n22513, n22514, n22515, n22516, n22517, n22518, n22519, 
      n22520, n22521, n22522, n22523, n22524, n22525, n22526, n22527, n22528, 
      n22529, n22530, n22531, n22532, n22533, n22534, n22535, n22536, n22537, 
      n22538, n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546, 
      n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555, 
      n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563, n22564, 
      n22565, n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573, 
      n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581 : 
      std_logic;

begin
   
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n7453, CK => CLK, Q => 
                           n19996, QN => n8471);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n7452, CK => CLK, Q => 
                           n19994, QN => n8439);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n7451, CK => CLK, Q => 
                           n19992, QN => n8407);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n7450, CK => CLK, Q => 
                           n19990, QN => n8375);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n7449, CK => CLK, Q => 
                           n19988, QN => n8343);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n7448, CK => CLK, Q => 
                           n19986, QN => n8311);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n7447, CK => CLK, Q => 
                           n19984, QN => n8279);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n7446, CK => CLK, Q => 
                           n19982, QN => n8247);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n7445, CK => CLK, Q => 
                           n19980, QN => n8215);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n7444, CK => CLK, Q => 
                           n19978, QN => n8183);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n7443, CK => CLK, Q => 
                           n19691, QN => n8151);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n7442, CK => CLK, Q => 
                           n19975, QN => n8119);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n7441, CK => CLK, Q => 
                           n19690, QN => n8087);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n7440, CK => CLK, Q => 
                           n19998, QN => n8055);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n7439, CK => CLK, Q => 
                           n19971, QN => n8023);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n7438, CK => CLK, Q => 
                           n19969, QN => n7991);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n7437, CK => CLK, Q => 
                           n19967, QN => n7959);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n7436, CK => CLK, Q => 
                           n19965, QN => n7927);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n7435, CK => CLK, Q => 
                           n19963, QN => n7895);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n7434, CK => CLK, Q => 
                           n19961, QN => n7863);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n7433, CK => CLK, Q => 
                           n19959, QN => n7831);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n7432, CK => CLK, Q => 
                           n19957, QN => n7799);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n7431, CK => CLK, Q => n19955
                           , QN => n7767);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n7430, CK => CLK, Q => n19953
                           , QN => n7735);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n7429, CK => CLK, Q => n19951
                           , QN => n7703);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n7428, CK => CLK, Q => n19949
                           , QN => n7671);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n7427, CK => CLK, Q => n19947
                           , QN => n7639);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n7426, CK => CLK, Q => n19945
                           , QN => n7607);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n7425, CK => CLK, Q => n19943
                           , QN => n7575);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n7424, CK => CLK, Q => n19941
                           , QN => n7543);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n7423, CK => CLK, Q => n19939
                           , QN => n7511);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n7422, CK => CLK, Q => n19937
                           , QN => n7479);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n7421, CK => CLK, Q => 
                           n19997, QN => n8470);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n7420, CK => CLK, Q => 
                           n19995, QN => n8438);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n7419, CK => CLK, Q => 
                           n19993, QN => n8406);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n7418, CK => CLK, Q => 
                           n19991, QN => n8374);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n7417, CK => CLK, Q => 
                           n19989, QN => n8342);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n7416, CK => CLK, Q => 
                           n19987, QN => n8310);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n7415, CK => CLK, Q => 
                           n19985, QN => n8278);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n7414, CK => CLK, Q => 
                           n19983, QN => n8246);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n7413, CK => CLK, Q => 
                           n19981, QN => n8214);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n7412, CK => CLK, Q => 
                           n19979, QN => n8182);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n7411, CK => CLK, Q => 
                           n19977, QN => n8150);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n7410, CK => CLK, Q => 
                           n19976, QN => n8118);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n7409, CK => CLK, Q => 
                           n19974, QN => n8086);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n7408, CK => CLK, Q => 
                           n19973, QN => n8054);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n7407, CK => CLK, Q => 
                           n19972, QN => n8022);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n7406, CK => CLK, Q => 
                           n19970, QN => n7990);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n7405, CK => CLK, Q => 
                           n19968, QN => n7958);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n7404, CK => CLK, Q => 
                           n19966, QN => n7926);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n7403, CK => CLK, Q => 
                           n19964, QN => n7894);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n7402, CK => CLK, Q => 
                           n19962, QN => n7862);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n7401, CK => CLK, Q => 
                           n19960, QN => n7830);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n7400, CK => CLK, Q => 
                           n19958, QN => n7798);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n7399, CK => CLK, Q => n19956
                           , QN => n7766);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n7398, CK => CLK, Q => n19954
                           , QN => n7734);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n7397, CK => CLK, Q => n19952
                           , QN => n7702);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n7396, CK => CLK, Q => n19950
                           , QN => n7670);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n7395, CK => CLK, Q => n19948
                           , QN => n7638);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n7394, CK => CLK, Q => n19946
                           , QN => n7606);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n7393, CK => CLK, Q => n19944
                           , QN => n7574);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n7392, CK => CLK, Q => n19942
                           , QN => n7542);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n7391, CK => CLK, Q => n19940
                           , QN => n7510);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n7390, CK => CLK, Q => n19938
                           , QN => n7478);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n7349, CK => CLK, Q => n8526
                           , QN => n20211);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n7348, CK => CLK, Q => n8528
                           , QN => n20210);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n7347, CK => CLK, Q => n8530
                           , QN => n20209);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n7346, CK => CLK, Q => n8532
                           , QN => n20208);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n7345, CK => CLK, Q => n8534
                           , QN => n20207);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n7344, CK => CLK, Q => n8536
                           , QN => n20206);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n7343, CK => CLK, Q => n8538
                           , QN => n20205);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n7342, CK => CLK, Q => n8540
                           , QN => n20204);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n7341, CK => CLK, Q => n8542
                           , QN => n20203);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n7340, CK => CLK, Q => n8544
                           , QN => n20202);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n7339, CK => CLK, Q => n8546
                           , QN => n20201);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n7338, CK => CLK, Q => n8548
                           , QN => n20200);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n7337, CK => CLK, Q => n8550
                           , QN => n20199);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n7336, CK => CLK, Q => n8552
                           , QN => n20198);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n7335, CK => CLK, Q => n8554,
                           QN => n20197);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n7334, CK => CLK, Q => n8556,
                           QN => n20196);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n7333, CK => CLK, Q => n8558,
                           QN => n20195);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n7332, CK => CLK, Q => n8560,
                           QN => n20194);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n7331, CK => CLK, Q => n8562,
                           QN => n20193);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n7330, CK => CLK, Q => n8564,
                           QN => n20192);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n7329, CK => CLK, Q => n8566,
                           QN => n20191);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n7328, CK => CLK, Q => n8568,
                           QN => n20190);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n7327, CK => CLK, Q => n8570,
                           QN => n20189);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n7326, CK => CLK, Q => n8572,
                           QN => n20096);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n7317, CK => CLK, Q => n9734
                           , QN => n15239);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n7316, CK => CLK, Q => n9735
                           , QN => n15240);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n7315, CK => CLK, Q => n9736
                           , QN => n15241);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n7314, CK => CLK, Q => n9737
                           , QN => n15242);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n7313, CK => CLK, Q => n9738
                           , QN => n15243);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n7312, CK => CLK, Q => n9739
                           , QN => n15244);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n7311, CK => CLK, Q => n9740
                           , QN => n15245);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n7310, CK => CLK, Q => n9741
                           , QN => n15246);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n7309, CK => CLK, Q => n9742
                           , QN => n15247);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n7308, CK => CLK, Q => n9743
                           , QN => n15248);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n7307, CK => CLK, Q => n9744
                           , QN => n15249);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n7306, CK => CLK, Q => n9745
                           , QN => n15250);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n7305, CK => CLK, Q => n9746
                           , QN => n15251);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n7304, CK => CLK, Q => n9747
                           , QN => n15252);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n7303, CK => CLK, Q => n9748,
                           QN => n15253);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n7302, CK => CLK, Q => n9749,
                           QN => n15254);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n7301, CK => CLK, Q => n9750,
                           QN => n15255);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n7300, CK => CLK, Q => n9751,
                           QN => n15256);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n7299, CK => CLK, Q => n9752,
                           QN => n15257);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n7298, CK => CLK, Q => n9753,
                           QN => n15258);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n7297, CK => CLK, Q => n9754,
                           QN => n15259);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n7296, CK => CLK, Q => n9755,
                           QN => n15260);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n7295, CK => CLK, Q => n9756,
                           QN => n15261);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n7294, CK => CLK, Q => n9757,
                           QN => n15262);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n7285, CK => CLK, Q => n9766
                           , QN => n15274);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n7284, CK => CLK, Q => n9767
                           , QN => n15275);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n7283, CK => CLK, Q => n9768
                           , QN => n15276);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n7282, CK => CLK, Q => n9769
                           , QN => n15277);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n7281, CK => CLK, Q => n9770
                           , QN => n15278);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n7280, CK => CLK, Q => n9771
                           , QN => n15279);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n7279, CK => CLK, Q => n9772
                           , QN => n15280);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n7278, CK => CLK, Q => n9773
                           , QN => n15281);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n7277, CK => CLK, Q => n9774
                           , QN => n15282);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n7276, CK => CLK, Q => n9775
                           , QN => n15283);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n7275, CK => CLK, Q => n9776
                           , QN => n15284);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n7274, CK => CLK, Q => n9777
                           , QN => n15285);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n7273, CK => CLK, Q => n9778
                           , QN => n15286);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n7272, CK => CLK, Q => n9779
                           , QN => n15287);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n7271, CK => CLK, Q => n9780,
                           QN => n15288);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n7270, CK => CLK, Q => n9781,
                           QN => n15289);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n7269, CK => CLK, Q => n9782,
                           QN => n15290);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n7268, CK => CLK, Q => n9783,
                           QN => n15291);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n7267, CK => CLK, Q => n9784,
                           QN => n15292);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n7266, CK => CLK, Q => n9785,
                           QN => n15293);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n7265, CK => CLK, Q => n9786,
                           QN => n15294);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n7264, CK => CLK, Q => n9787,
                           QN => n15295);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n7263, CK => CLK, Q => n9788,
                           QN => n15296);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n7262, CK => CLK, Q => n9789,
                           QN => n15297);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n7253, CK => CLK, Q => n8527
                           , QN => n20188);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n7252, CK => CLK, Q => n8529
                           , QN => n20187);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n7251, CK => CLK, Q => n8531
                           , QN => n20186);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n7250, CK => CLK, Q => n8533
                           , QN => n20185);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n7249, CK => CLK, Q => n8535
                           , QN => n20184);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n7248, CK => CLK, Q => n8537
                           , QN => n20183);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n7247, CK => CLK, Q => n8539
                           , QN => n20182);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n7246, CK => CLK, Q => n8541
                           , QN => n20181);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n7245, CK => CLK, Q => n8543
                           , QN => n20180);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n7244, CK => CLK, Q => n8545
                           , QN => n20179);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n7243, CK => CLK, Q => n8547
                           , QN => n20178);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n7242, CK => CLK, Q => n8549
                           , QN => n20177);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n7241, CK => CLK, Q => n8551
                           , QN => n20176);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n7240, CK => CLK, Q => n8553
                           , QN => n20175);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n7239, CK => CLK, Q => n8555,
                           QN => n20174);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n7238, CK => CLK, Q => n8557,
                           QN => n20173);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n7237, CK => CLK, Q => n8559,
                           QN => n20172);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n7236, CK => CLK, Q => n8561,
                           QN => n20171);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n7235, CK => CLK, Q => n8563,
                           QN => n20170);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n7234, CK => CLK, Q => n8565,
                           QN => n20169);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n7233, CK => CLK, Q => n8567,
                           QN => n20168);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n7232, CK => CLK, Q => n8569,
                           QN => n20167);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n7231, CK => CLK, Q => n8571,
                           QN => n20166);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n7230, CK => CLK, Q => n8573,
                           QN => n15331);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n7221, CK => CLK, Q => n8975
                           , QN => n20045);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n7220, CK => CLK, Q => n8977
                           , QN => n20044);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n7219, CK => CLK, Q => n8979
                           , QN => n20043);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n7218, CK => CLK, Q => n8981
                           , QN => n20042);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n7217, CK => CLK, Q => n8983
                           , QN => n20041);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n7216, CK => CLK, Q => n8985
                           , QN => n20040);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n7215, CK => CLK, Q => n8987
                           , QN => n20039);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n7214, CK => CLK, Q => n8989
                           , QN => n20038);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n7213, CK => CLK, Q => n8991
                           , QN => n20037);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n7212, CK => CLK, Q => n8993
                           , QN => n20036);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n7211, CK => CLK, Q => n8995
                           , QN => n20035);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n7210, CK => CLK, Q => n8997
                           , QN => n20034);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n7209, CK => CLK, Q => n8999
                           , QN => n20033);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n7208, CK => CLK, Q => n9001
                           , QN => n20032);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n7207, CK => CLK, Q => n9003,
                           QN => n20031);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n7206, CK => CLK, Q => n9005,
                           QN => n20030);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n7205, CK => CLK, Q => n9007,
                           QN => n20029);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n7204, CK => CLK, Q => n9009,
                           QN => n20028);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n7203, CK => CLK, Q => n9011,
                           QN => n20027);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n7202, CK => CLK, Q => n9013,
                           QN => n20026);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n7201, CK => CLK, Q => n9015,
                           QN => n20025);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n7200, CK => CLK, Q => n9017,
                           QN => n20024);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n7199, CK => CLK, Q => n9019,
                           QN => n20023);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n7198, CK => CLK, Q => n9021,
                           QN => n15365);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n7189, CK => CLK, Q => n9116
                           , QN => n15377);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n7188, CK => CLK, Q => n9127
                           , QN => n15378);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n7187, CK => CLK, Q => n9138
                           , QN => n15379);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n7186, CK => CLK, Q => n9149
                           , QN => n15380);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n7185, CK => CLK, Q => n9160
                           , QN => n15381);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n7184, CK => CLK, Q => n9171
                           , QN => n15382);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n7183, CK => CLK, Q => n9182
                           , QN => n15383);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n7182, CK => CLK, Q => n9193
                           , QN => n15384);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n7181, CK => CLK, Q => n9204
                           , QN => n15385);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n7180, CK => CLK, Q => n9215
                           , QN => n15386);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n7179, CK => CLK, Q => n9226
                           , QN => n15387);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n7178, CK => CLK, Q => n9237
                           , QN => n15388);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n7177, CK => CLK, Q => n9248
                           , QN => n15389);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n7176, CK => CLK, Q => n9259
                           , QN => n15390);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n7175, CK => CLK, Q => n9270,
                           QN => n15391);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n7174, CK => CLK, Q => n9281,
                           QN => n15392);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n7173, CK => CLK, Q => n9292,
                           QN => n15393);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n7172, CK => CLK, Q => n9303,
                           QN => n15394);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n7171, CK => CLK, Q => n9314,
                           QN => n15395);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n7170, CK => CLK, Q => n9325,
                           QN => n15396);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n7169, CK => CLK, Q => n9336,
                           QN => n15397);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n7168, CK => CLK, Q => n9347,
                           QN => n15398);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n7167, CK => CLK, Q => n9358,
                           QN => n15399);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n7166, CK => CLK, Q => n9369,
                           QN => n15400);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n7157, CK => CLK, Q => n9120
                           , QN => n15412);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n7156, CK => CLK, Q => n9131
                           , QN => n15413);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n7155, CK => CLK, Q => n9142
                           , QN => n15414);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n7154, CK => CLK, Q => n9153
                           , QN => n15415);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n7153, CK => CLK, Q => n9164
                           , QN => n15416);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n7152, CK => CLK, Q => n9175
                           , QN => n15417);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n7151, CK => CLK, Q => n9186
                           , QN => n15418);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n7150, CK => CLK, Q => n9197
                           , QN => n15419);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n7149, CK => CLK, Q => n9208
                           , QN => n15420);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n7148, CK => CLK, Q => n9219
                           , QN => n15421);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n7147, CK => CLK, Q => n9230
                           , QN => n15422);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n7146, CK => CLK, Q => n9241
                           , QN => n15423);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n7145, CK => CLK, Q => n9252
                           , QN => n15424);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n7144, CK => CLK, Q => n9263
                           , QN => n15425);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n7143, CK => CLK, Q => n9274,
                           QN => n15426);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n7142, CK => CLK, Q => n9285,
                           QN => n15427);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n7141, CK => CLK, Q => n9296,
                           QN => n15428);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n7140, CK => CLK, Q => n9307,
                           QN => n15429);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n7139, CK => CLK, Q => n9318,
                           QN => n15430);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n7138, CK => CLK, Q => n9329,
                           QN => n15431);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n7137, CK => CLK, Q => n9340,
                           QN => n15432);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n7136, CK => CLK, Q => n9351,
                           QN => n15433);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n7135, CK => CLK, Q => n9362,
                           QN => n15434);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n7134, CK => CLK, Q => n9373,
                           QN => n15435);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n7125, CK => CLK, Q => 
                           n9574, QN => n15446);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n7124, CK => CLK, Q => 
                           n9575, QN => n15447);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n7123, CK => CLK, Q => 
                           n9576, QN => n15448);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n7122, CK => CLK, Q => 
                           n9577, QN => n15449);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n7121, CK => CLK, Q => 
                           n9578, QN => n15450);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n7120, CK => CLK, Q => 
                           n9579, QN => n15451);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n7119, CK => CLK, Q => 
                           n9580, QN => n15452);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n7118, CK => CLK, Q => 
                           n9581, QN => n15453);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n7117, CK => CLK, Q => 
                           n9582, QN => n15454);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n7116, CK => CLK, Q => 
                           n9583, QN => n15455);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n7115, CK => CLK, Q => 
                           n9584, QN => n15456);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n7114, CK => CLK, Q => 
                           n9585, QN => n15457);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n7113, CK => CLK, Q => 
                           n9586, QN => n15458);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n7112, CK => CLK, Q => 
                           n9587, QN => n15459);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n7111, CK => CLK, Q => n9588
                           , QN => n15460);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n7110, CK => CLK, Q => n9589
                           , QN => n15461);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n7109, CK => CLK, Q => n9590
                           , QN => n15462);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n7108, CK => CLK, Q => n9591
                           , QN => n15463);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n7107, CK => CLK, Q => n9592
                           , QN => n15464);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n7106, CK => CLK, Q => n9593
                           , QN => n15465);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n7105, CK => CLK, Q => n9594
                           , QN => n15466);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n7104, CK => CLK, Q => n9595
                           , QN => n15467);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n7103, CK => CLK, Q => n9596
                           , QN => n15468);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n7102, CK => CLK, Q => n9597
                           , QN => n15469);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n7093, CK => CLK, Q => 
                           n9414, QN => n15480);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n7092, CK => CLK, Q => 
                           n9415, QN => n15481);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n7091, CK => CLK, Q => 
                           n9416, QN => n15482);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n7090, CK => CLK, Q => 
                           n9417, QN => n15483);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n7089, CK => CLK, Q => 
                           n9418, QN => n15484);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n7088, CK => CLK, Q => 
                           n9419, QN => n15485);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n7087, CK => CLK, Q => 
                           n9420, QN => n15486);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n7086, CK => CLK, Q => 
                           n9421, QN => n15487);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n7085, CK => CLK, Q => 
                           n9422, QN => n15488);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n7084, CK => CLK, Q => 
                           n9423, QN => n15489);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n7083, CK => CLK, Q => 
                           n9424, QN => n15490);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n7082, CK => CLK, Q => 
                           n9425, QN => n15491);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n7081, CK => CLK, Q => 
                           n9426, QN => n15492);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n7080, CK => CLK, Q => 
                           n9427, QN => n15493);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n7079, CK => CLK, Q => n9428
                           , QN => n15494);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n7078, CK => CLK, Q => n9429
                           , QN => n15495);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n7077, CK => CLK, Q => n9430
                           , QN => n15496);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n7076, CK => CLK, Q => n9431
                           , QN => n15497);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n7075, CK => CLK, Q => n9432
                           , QN => n15498);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n7074, CK => CLK, Q => n9433
                           , QN => n15499);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n7073, CK => CLK, Q => n9434
                           , QN => n15500);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n7072, CK => CLK, Q => n9435
                           , QN => n15501);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n7071, CK => CLK, Q => n9436
                           , QN => n15502);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n7070, CK => CLK, Q => n9437
                           , QN => n15503);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n7061, CK => CLK, Q => 
                           n8668, QN => n20307);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n7060, CK => CLK, Q => 
                           n8679, QN => n20306);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n7059, CK => CLK, Q => 
                           n8690, QN => n20305);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n7058, CK => CLK, Q => 
                           n8701, QN => n20304);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n7057, CK => CLK, Q => 
                           n8712, QN => n20303);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n7056, CK => CLK, Q => 
                           n8723, QN => n20302);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n7055, CK => CLK, Q => 
                           n8734, QN => n20301);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n7054, CK => CLK, Q => 
                           n8745, QN => n20300);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n7053, CK => CLK, Q => 
                           n8756, QN => n20299);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n7052, CK => CLK, Q => 
                           n8767, QN => n20298);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n7051, CK => CLK, Q => 
                           n8778, QN => n20297);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n7050, CK => CLK, Q => 
                           n8789, QN => n20296);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n7049, CK => CLK, Q => 
                           n8800, QN => n20295);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n7048, CK => CLK, Q => 
                           n8811, QN => n20294);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n7047, CK => CLK, Q => n8822
                           , QN => n20293);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n7046, CK => CLK, Q => n8833
                           , QN => n20292);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n7045, CK => CLK, Q => n8844
                           , QN => n20291);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n7044, CK => CLK, Q => n8855
                           , QN => n20290);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n7043, CK => CLK, Q => n8866
                           , QN => n20289);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n7042, CK => CLK, Q => n8877
                           , QN => n20288);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n7041, CK => CLK, Q => n8888
                           , QN => n20287);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n7040, CK => CLK, Q => n8899
                           , QN => n20286);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n7039, CK => CLK, Q => n8910
                           , QN => n20285);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n7038, CK => CLK, Q => n8921
                           , QN => n20284);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n7029, CK => CLK, Q => 
                           n8672, QN => n20283);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n7028, CK => CLK, Q => 
                           n8683, QN => n20282);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n7027, CK => CLK, Q => 
                           n8694, QN => n20281);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n7026, CK => CLK, Q => 
                           n8705, QN => n20280);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n7025, CK => CLK, Q => 
                           n8716, QN => n20279);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n7024, CK => CLK, Q => 
                           n8727, QN => n20278);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n7023, CK => CLK, Q => 
                           n8738, QN => n20277);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n7022, CK => CLK, Q => 
                           n8749, QN => n20276);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n7021, CK => CLK, Q => 
                           n8760, QN => n20275);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n7020, CK => CLK, Q => 
                           n8771, QN => n20274);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n7019, CK => CLK, Q => 
                           n8782, QN => n20273);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n7018, CK => CLK, Q => 
                           n8793, QN => n20272);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n7017, CK => CLK, Q => 
                           n8804, QN => n20271);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n7016, CK => CLK, Q => 
                           n8815, QN => n20270);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n7015, CK => CLK, Q => n8826
                           , QN => n20269);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n7014, CK => CLK, Q => n8837
                           , QN => n20268);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n7013, CK => CLK, Q => n8848
                           , QN => n20267);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n7012, CK => CLK, Q => n8859
                           , QN => n20266);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n7011, CK => CLK, Q => n8870
                           , QN => n20265);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n7010, CK => CLK, Q => n8881
                           , QN => n20264);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n7009, CK => CLK, Q => n8892
                           , QN => n20263);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n7008, CK => CLK, Q => n8903
                           , QN => n20262);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n7007, CK => CLK, Q => n8914
                           , QN => n20261);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n7006, CK => CLK, Q => n8925
                           , QN => n20260);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n6997, CK => CLK, Q => 
                           n9382, QN => n15584);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n6996, CK => CLK, Q => 
                           n9383, QN => n15585);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n6995, CK => CLK, Q => 
                           n9384, QN => n15586);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n6994, CK => CLK, Q => 
                           n9385, QN => n15587);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n6993, CK => CLK, Q => 
                           n9386, QN => n15588);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n6992, CK => CLK, Q => 
                           n9387, QN => n15589);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n6991, CK => CLK, Q => 
                           n9388, QN => n15590);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n6990, CK => CLK, Q => 
                           n9389, QN => n15591);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n6989, CK => CLK, Q => 
                           n9390, QN => n15592);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n6988, CK => CLK, Q => 
                           n9391, QN => n15593);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n6987, CK => CLK, Q => 
                           n9392, QN => n15594);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n6986, CK => CLK, Q => 
                           n9393, QN => n15595);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n6985, CK => CLK, Q => 
                           n9394, QN => n15596);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n6984, CK => CLK, Q => 
                           n9395, QN => n15597);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n6983, CK => CLK, Q => n9396
                           , QN => n15598);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n6982, CK => CLK, Q => n9397
                           , QN => n15599);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n6981, CK => CLK, Q => n9398
                           , QN => n15600);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n6980, CK => CLK, Q => n9399
                           , QN => n15601);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n6979, CK => CLK, Q => n9400
                           , QN => n15602);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n6978, CK => CLK, Q => n9401
                           , QN => n15603);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n6977, CK => CLK, Q => n9402
                           , QN => n15604);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n6976, CK => CLK, Q => n9403
                           , QN => n15605);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n6975, CK => CLK, Q => n9404
                           , QN => n15606);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n6974, CK => CLK, Q => n9405
                           , QN => n15607);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n6965, CK => CLK, Q => 
                           n8934, QN => n20165);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n6964, CK => CLK, Q => 
                           n8935, QN => n20164);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n6963, CK => CLK, Q => 
                           n8936, QN => n20163);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n6962, CK => CLK, Q => 
                           n8937, QN => n20162);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n6961, CK => CLK, Q => 
                           n8938, QN => n20161);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n6960, CK => CLK, Q => 
                           n8939, QN => n20160);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n6959, CK => CLK, Q => 
                           n8940, QN => n20159);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n6958, CK => CLK, Q => 
                           n8941, QN => n20158);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n6957, CK => CLK, Q => 
                           n8942, QN => n20157);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n6956, CK => CLK, Q => 
                           n8943, QN => n20156);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n6955, CK => CLK, Q => 
                           n8944, QN => n20155);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n6954, CK => CLK, Q => 
                           n8945, QN => n20154);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n6953, CK => CLK, Q => 
                           n8946, QN => n20153);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n6952, CK => CLK, Q => 
                           n8947, QN => n20152);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n6951, CK => CLK, Q => n8948
                           , QN => n20151);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n6950, CK => CLK, Q => n8949
                           , QN => n20150);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n6949, CK => CLK, Q => n8950
                           , QN => n20149);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n6948, CK => CLK, Q => n8951
                           , QN => n20148);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n6947, CK => CLK, Q => n8952
                           , QN => n20147);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n6946, CK => CLK, Q => n8953
                           , QN => n20146);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n6945, CK => CLK, Q => n8954
                           , QN => n20145);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n6944, CK => CLK, Q => n8955
                           , QN => n20144);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n6943, CK => CLK, Q => n8956
                           , QN => n20143);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n6942, CK => CLK, Q => n8957
                           , QN => n15641);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n6933, CK => CLK, Q => 
                           n9115, QN => n15656);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n6932, CK => CLK, Q => 
                           n9126, QN => n15657);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n6931, CK => CLK, Q => 
                           n9137, QN => n15658);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n6930, CK => CLK, Q => 
                           n9148, QN => n15659);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n6929, CK => CLK, Q => 
                           n9159, QN => n15660);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n6928, CK => CLK, Q => 
                           n9170, QN => n15661);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n6927, CK => CLK, Q => 
                           n9181, QN => n15662);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n6926, CK => CLK, Q => 
                           n9192, QN => n15663);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n6925, CK => CLK, Q => 
                           n9203, QN => n15664);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n6924, CK => CLK, Q => 
                           n9214, QN => n15665);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n6923, CK => CLK, Q => 
                           n9225, QN => n15666);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n6922, CK => CLK, Q => 
                           n9236, QN => n15667);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n6921, CK => CLK, Q => 
                           n9247, QN => n15668);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n6920, CK => CLK, Q => 
                           n9258, QN => n15669);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n6919, CK => CLK, Q => n9269
                           , QN => n15670);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n6918, CK => CLK, Q => n9280
                           , QN => n15671);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n6917, CK => CLK, Q => n9291
                           , QN => n15672);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n6916, CK => CLK, Q => n9302
                           , QN => n15673);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n6915, CK => CLK, Q => n9313
                           , QN => n15674);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n6914, CK => CLK, Q => n9324
                           , QN => n15675);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n6913, CK => CLK, Q => n9335
                           , QN => n15676);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n6912, CK => CLK, Q => n9346
                           , QN => n15677);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n6911, CK => CLK, Q => n9357
                           , QN => n15678);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n6910, CK => CLK, Q => n9368
                           , QN => n15679);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n6901, CK => CLK, Q => 
                           n9119, QN => n15691);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n6900, CK => CLK, Q => 
                           n9130, QN => n15692);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n6899, CK => CLK, Q => 
                           n9141, QN => n15693);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n6898, CK => CLK, Q => 
                           n9152, QN => n15694);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n6897, CK => CLK, Q => 
                           n9163, QN => n15695);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n6896, CK => CLK, Q => 
                           n9174, QN => n15696);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n6895, CK => CLK, Q => 
                           n9185, QN => n15697);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n6894, CK => CLK, Q => 
                           n9196, QN => n15698);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n6893, CK => CLK, Q => 
                           n9207, QN => n15699);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n6892, CK => CLK, Q => 
                           n9218, QN => n15700);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n6891, CK => CLK, Q => 
                           n9229, QN => n15701);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n6890, CK => CLK, Q => 
                           n9240, QN => n15702);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n6889, CK => CLK, Q => 
                           n9251, QN => n15703);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n6888, CK => CLK, Q => 
                           n9262, QN => n15704);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n6887, CK => CLK, Q => n9273
                           , QN => n15705);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n6886, CK => CLK, Q => n9284
                           , QN => n15706);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n6885, CK => CLK, Q => n9295
                           , QN => n15707);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n6884, CK => CLK, Q => n9306
                           , QN => n15708);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n6883, CK => CLK, Q => n9317
                           , QN => n15709);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n6882, CK => CLK, Q => n9328
                           , QN => n15710);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n6881, CK => CLK, Q => n9339
                           , QN => n15711);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n6880, CK => CLK, Q => n9350
                           , QN => n15712);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n6879, CK => CLK, Q => n9361
                           , QN => n15713);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n6878, CK => CLK, Q => n9372
                           , QN => n15714);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n6869, CK => CLK, Q => 
                           n9446, QN => n20142);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n6868, CK => CLK, Q => 
                           n9447, QN => n20141);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n6867, CK => CLK, Q => 
                           n9448, QN => n20140);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n6866, CK => CLK, Q => 
                           n9449, QN => n20139);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n6865, CK => CLK, Q => 
                           n9450, QN => n20138);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n6864, CK => CLK, Q => 
                           n9451, QN => n20137);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n6863, CK => CLK, Q => 
                           n9452, QN => n20136);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n6862, CK => CLK, Q => 
                           n9453, QN => n20135);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n6861, CK => CLK, Q => 
                           n9454, QN => n20134);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n6860, CK => CLK, Q => 
                           n9455, QN => n20133);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n6859, CK => CLK, Q => 
                           n9456, QN => n20132);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n6858, CK => CLK, Q => 
                           n9457, QN => n20131);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n6857, CK => CLK, Q => 
                           n9458, QN => n20130);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n6856, CK => CLK, Q => 
                           n9459, QN => n20129);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n6855, CK => CLK, Q => n9460
                           , QN => n20128);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n6854, CK => CLK, Q => n9461
                           , QN => n20127);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n6853, CK => CLK, Q => n9462
                           , QN => n20126);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n6852, CK => CLK, Q => n9463
                           , QN => n20125);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n6851, CK => CLK, Q => n9464
                           , QN => n20124);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n6850, CK => CLK, Q => n9465
                           , QN => n20123);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n6849, CK => CLK, Q => n9466
                           , QN => n20122);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n6848, CK => CLK, Q => n9467
                           , QN => n20121);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n6847, CK => CLK, Q => n9468
                           , QN => n20120);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n6846, CK => CLK, Q => n9469
                           , QN => n15748);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n6845, CK => CLK, Q => 
                           n19768, QN => n5053);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n6844, CK => CLK, Q => 
                           n19766, QN => n5052);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n6843, CK => CLK, Q => 
                           n19780, QN => n5051);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n6842, CK => CLK, Q => 
                           n19779, QN => n5050);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n6841, CK => CLK, Q => 
                           n19778, QN => n5049);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n6840, CK => CLK, Q => 
                           n19776, QN => n5048);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n6839, CK => CLK, Q => 
                           n19774, QN => n5047);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n6838, CK => CLK, Q => 
                           n19772, QN => n5046);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n6837, CK => CLK, Q => 
                           n19685, QN => n5045);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n6836, CK => CLK, Q => 
                           n19684, QN => n5044);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n6835, CK => CLK, Q => 
                           n19762, QN => n5043);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n6834, CK => CLK, Q => 
                           n19761, QN => n5042);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n6833, CK => CLK, Q => 
                           n19760, QN => n5041);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n6832, CK => CLK, Q => 
                           n19758, QN => n5040);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n6831, CK => CLK, Q => 
                           n19756, QN => n5039);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n6830, CK => CLK, Q => 
                           n19754, QN => n5038);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n6829, CK => CLK, Q => 
                           n19752, QN => n5037);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n6828, CK => CLK, Q => 
                           n19750, QN => n5036);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n6827, CK => CLK, Q => 
                           n19748, QN => n5035);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n6826, CK => CLK, Q => 
                           n19746, QN => n5034);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n6825, CK => CLK, Q => 
                           n19744, QN => n5033);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n6824, CK => CLK, Q => 
                           n19742, QN => n5032);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n6823, CK => CLK, Q => 
                           n19740, QN => n5031);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n6822, CK => CLK, Q => 
                           n19738, QN => n5030);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n6821, CK => CLK, Q => 
                           n19736, QN => n5029);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n6820, CK => CLK, Q => 
                           n19734, QN => n5028);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n6819, CK => CLK, Q => 
                           n19732, QN => n5027);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n6818, CK => CLK, Q => 
                           n19730, QN => n5026);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n6817, CK => CLK, Q => 
                           n19728, QN => n5025);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n6816, CK => CLK, Q => 
                           n19726, QN => n5024);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n6815, CK => CLK, Q => 
                           n19724, QN => n5023);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n6814, CK => CLK, Q => 
                           n19999, QN => n5022);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n6805, CK => CLK, Q => 
                           n8667, QN => n15762);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n6804, CK => CLK, Q => 
                           n8678, QN => n15763);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n6803, CK => CLK, Q => 
                           n8689, QN => n15764);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n6802, CK => CLK, Q => 
                           n8700, QN => n15765);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n6801, CK => CLK, Q => 
                           n8711, QN => n15766);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n6800, CK => CLK, Q => 
                           n8722, QN => n15767);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n6799, CK => CLK, Q => 
                           n8733, QN => n15768);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n6798, CK => CLK, Q => 
                           n8744, QN => n15769);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n6797, CK => CLK, Q => 
                           n8755, QN => n15770);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n6796, CK => CLK, Q => 
                           n8766, QN => n15771);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n6795, CK => CLK, Q => 
                           n8777, QN => n15772);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n6794, CK => CLK, Q => 
                           n8788, QN => n15773);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n6793, CK => CLK, Q => 
                           n8799, QN => n15774);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n6792, CK => CLK, Q => 
                           n8810, QN => n15775);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n6791, CK => CLK, Q => n8821
                           , QN => n15776);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n6790, CK => CLK, Q => n8832
                           , QN => n15777);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n6789, CK => CLK, Q => n8843
                           , QN => n15778);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n6788, CK => CLK, Q => n8854
                           , QN => n15779);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n6787, CK => CLK, Q => n8865
                           , QN => n15780);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n6786, CK => CLK, Q => n8876
                           , QN => n15781);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n6785, CK => CLK, Q => n8887
                           , QN => n15782);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n6784, CK => CLK, Q => n8898
                           , QN => n15783);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n6783, CK => CLK, Q => n8909
                           , QN => n15784);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n6782, CK => CLK, Q => n8920
                           , QN => n15785);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n6773, CK => CLK, Q => 
                           n8671, QN => n15797);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n6772, CK => CLK, Q => 
                           n8682, QN => n15798);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n6771, CK => CLK, Q => 
                           n8693, QN => n15799);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n6770, CK => CLK, Q => 
                           n8704, QN => n15800);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n6769, CK => CLK, Q => 
                           n8715, QN => n15801);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n6768, CK => CLK, Q => 
                           n8726, QN => n15802);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n6767, CK => CLK, Q => 
                           n8737, QN => n15803);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n6766, CK => CLK, Q => 
                           n8748, QN => n15804);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n6765, CK => CLK, Q => 
                           n8759, QN => n15805);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n6764, CK => CLK, Q => 
                           n8770, QN => n15806);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n6763, CK => CLK, Q => 
                           n8781, QN => n15807);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n6762, CK => CLK, Q => 
                           n8792, QN => n15808);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n6761, CK => CLK, Q => 
                           n8803, QN => n15809);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n6760, CK => CLK, Q => 
                           n8814, QN => n15810);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n6759, CK => CLK, Q => n8825
                           , QN => n15811);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n6758, CK => CLK, Q => n8836
                           , QN => n15812);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n6757, CK => CLK, Q => n8847
                           , QN => n15813);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n6756, CK => CLK, Q => n8858
                           , QN => n15814);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n6755, CK => CLK, Q => n8869
                           , QN => n15815);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n6754, CK => CLK, Q => n8880
                           , QN => n15816);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n6753, CK => CLK, Q => n8891
                           , QN => n15817);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n6752, CK => CLK, Q => n8902
                           , QN => n15818);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n6751, CK => CLK, Q => n8913
                           , QN => n15819);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n6750, CK => CLK, Q => n8924
                           , QN => n15820);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n6741, CK => CLK, Q => 
                           n9478, QN => n15831);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n6740, CK => CLK, Q => 
                           n9479, QN => n15832);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n6739, CK => CLK, Q => 
                           n9480, QN => n15833);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n6738, CK => CLK, Q => 
                           n9481, QN => n15834);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n6737, CK => CLK, Q => 
                           n9482, QN => n15835);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n6736, CK => CLK, Q => 
                           n9483, QN => n15836);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           n9484, QN => n15837);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           n9485, QN => n15838);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => 
                           n9486, QN => n15839);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => 
                           n9487, QN => n15840);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => 
                           n9488, QN => n15841);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => 
                           n9489, QN => n15842);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n6729, CK => CLK, Q => 
                           n9490, QN => n15843);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n6728, CK => CLK, Q => 
                           n9491, QN => n15844);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n6727, CK => CLK, Q => n9492
                           , QN => n15845);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n6726, CK => CLK, Q => n9493
                           , QN => n15846);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n6725, CK => CLK, Q => n9494
                           , QN => n15847);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n6724, CK => CLK, Q => n9495
                           , QN => n15848);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n6723, CK => CLK, Q => n9496
                           , QN => n15849);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n6722, CK => CLK, Q => n9497
                           , QN => n15850);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n6721, CK => CLK, Q => n9498
                           , QN => n15851);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n6720, CK => CLK, Q => n9499
                           , QN => n15852);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n6719, CK => CLK, Q => n9500
                           , QN => n15853);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n6718, CK => CLK, Q => n9501
                           , QN => n15854);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n6685, CK => CLK, Q => 
                           n19873, QN => n8467);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n6684, CK => CLK, Q => 
                           n19871, QN => n8435);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n6683, CK => CLK, Q => 
                           n19869, QN => n8403);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n6682, CK => CLK, Q => 
                           n19867, QN => n8371);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n6681, CK => CLK, Q => 
                           n19865, QN => n8339);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n6680, CK => CLK, Q => 
                           n19863, QN => n8307);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n6679, CK => CLK, Q => 
                           n19861, QN => n8275);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n6678, CK => CLK, Q => 
                           n19859, QN => n8243);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n6677, CK => CLK, Q => 
                           n19857, QN => n8211);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n6676, CK => CLK, Q => 
                           n19855, QN => n8179);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n6675, CK => CLK, Q => 
                           n19853, QN => n8147);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n6674, CK => CLK, Q => 
                           n19688, QN => n8115);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n6673, CK => CLK, Q => 
                           n19851, QN => n8083);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n6672, CK => CLK, Q => 
                           n19849, QN => n8051);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n6671, CK => CLK, Q => 
                           n19847, QN => n8019);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n6670, CK => CLK, Q => 
                           n19845, QN => n7987);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n6669, CK => CLK, Q => 
                           n19843, QN => n7955);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n6668, CK => CLK, Q => 
                           n19841, QN => n7923);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n6667, CK => CLK, Q => 
                           n19839, QN => n7891);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n6666, CK => CLK, Q => 
                           n19837, QN => n7859);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n6665, CK => CLK, Q => 
                           n19835, QN => n7827);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n6664, CK => CLK, Q => 
                           n19833, QN => n7795);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n6663, CK => CLK, Q => 
                           n19831, QN => n7763);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n6662, CK => CLK, Q => 
                           n19829, QN => n7731);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n6661, CK => CLK, Q => 
                           n19827, QN => n7699);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n6660, CK => CLK, Q => 
                           n19825, QN => n7667);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n6659, CK => CLK, Q => 
                           n19823, QN => n7635);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n6658, CK => CLK, Q => 
                           n19821, QN => n7603);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n6657, CK => CLK, Q => 
                           n19819, QN => n7571);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n6656, CK => CLK, Q => 
                           n19817, QN => n7539);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n6655, CK => CLK, Q => 
                           n19815, QN => n7507);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n6654, CK => CLK, Q => 
                           n19813, QN => n7475);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n6653, CK => CLK, Q => 
                           n19874, QN => n8466);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n6652, CK => CLK, Q => 
                           n19872, QN => n8434);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n6651, CK => CLK, Q => 
                           n19870, QN => n8402);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n6650, CK => CLK, Q => 
                           n19868, QN => n8370);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n6649, CK => CLK, Q => 
                           n19866, QN => n8338);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n6648, CK => CLK, Q => 
                           n19864, QN => n8306);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n6647, CK => CLK, Q => 
                           n19862, QN => n8274);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n6646, CK => CLK, Q => 
                           n19860, QN => n8242);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n6645, CK => CLK, Q => 
                           n19858, QN => n8210);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n6644, CK => CLK, Q => 
                           n19856, QN => n8178);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n6643, CK => CLK, Q => 
                           n19854, QN => n8146);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n6642, CK => CLK, Q => 
                           n19680, QN => n8114);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n6641, CK => CLK, Q => 
                           n19852, QN => n8082);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n6640, CK => CLK, Q => 
                           n19850, QN => n8050);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n6639, CK => CLK, Q => 
                           n19848, QN => n8018);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n6638, CK => CLK, Q => 
                           n19846, QN => n7986);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n6637, CK => CLK, Q => 
                           n19844, QN => n7954);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n6636, CK => CLK, Q => 
                           n19842, QN => n7922);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n6635, CK => CLK, Q => 
                           n19840, QN => n7890);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n6634, CK => CLK, Q => 
                           n19838, QN => n7858);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n6633, CK => CLK, Q => 
                           n19836, QN => n7826);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n6632, CK => CLK, Q => 
                           n19834, QN => n7794);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n6631, CK => CLK, Q => 
                           n19832, QN => n7762);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n6630, CK => CLK, Q => 
                           n19830, QN => n7730);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n6629, CK => CLK, Q => 
                           n19828, QN => n7698);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n6628, CK => CLK, Q => 
                           n19826, QN => n7666);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n6627, CK => CLK, Q => 
                           n19824, QN => n7634);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n6626, CK => CLK, Q => 
                           n19822, QN => n7602);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n6625, CK => CLK, Q => 
                           n19820, QN => n7570);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n6624, CK => CLK, Q => 
                           n19818, QN => n7538);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n6623, CK => CLK, Q => 
                           n19816, QN => n7506);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n6622, CK => CLK, Q => 
                           n19814, QN => n7474);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n6613, CK => CLK, Q => 
                           n9638, QN => n15904);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n6612, CK => CLK, Q => 
                           n9639, QN => n15905);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n6611, CK => CLK, Q => 
                           n9640, QN => n15906);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n6610, CK => CLK, Q => 
                           n9641, QN => n15907);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n6609, CK => CLK, Q => 
                           n9642, QN => n15908);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n6608, CK => CLK, Q => 
                           n9643, QN => n15909);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n6607, CK => CLK, Q => 
                           n9644, QN => n15910);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n6606, CK => CLK, Q => 
                           n9645, QN => n15911);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n6605, CK => CLK, Q => 
                           n9646, QN => n15912);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n6604, CK => CLK, Q => 
                           n9647, QN => n15913);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n6603, CK => CLK, Q => 
                           n9648, QN => n15914);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n6602, CK => CLK, Q => 
                           n9649, QN => n15915);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n6601, CK => CLK, Q => 
                           n9650, QN => n15916);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n6600, CK => CLK, Q => 
                           n9651, QN => n15917);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n6599, CK => CLK, Q => n9652
                           , QN => n15918);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n6598, CK => CLK, Q => n9653
                           , QN => n15919);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n6597, CK => CLK, Q => n9654
                           , QN => n15920);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n6596, CK => CLK, Q => n9655
                           , QN => n15921);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n6595, CK => CLK, Q => n9656
                           , QN => n15922);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n6594, CK => CLK, Q => n9657
                           , QN => n15923);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n6593, CK => CLK, Q => n9658
                           , QN => n15924);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n6592, CK => CLK, Q => n9659
                           , QN => n15925);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n6591, CK => CLK, Q => n9660
                           , QN => n15926);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n6590, CK => CLK, Q => n9661
                           , QN => n15927);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n6549, CK => CLK, Q => 
                           n9798, QN => n20095);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n6548, CK => CLK, Q => 
                           n9799, QN => n20094);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n6547, CK => CLK, Q => 
                           n9800, QN => n20093);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n6546, CK => CLK, Q => 
                           n9801, QN => n20092);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n6545, CK => CLK, Q => 
                           n9802, QN => n20091);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n6544, CK => CLK, Q => 
                           n9803, QN => n20090);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n6543, CK => CLK, Q => 
                           n9804, QN => n20089);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n6542, CK => CLK, Q => 
                           n9805, QN => n20088);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n6541, CK => CLK, Q => 
                           n9806, QN => n20087);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n6540, CK => CLK, Q => 
                           n9807, QN => n20086);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n6539, CK => CLK, Q => 
                           n9808, QN => n20085);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n6538, CK => CLK, Q => 
                           n9809, QN => n20084);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n6537, CK => CLK, Q => 
                           n9810, QN => n20083);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n6536, CK => CLK, Q => 
                           n9811, QN => n20082);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n6535, CK => CLK, Q => n9812
                           , QN => n20081);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n6534, CK => CLK, Q => n9813
                           , QN => n20080);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n6533, CK => CLK, Q => n9814
                           , QN => n20079);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n6532, CK => CLK, Q => n9815
                           , QN => n20078);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n6531, CK => CLK, Q => n9816
                           , QN => n20077);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n6530, CK => CLK, Q => n9817
                           , QN => n20076);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n6529, CK => CLK, Q => n9818
                           , QN => n20075);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n6528, CK => CLK, Q => n9819
                           , QN => n20074);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n6527, CK => CLK, Q => n9820
                           , QN => n20073);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n6526, CK => CLK, Q => n9821
                           , QN => n20072);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n6517, CK => CLK, Q => 
                           n9830, QN => n20071);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n6516, CK => CLK, Q => 
                           n9831, QN => n20070);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n6515, CK => CLK, Q => 
                           n9832, QN => n20069);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n6514, CK => CLK, Q => 
                           n9833, QN => n20068);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n6513, CK => CLK, Q => 
                           n9834, QN => n20067);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n6512, CK => CLK, Q => 
                           n9835, QN => n20066);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n6511, CK => CLK, Q => 
                           n9836, QN => n20065);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n6510, CK => CLK, Q => 
                           n9837, QN => n20064);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n6509, CK => CLK, Q => 
                           n9838, QN => n20063);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n6508, CK => CLK, Q => 
                           n9839, QN => n20062);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n6507, CK => CLK, Q => 
                           n9840, QN => n20061);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n6506, CK => CLK, Q => 
                           n9841, QN => n20060);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n6505, CK => CLK, Q => 
                           n9842, QN => n20059);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n6504, CK => CLK, Q => 
                           n9843, QN => n20058);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n6503, CK => CLK, Q => n9844
                           , QN => n20057);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n6502, CK => CLK, Q => n9845
                           , QN => n20056);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n6501, CK => CLK, Q => n9846
                           , QN => n20055);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n6500, CK => CLK, Q => n9847
                           , QN => n20054);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n6499, CK => CLK, Q => n9848
                           , QN => n20053);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n6498, CK => CLK, Q => n9849
                           , QN => n20052);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n6497, CK => CLK, Q => n9850
                           , QN => n20051);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n6496, CK => CLK, Q => n9851
                           , QN => n20050);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n6495, CK => CLK, Q => n9852
                           , QN => n20049);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n6494, CK => CLK, Q => n9853
                           , QN => n20048);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n6485, CK => CLK, Q => 
                           n9542, QN => n16041);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n6484, CK => CLK, Q => 
                           n9543, QN => n16042);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n6483, CK => CLK, Q => 
                           n9544, QN => n16043);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n6482, CK => CLK, Q => 
                           n9545, QN => n16044);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n6481, CK => CLK, Q => 
                           n9546, QN => n16045);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n6480, CK => CLK, Q => 
                           n9547, QN => n16046);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n6479, CK => CLK, Q => 
                           n9548, QN => n16047);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n6478, CK => CLK, Q => 
                           n9549, QN => n16048);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n6477, CK => CLK, Q => 
                           n9550, QN => n16049);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n6476, CK => CLK, Q => 
                           n9551, QN => n16050);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n6475, CK => CLK, Q => 
                           n9552, QN => n16051);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n6474, CK => CLK, Q => 
                           n9553, QN => n16052);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n6473, CK => CLK, Q => 
                           n9554, QN => n16053);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n6472, CK => CLK, Q => 
                           n9555, QN => n16054);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n6471, CK => CLK, Q => n9556
                           , QN => n16055);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n6470, CK => CLK, Q => n9557
                           , QN => n16056);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n6469, CK => CLK, Q => n9558
                           , QN => n16057);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n6468, CK => CLK, Q => n9559
                           , QN => n16058);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n6467, CK => CLK, Q => n9560
                           , QN => n16059);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n6466, CK => CLK, Q => n9561
                           , QN => n16060);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n6465, CK => CLK, Q => n9562
                           , QN => n16061);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n6464, CK => CLK, Q => n9563
                           , QN => n16062);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n6463, CK => CLK, Q => n9564
                           , QN => n16063);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n6462, CK => CLK, Q => n9565
                           , QN => n16064);
   REGISTERS_reg_32_23_inst : DFF_X1 port map( D => n6421, CK => CLK, Q => 
                           n8665, QN => n16109);
   REGISTERS_reg_32_22_inst : DFF_X1 port map( D => n6420, CK => CLK, Q => 
                           n8676, QN => n16110);
   REGISTERS_reg_32_21_inst : DFF_X1 port map( D => n6419, CK => CLK, Q => 
                           n8687, QN => n16111);
   REGISTERS_reg_32_20_inst : DFF_X1 port map( D => n6418, CK => CLK, Q => 
                           n8698, QN => n16112);
   REGISTERS_reg_32_19_inst : DFF_X1 port map( D => n6417, CK => CLK, Q => 
                           n8709, QN => n16113);
   REGISTERS_reg_32_18_inst : DFF_X1 port map( D => n6416, CK => CLK, Q => 
                           n8720, QN => n16114);
   REGISTERS_reg_32_17_inst : DFF_X1 port map( D => n6415, CK => CLK, Q => 
                           n8731, QN => n16115);
   REGISTERS_reg_32_16_inst : DFF_X1 port map( D => n6414, CK => CLK, Q => 
                           n8742, QN => n16116);
   REGISTERS_reg_32_15_inst : DFF_X1 port map( D => n6413, CK => CLK, Q => 
                           n8753, QN => n16117);
   REGISTERS_reg_32_14_inst : DFF_X1 port map( D => n6412, CK => CLK, Q => 
                           n8764, QN => n16118);
   REGISTERS_reg_32_13_inst : DFF_X1 port map( D => n6411, CK => CLK, Q => 
                           n8775, QN => n16119);
   REGISTERS_reg_32_12_inst : DFF_X1 port map( D => n6410, CK => CLK, Q => 
                           n8786, QN => n16120);
   REGISTERS_reg_32_11_inst : DFF_X1 port map( D => n6409, CK => CLK, Q => 
                           n8797, QN => n16121);
   REGISTERS_reg_32_10_inst : DFF_X1 port map( D => n6408, CK => CLK, Q => 
                           n8808, QN => n16122);
   REGISTERS_reg_32_9_inst : DFF_X1 port map( D => n6407, CK => CLK, Q => n8819
                           , QN => n16123);
   REGISTERS_reg_32_8_inst : DFF_X1 port map( D => n6406, CK => CLK, Q => n8830
                           , QN => n16124);
   REGISTERS_reg_32_7_inst : DFF_X1 port map( D => n6405, CK => CLK, Q => n8841
                           , QN => n16125);
   REGISTERS_reg_32_6_inst : DFF_X1 port map( D => n6404, CK => CLK, Q => n8852
                           , QN => n16126);
   REGISTERS_reg_32_5_inst : DFF_X1 port map( D => n6403, CK => CLK, Q => n8863
                           , QN => n16127);
   REGISTERS_reg_32_4_inst : DFF_X1 port map( D => n6402, CK => CLK, Q => n8874
                           , QN => n16128);
   REGISTERS_reg_32_3_inst : DFF_X1 port map( D => n6401, CK => CLK, Q => n8885
                           , QN => n16129);
   REGISTERS_reg_32_2_inst : DFF_X1 port map( D => n6400, CK => CLK, Q => n8896
                           , QN => n16130);
   REGISTERS_reg_32_1_inst : DFF_X1 port map( D => n6399, CK => CLK, Q => n8907
                           , QN => n16131);
   REGISTERS_reg_32_0_inst : DFF_X1 port map( D => n6398, CK => CLK, Q => n8918
                           , QN => n16132);
   REGISTERS_reg_33_20_inst : DFF_X1 port map( D => n6386, CK => CLK, Q => 
                           n8702, QN => n16147);
   REGISTERS_reg_33_19_inst : DFF_X1 port map( D => n6385, CK => CLK, Q => 
                           n8713, QN => n16148);
   REGISTERS_reg_33_18_inst : DFF_X1 port map( D => n6384, CK => CLK, Q => 
                           n8724, QN => n16149);
   REGISTERS_reg_33_17_inst : DFF_X1 port map( D => n6383, CK => CLK, Q => 
                           n8735, QN => n16150);
   REGISTERS_reg_33_16_inst : DFF_X1 port map( D => n6382, CK => CLK, Q => 
                           n8746, QN => n16151);
   REGISTERS_reg_33_15_inst : DFF_X1 port map( D => n6381, CK => CLK, Q => 
                           n8757, QN => n16152);
   REGISTERS_reg_33_14_inst : DFF_X1 port map( D => n6380, CK => CLK, Q => 
                           n8768, QN => n16153);
   REGISTERS_reg_33_13_inst : DFF_X1 port map( D => n6379, CK => CLK, Q => 
                           n8779, QN => n16154);
   REGISTERS_reg_33_12_inst : DFF_X1 port map( D => n6378, CK => CLK, Q => 
                           n8790, QN => n16155);
   REGISTERS_reg_33_11_inst : DFF_X1 port map( D => n6377, CK => CLK, Q => 
                           n8801, QN => n16156);
   REGISTERS_reg_33_10_inst : DFF_X1 port map( D => n6376, CK => CLK, Q => 
                           n8812, QN => n16157);
   REGISTERS_reg_33_9_inst : DFF_X1 port map( D => n6375, CK => CLK, Q => n8823
                           , QN => n16158);
   REGISTERS_reg_33_8_inst : DFF_X1 port map( D => n6374, CK => CLK, Q => n8834
                           , QN => n16159);
   REGISTERS_reg_33_7_inst : DFF_X1 port map( D => n6373, CK => CLK, Q => n8845
                           , QN => n16160);
   REGISTERS_reg_33_6_inst : DFF_X1 port map( D => n6372, CK => CLK, Q => n8856
                           , QN => n16161);
   REGISTERS_reg_33_5_inst : DFF_X1 port map( D => n6371, CK => CLK, Q => n8867
                           , QN => n16162);
   REGISTERS_reg_33_4_inst : DFF_X1 port map( D => n6370, CK => CLK, Q => n8878
                           , QN => n16163);
   REGISTERS_reg_33_3_inst : DFF_X1 port map( D => n6369, CK => CLK, Q => n8889
                           , QN => n16164);
   REGISTERS_reg_33_2_inst : DFF_X1 port map( D => n6368, CK => CLK, Q => n8900
                           , QN => n16165);
   REGISTERS_reg_33_1_inst : DFF_X1 port map( D => n6367, CK => CLK, Q => n8911
                           , QN => n16166);
   REGISTERS_reg_33_0_inst : DFF_X1 port map( D => n6366, CK => CLK, Q => n8922
                           , QN => n16167);
   REGISTERS_reg_34_31_inst : DFF_X1 port map( D => n6365, CK => CLK, Q => 
                           n19767, QN => n4829);
   REGISTERS_reg_34_30_inst : DFF_X1 port map( D => n6364, CK => CLK, Q => 
                           n19765, QN => n4828);
   REGISTERS_reg_34_29_inst : DFF_X1 port map( D => n6363, CK => CLK, Q => 
                           n19764, QN => n4827);
   REGISTERS_reg_34_28_inst : DFF_X1 port map( D => n6362, CK => CLK, Q => 
                           n19763, QN => n4826);
   REGISTERS_reg_34_27_inst : DFF_X1 port map( D => n6361, CK => CLK, Q => 
                           n19777, QN => n4825);
   REGISTERS_reg_34_26_inst : DFF_X1 port map( D => n6360, CK => CLK, Q => 
                           n19775, QN => n4824);
   REGISTERS_reg_34_25_inst : DFF_X1 port map( D => n6359, CK => CLK, Q => 
                           n19773, QN => n4823);
   REGISTERS_reg_34_24_inst : DFF_X1 port map( D => n6358, CK => CLK, Q => 
                           n19771, QN => n4822);
   REGISTERS_reg_34_23_inst : DFF_X1 port map( D => n6357, CK => CLK, Q => 
                           n19770, QN => n4821);
   REGISTERS_reg_34_22_inst : DFF_X1 port map( D => n6356, CK => CLK, Q => 
                           n19769, QN => n4820);
   REGISTERS_reg_34_21_inst : DFF_X1 port map( D => n6355, CK => CLK, Q => 
                           n19683, QN => n4819);
   REGISTERS_reg_34_20_inst : DFF_X1 port map( D => n6354, CK => CLK, Q => 
                           n19682, QN => n4818);
   REGISTERS_reg_34_19_inst : DFF_X1 port map( D => n6353, CK => CLK, Q => 
                           n19759, QN => n4817);
   REGISTERS_reg_34_18_inst : DFF_X1 port map( D => n6352, CK => CLK, Q => 
                           n19757, QN => n4816);
   REGISTERS_reg_34_17_inst : DFF_X1 port map( D => n6351, CK => CLK, Q => 
                           n19755, QN => n4815);
   REGISTERS_reg_34_16_inst : DFF_X1 port map( D => n6350, CK => CLK, Q => 
                           n19753, QN => n4814);
   REGISTERS_reg_34_15_inst : DFF_X1 port map( D => n6349, CK => CLK, Q => 
                           n19751, QN => n4813);
   REGISTERS_reg_34_14_inst : DFF_X1 port map( D => n6348, CK => CLK, Q => 
                           n19749, QN => n4812);
   REGISTERS_reg_34_13_inst : DFF_X1 port map( D => n6347, CK => CLK, Q => 
                           n19747, QN => n4811);
   REGISTERS_reg_34_12_inst : DFF_X1 port map( D => n6346, CK => CLK, Q => 
                           n19745, QN => n4810);
   REGISTERS_reg_34_11_inst : DFF_X1 port map( D => n6345, CK => CLK, Q => 
                           n19743, QN => n4809);
   REGISTERS_reg_34_10_inst : DFF_X1 port map( D => n6344, CK => CLK, Q => 
                           n19741, QN => n4808);
   REGISTERS_reg_34_9_inst : DFF_X1 port map( D => n6343, CK => CLK, Q => 
                           n19739, QN => n4807);
   REGISTERS_reg_34_8_inst : DFF_X1 port map( D => n6342, CK => CLK, Q => 
                           n19737, QN => n4806);
   REGISTERS_reg_34_7_inst : DFF_X1 port map( D => n6341, CK => CLK, Q => 
                           n19735, QN => n4805);
   REGISTERS_reg_34_6_inst : DFF_X1 port map( D => n6340, CK => CLK, Q => 
                           n19733, QN => n4804);
   REGISTERS_reg_34_5_inst : DFF_X1 port map( D => n6339, CK => CLK, Q => 
                           n19731, QN => n4803);
   REGISTERS_reg_34_4_inst : DFF_X1 port map( D => n6338, CK => CLK, Q => 
                           n19729, QN => n4802);
   REGISTERS_reg_34_3_inst : DFF_X1 port map( D => n6337, CK => CLK, Q => 
                           n19727, QN => n4801);
   REGISTERS_reg_34_2_inst : DFF_X1 port map( D => n6336, CK => CLK, Q => 
                           n19725, QN => n4800);
   REGISTERS_reg_34_1_inst : DFF_X1 port map( D => n6335, CK => CLK, Q => 
                           n19723, QN => n4799);
   REGISTERS_reg_34_0_inst : DFF_X1 port map( D => n6334, CK => CLK, Q => 
                           n19812, QN => n4798);
   REGISTERS_reg_40_31_inst : DFF_X1 port map( D => n6173, CK => CLK, Q => 
                           n19933, QN => n8459);
   REGISTERS_reg_40_30_inst : DFF_X1 port map( D => n6172, CK => CLK, Q => 
                           n19931, QN => n8427);
   REGISTERS_reg_40_29_inst : DFF_X1 port map( D => n6171, CK => CLK, Q => 
                           n19929, QN => n8395);
   REGISTERS_reg_40_28_inst : DFF_X1 port map( D => n6170, CK => CLK, Q => 
                           n19927, QN => n8363);
   REGISTERS_reg_40_27_inst : DFF_X1 port map( D => n6169, CK => CLK, Q => 
                           n19925, QN => n8331);
   REGISTERS_reg_40_26_inst : DFF_X1 port map( D => n6168, CK => CLK, Q => 
                           n19923, QN => n8299);
   REGISTERS_reg_40_25_inst : DFF_X1 port map( D => n6167, CK => CLK, Q => 
                           n19921, QN => n8267);
   REGISTERS_reg_40_24_inst : DFF_X1 port map( D => n6166, CK => CLK, Q => 
                           n19919, QN => n8235);
   REGISTERS_reg_40_23_inst : DFF_X1 port map( D => n6165, CK => CLK, Q => 
                           n19917, QN => n8203);
   REGISTERS_reg_40_22_inst : DFF_X1 port map( D => n6164, CK => CLK, Q => 
                           n19915, QN => n8171);
   REGISTERS_reg_40_21_inst : DFF_X1 port map( D => n6163, CK => CLK, Q => 
                           n19936, QN => n8139);
   REGISTERS_reg_40_20_inst : DFF_X1 port map( D => n6162, CK => CLK, Q => 
                           n19689, QN => n8107);
   REGISTERS_reg_40_19_inst : DFF_X1 port map( D => n6161, CK => CLK, Q => 
                           n19687, QN => n8075);
   REGISTERS_reg_40_18_inst : DFF_X1 port map( D => n6160, CK => CLK, Q => 
                           n19935, QN => n8043);
   REGISTERS_reg_40_17_inst : DFF_X1 port map( D => n6159, CK => CLK, Q => 
                           n19909, QN => n8011);
   REGISTERS_reg_40_16_inst : DFF_X1 port map( D => n6158, CK => CLK, Q => 
                           n19907, QN => n7979);
   REGISTERS_reg_40_15_inst : DFF_X1 port map( D => n6157, CK => CLK, Q => 
                           n19905, QN => n7947);
   REGISTERS_reg_40_14_inst : DFF_X1 port map( D => n6156, CK => CLK, Q => 
                           n19903, QN => n7915);
   REGISTERS_reg_40_13_inst : DFF_X1 port map( D => n6155, CK => CLK, Q => 
                           n19901, QN => n7883);
   REGISTERS_reg_40_12_inst : DFF_X1 port map( D => n6154, CK => CLK, Q => 
                           n19899, QN => n7851);
   REGISTERS_reg_40_11_inst : DFF_X1 port map( D => n6153, CK => CLK, Q => 
                           n19897, QN => n7819);
   REGISTERS_reg_40_10_inst : DFF_X1 port map( D => n6152, CK => CLK, Q => 
                           n19895, QN => n7787);
   REGISTERS_reg_40_9_inst : DFF_X1 port map( D => n6151, CK => CLK, Q => 
                           n19893, QN => n7755);
   REGISTERS_reg_40_8_inst : DFF_X1 port map( D => n6150, CK => CLK, Q => 
                           n19891, QN => n7723);
   REGISTERS_reg_40_7_inst : DFF_X1 port map( D => n6149, CK => CLK, Q => 
                           n19889, QN => n7691);
   REGISTERS_reg_40_6_inst : DFF_X1 port map( D => n6148, CK => CLK, Q => 
                           n19887, QN => n7659);
   REGISTERS_reg_40_5_inst : DFF_X1 port map( D => n6147, CK => CLK, Q => 
                           n19885, QN => n7627);
   REGISTERS_reg_40_4_inst : DFF_X1 port map( D => n6146, CK => CLK, Q => 
                           n19883, QN => n7595);
   REGISTERS_reg_40_3_inst : DFF_X1 port map( D => n6145, CK => CLK, Q => 
                           n19881, QN => n7563);
   REGISTERS_reg_40_2_inst : DFF_X1 port map( D => n6144, CK => CLK, Q => 
                           n19879, QN => n7531);
   REGISTERS_reg_40_1_inst : DFF_X1 port map( D => n6143, CK => CLK, Q => 
                           n19877, QN => n7499);
   REGISTERS_reg_40_0_inst : DFF_X1 port map( D => n6142, CK => CLK, Q => 
                           n19875, QN => n7467);
   REGISTERS_reg_41_31_inst : DFF_X1 port map( D => n6141, CK => CLK, Q => 
                           n19934, QN => n8458);
   REGISTERS_reg_41_30_inst : DFF_X1 port map( D => n6140, CK => CLK, Q => 
                           n19932, QN => n8426);
   REGISTERS_reg_41_29_inst : DFF_X1 port map( D => n6139, CK => CLK, Q => 
                           n19930, QN => n8394);
   REGISTERS_reg_41_28_inst : DFF_X1 port map( D => n6138, CK => CLK, Q => 
                           n19928, QN => n8362);
   REGISTERS_reg_41_27_inst : DFF_X1 port map( D => n6137, CK => CLK, Q => 
                           n19926, QN => n8330);
   REGISTERS_reg_41_26_inst : DFF_X1 port map( D => n6136, CK => CLK, Q => 
                           n19924, QN => n8298);
   REGISTERS_reg_41_25_inst : DFF_X1 port map( D => n6135, CK => CLK, Q => 
                           n19922, QN => n8266);
   REGISTERS_reg_41_24_inst : DFF_X1 port map( D => n6134, CK => CLK, Q => 
                           n19920, QN => n8234);
   REGISTERS_reg_41_23_inst : DFF_X1 port map( D => n6133, CK => CLK, Q => 
                           n19918, QN => n8202);
   REGISTERS_reg_41_22_inst : DFF_X1 port map( D => n6132, CK => CLK, Q => 
                           n19916, QN => n8170);
   REGISTERS_reg_41_21_inst : DFF_X1 port map( D => n6131, CK => CLK, Q => 
                           n19914, QN => n8138);
   REGISTERS_reg_41_20_inst : DFF_X1 port map( D => n6130, CK => CLK, Q => 
                           n19913, QN => n8106);
   REGISTERS_reg_41_19_inst : DFF_X1 port map( D => n6129, CK => CLK, Q => 
                           n19912, QN => n8074);
   REGISTERS_reg_41_18_inst : DFF_X1 port map( D => n6128, CK => CLK, Q => 
                           n19911, QN => n8042);
   REGISTERS_reg_41_17_inst : DFF_X1 port map( D => n6127, CK => CLK, Q => 
                           n19910, QN => n8010);
   REGISTERS_reg_41_16_inst : DFF_X1 port map( D => n6126, CK => CLK, Q => 
                           n19908, QN => n7978);
   REGISTERS_reg_41_15_inst : DFF_X1 port map( D => n6125, CK => CLK, Q => 
                           n19906, QN => n7946);
   REGISTERS_reg_41_14_inst : DFF_X1 port map( D => n6124, CK => CLK, Q => 
                           n19904, QN => n7914);
   REGISTERS_reg_41_13_inst : DFF_X1 port map( D => n6123, CK => CLK, Q => 
                           n19902, QN => n7882);
   REGISTERS_reg_41_12_inst : DFF_X1 port map( D => n6122, CK => CLK, Q => 
                           n19900, QN => n7850);
   REGISTERS_reg_41_11_inst : DFF_X1 port map( D => n6121, CK => CLK, Q => 
                           n19898, QN => n7818);
   REGISTERS_reg_41_10_inst : DFF_X1 port map( D => n6120, CK => CLK, Q => 
                           n19896, QN => n7786);
   REGISTERS_reg_41_9_inst : DFF_X1 port map( D => n6119, CK => CLK, Q => 
                           n19894, QN => n7754);
   REGISTERS_reg_41_8_inst : DFF_X1 port map( D => n6118, CK => CLK, Q => 
                           n19892, QN => n7722);
   REGISTERS_reg_41_7_inst : DFF_X1 port map( D => n6117, CK => CLK, Q => 
                           n19890, QN => n7690);
   REGISTERS_reg_41_6_inst : DFF_X1 port map( D => n6116, CK => CLK, Q => 
                           n19888, QN => n7658);
   REGISTERS_reg_41_5_inst : DFF_X1 port map( D => n6115, CK => CLK, Q => 
                           n19886, QN => n7626);
   REGISTERS_reg_41_4_inst : DFF_X1 port map( D => n6114, CK => CLK, Q => 
                           n19884, QN => n7594);
   REGISTERS_reg_41_3_inst : DFF_X1 port map( D => n6113, CK => CLK, Q => 
                           n19882, QN => n7562);
   REGISTERS_reg_41_2_inst : DFF_X1 port map( D => n6112, CK => CLK, Q => 
                           n19880, QN => n7530);
   REGISTERS_reg_41_1_inst : DFF_X1 port map( D => n6111, CK => CLK, Q => 
                           n19878, QN => n7498);
   REGISTERS_reg_41_0_inst : DFF_X1 port map( D => n6110, CK => CLK, Q => 
                           n19876, QN => n7466);
   REGISTERS_reg_42_31_inst : DFF_X1 port map( D => n6109, CK => CLK, Q => 
                           n19722, QN => n4701);
   REGISTERS_reg_42_30_inst : DFF_X1 port map( D => n6108, CK => CLK, Q => 
                           n19721, QN => n4700);
   REGISTERS_reg_42_29_inst : DFF_X1 port map( D => n6107, CK => CLK, Q => 
                           n19720, QN => n4699);
   REGISTERS_reg_42_28_inst : DFF_X1 port map( D => n6106, CK => CLK, Q => 
                           n19719, QN => n4698);
   REGISTERS_reg_42_27_inst : DFF_X1 port map( D => n6105, CK => CLK, Q => 
                           n19718, QN => n4697);
   REGISTERS_reg_42_26_inst : DFF_X1 port map( D => n6104, CK => CLK, Q => 
                           n19717, QN => n4696);
   REGISTERS_reg_42_25_inst : DFF_X1 port map( D => n6103, CK => CLK, Q => 
                           n19716, QN => n4695);
   REGISTERS_reg_42_24_inst : DFF_X1 port map( D => n6102, CK => CLK, Q => 
                           n19715, QN => n4694);
   REGISTERS_reg_42_23_inst : DFF_X1 port map( D => n6101, CK => CLK, Q => 
                           n19714, QN => n4693);
   REGISTERS_reg_42_22_inst : DFF_X1 port map( D => n6100, CK => CLK, Q => 
                           n19713, QN => n4692);
   REGISTERS_reg_42_21_inst : DFF_X1 port map( D => n6099, CK => CLK, Q => 
                           n19681, QN => n4691);
   REGISTERS_reg_42_20_inst : DFF_X1 port map( D => n6098, CK => CLK, Q => 
                           n19712, QN => n4690);
   REGISTERS_reg_42_19_inst : DFF_X1 port map( D => n6097, CK => CLK, Q => 
                           n19711, QN => n4689);
   REGISTERS_reg_42_18_inst : DFF_X1 port map( D => n6096, CK => CLK, Q => 
                           n19710, QN => n4688);
   REGISTERS_reg_42_17_inst : DFF_X1 port map( D => n6095, CK => CLK, Q => 
                           n19709, QN => n4687);
   REGISTERS_reg_42_16_inst : DFF_X1 port map( D => n6094, CK => CLK, Q => 
                           n19708, QN => n4686);
   REGISTERS_reg_42_15_inst : DFF_X1 port map( D => n6093, CK => CLK, Q => 
                           n19707, QN => n4685);
   REGISTERS_reg_42_14_inst : DFF_X1 port map( D => n6092, CK => CLK, Q => 
                           n19706, QN => n4684);
   REGISTERS_reg_42_13_inst : DFF_X1 port map( D => n6091, CK => CLK, Q => 
                           n19705, QN => n4683);
   REGISTERS_reg_42_12_inst : DFF_X1 port map( D => n6090, CK => CLK, Q => 
                           n19704, QN => n4682);
   REGISTERS_reg_42_11_inst : DFF_X1 port map( D => n6089, CK => CLK, Q => 
                           n19703, QN => n4681);
   REGISTERS_reg_42_10_inst : DFF_X1 port map( D => n6088, CK => CLK, Q => 
                           n19702, QN => n4680);
   REGISTERS_reg_42_9_inst : DFF_X1 port map( D => n6087, CK => CLK, Q => 
                           n19701, QN => n4679);
   REGISTERS_reg_42_8_inst : DFF_X1 port map( D => n6086, CK => CLK, Q => 
                           n19700, QN => n4678);
   REGISTERS_reg_42_7_inst : DFF_X1 port map( D => n6085, CK => CLK, Q => 
                           n19699, QN => n4677);
   REGISTERS_reg_42_6_inst : DFF_X1 port map( D => n6084, CK => CLK, Q => 
                           n19698, QN => n4676);
   REGISTERS_reg_42_5_inst : DFF_X1 port map( D => n6083, CK => CLK, Q => 
                           n19697, QN => n4675);
   REGISTERS_reg_42_4_inst : DFF_X1 port map( D => n6082, CK => CLK, Q => 
                           n19696, QN => n4674);
   REGISTERS_reg_42_3_inst : DFF_X1 port map( D => n6081, CK => CLK, Q => 
                           n19695, QN => n4673);
   REGISTERS_reg_42_2_inst : DFF_X1 port map( D => n6080, CK => CLK, Q => 
                           n19694, QN => n4672);
   REGISTERS_reg_42_1_inst : DFF_X1 port map( D => n6079, CK => CLK, Q => 
                           n19693, QN => n4671);
   REGISTERS_reg_42_0_inst : DFF_X1 port map( D => n6078, CK => CLK, Q => 
                           n19692, QN => n4670);
   REGISTERS_reg_48_23_inst : DFF_X1 port map( D => n5909, CK => CLK, Q => 
                           n9958, QN => n16530);
   REGISTERS_reg_48_22_inst : DFF_X1 port map( D => n5908, CK => CLK, Q => 
                           n9959, QN => n16531);
   REGISTERS_reg_48_21_inst : DFF_X1 port map( D => n5907, CK => CLK, Q => 
                           n9960, QN => n16532);
   REGISTERS_reg_48_20_inst : DFF_X1 port map( D => n5906, CK => CLK, Q => 
                           n9961, QN => n16533);
   REGISTERS_reg_48_19_inst : DFF_X1 port map( D => n5905, CK => CLK, Q => 
                           n9962, QN => n16534);
   REGISTERS_reg_48_18_inst : DFF_X1 port map( D => n5904, CK => CLK, Q => 
                           n9963, QN => n16535);
   REGISTERS_reg_48_17_inst : DFF_X1 port map( D => n5903, CK => CLK, Q => 
                           n9964, QN => n16536);
   REGISTERS_reg_48_16_inst : DFF_X1 port map( D => n5902, CK => CLK, Q => 
                           n9965, QN => n16537);
   REGISTERS_reg_48_15_inst : DFF_X1 port map( D => n5901, CK => CLK, Q => 
                           n9966, QN => n16538);
   REGISTERS_reg_48_14_inst : DFF_X1 port map( D => n5900, CK => CLK, Q => 
                           n9967, QN => n16539);
   REGISTERS_reg_48_13_inst : DFF_X1 port map( D => n5899, CK => CLK, Q => 
                           n9968, QN => n16540);
   REGISTERS_reg_48_12_inst : DFF_X1 port map( D => n5898, CK => CLK, Q => 
                           n9969, QN => n16541);
   REGISTERS_reg_48_11_inst : DFF_X1 port map( D => n5897, CK => CLK, Q => 
                           n9970, QN => n16542);
   REGISTERS_reg_48_10_inst : DFF_X1 port map( D => n5896, CK => CLK, Q => 
                           n9971, QN => n16543);
   REGISTERS_reg_48_9_inst : DFF_X1 port map( D => n5895, CK => CLK, Q => n9972
                           , QN => n16544);
   REGISTERS_reg_48_8_inst : DFF_X1 port map( D => n5894, CK => CLK, Q => n9973
                           , QN => n16545);
   REGISTERS_reg_48_7_inst : DFF_X1 port map( D => n5893, CK => CLK, Q => n9974
                           , QN => n16546);
   REGISTERS_reg_48_6_inst : DFF_X1 port map( D => n5892, CK => CLK, Q => n9975
                           , QN => n16547);
   REGISTERS_reg_48_5_inst : DFF_X1 port map( D => n5891, CK => CLK, Q => n9976
                           , QN => n16548);
   REGISTERS_reg_48_4_inst : DFF_X1 port map( D => n5890, CK => CLK, Q => n9977
                           , QN => n16549);
   REGISTERS_reg_48_3_inst : DFF_X1 port map( D => n5889, CK => CLK, Q => n9978
                           , QN => n16550);
   REGISTERS_reg_48_2_inst : DFF_X1 port map( D => n5888, CK => CLK, Q => n9979
                           , QN => n16551);
   REGISTERS_reg_48_1_inst : DFF_X1 port map( D => n5887, CK => CLK, Q => n9980
                           , QN => n16552);
   REGISTERS_reg_48_0_inst : DFF_X1 port map( D => n5886, CK => CLK, Q => n9981
                           , QN => n16553);
   REGISTERS_reg_49_23_inst : DFF_X1 port map( D => n5877, CK => CLK, Q => 
                           n9990, QN => n16565);
   REGISTERS_reg_49_22_inst : DFF_X1 port map( D => n5876, CK => CLK, Q => 
                           n9991, QN => n16566);
   REGISTERS_reg_49_21_inst : DFF_X1 port map( D => n5875, CK => CLK, Q => 
                           n9992, QN => n16567);
   REGISTERS_reg_49_20_inst : DFF_X1 port map( D => n5874, CK => CLK, Q => 
                           n9993, QN => n16568);
   REGISTERS_reg_49_19_inst : DFF_X1 port map( D => n5873, CK => CLK, Q => 
                           n9994, QN => n16569);
   REGISTERS_reg_49_18_inst : DFF_X1 port map( D => n5872, CK => CLK, Q => 
                           n9995, QN => n16570);
   REGISTERS_reg_49_17_inst : DFF_X1 port map( D => n5871, CK => CLK, Q => 
                           n9996, QN => n16571);
   REGISTERS_reg_49_16_inst : DFF_X1 port map( D => n5870, CK => CLK, Q => 
                           n9997, QN => n16572);
   REGISTERS_reg_49_15_inst : DFF_X1 port map( D => n5869, CK => CLK, Q => 
                           n9998, QN => n16573);
   REGISTERS_reg_49_14_inst : DFF_X1 port map( D => n5868, CK => CLK, Q => 
                           n9999, QN => n16574);
   REGISTERS_reg_49_13_inst : DFF_X1 port map( D => n5867, CK => CLK, Q => 
                           n10000, QN => n7870);
   REGISTERS_reg_49_12_inst : DFF_X1 port map( D => n5866, CK => CLK, Q => 
                           n10001, QN => n7838);
   REGISTERS_reg_49_11_inst : DFF_X1 port map( D => n5865, CK => CLK, Q => 
                           n10002, QN => n7806);
   REGISTERS_reg_49_10_inst : DFF_X1 port map( D => n5864, CK => CLK, Q => 
                           n10003, QN => n7774);
   REGISTERS_reg_49_9_inst : DFF_X1 port map( D => n5863, CK => CLK, Q => 
                           n10004, QN => n7742);
   REGISTERS_reg_49_8_inst : DFF_X1 port map( D => n5862, CK => CLK, Q => 
                           n10005, QN => n7710);
   REGISTERS_reg_49_7_inst : DFF_X1 port map( D => n5861, CK => CLK, Q => 
                           n10006, QN => n7678);
   REGISTERS_reg_49_6_inst : DFF_X1 port map( D => n5860, CK => CLK, Q => 
                           n10007, QN => n7646);
   REGISTERS_reg_49_5_inst : DFF_X1 port map( D => n5859, CK => CLK, Q => 
                           n10008, QN => n7614);
   REGISTERS_reg_49_4_inst : DFF_X1 port map( D => n5858, CK => CLK, Q => 
                           n10009, QN => n7582);
   REGISTERS_reg_49_3_inst : DFF_X1 port map( D => n5857, CK => CLK, Q => 
                           n10010, QN => n7550);
   REGISTERS_reg_49_2_inst : DFF_X1 port map( D => n5856, CK => CLK, Q => 
                           n10011, QN => n7518);
   REGISTERS_reg_49_1_inst : DFF_X1 port map( D => n5855, CK => CLK, Q => 
                           n10012, QN => n7486);
   REGISTERS_reg_49_0_inst : DFF_X1 port map( D => n5854, CK => CLK, Q => 
                           n10013, QN => n7454);
   REGISTERS_reg_50_23_inst : DFF_X1 port map( D => n5845, CK => CLK, Q => 
                           n8486, QN => n20022);
   REGISTERS_reg_50_22_inst : DFF_X1 port map( D => n5844, CK => CLK, Q => 
                           n8487, QN => n20021);
   REGISTERS_reg_50_21_inst : DFF_X1 port map( D => n5843, CK => CLK, Q => 
                           n8488, QN => n20020);
   REGISTERS_reg_50_20_inst : DFF_X1 port map( D => n5842, CK => CLK, Q => 
                           n8489, QN => n20019);
   REGISTERS_reg_50_19_inst : DFF_X1 port map( D => n5841, CK => CLK, Q => 
                           n8490, QN => n20018);
   REGISTERS_reg_50_18_inst : DFF_X1 port map( D => n5840, CK => CLK, Q => 
                           n8491, QN => n20017);
   REGISTERS_reg_50_17_inst : DFF_X1 port map( D => n5839, CK => CLK, Q => 
                           n8492, QN => n20016);
   REGISTERS_reg_50_16_inst : DFF_X1 port map( D => n5838, CK => CLK, Q => 
                           n8493, QN => n20015);
   REGISTERS_reg_50_15_inst : DFF_X1 port map( D => n5837, CK => CLK, Q => 
                           n8494, QN => n20014);
   REGISTERS_reg_50_14_inst : DFF_X1 port map( D => n5836, CK => CLK, Q => 
                           n8495, QN => n20013);
   REGISTERS_reg_50_13_inst : DFF_X1 port map( D => n5835, CK => CLK, Q => 
                           n8496, QN => n20012);
   REGISTERS_reg_50_12_inst : DFF_X1 port map( D => n5834, CK => CLK, Q => 
                           n8497, QN => n20011);
   REGISTERS_reg_50_11_inst : DFF_X1 port map( D => n5833, CK => CLK, Q => 
                           n8498, QN => n20010);
   REGISTERS_reg_50_10_inst : DFF_X1 port map( D => n5832, CK => CLK, Q => 
                           n8499, QN => n20009);
   REGISTERS_reg_50_9_inst : DFF_X1 port map( D => n5831, CK => CLK, Q => n8500
                           , QN => n20008);
   REGISTERS_reg_50_8_inst : DFF_X1 port map( D => n5830, CK => CLK, Q => n8501
                           , QN => n20007);
   REGISTERS_reg_50_7_inst : DFF_X1 port map( D => n5829, CK => CLK, Q => n8502
                           , QN => n20006);
   REGISTERS_reg_50_6_inst : DFF_X1 port map( D => n5828, CK => CLK, Q => n8503
                           , QN => n20005);
   REGISTERS_reg_50_5_inst : DFF_X1 port map( D => n5827, CK => CLK, Q => n8504
                           , QN => n20004);
   REGISTERS_reg_50_4_inst : DFF_X1 port map( D => n5826, CK => CLK, Q => n8505
                           , QN => n20003);
   REGISTERS_reg_50_3_inst : DFF_X1 port map( D => n5825, CK => CLK, Q => n8506
                           , QN => n20002);
   REGISTERS_reg_50_2_inst : DFF_X1 port map( D => n5824, CK => CLK, Q => n8507
                           , QN => n20001);
   REGISTERS_reg_50_1_inst : DFF_X1 port map( D => n5823, CK => CLK, Q => n8508
                           , QN => n20000);
   REGISTERS_reg_50_0_inst : DFF_X1 port map( D => n5822, CK => CLK, Q => n8509
                           , QN => n16608);
   REGISTERS_reg_51_31_inst : DFF_X1 port map( D => n5821, CK => CLK, Q => 
                           n10398, QN => n4541);
   REGISTERS_reg_51_30_inst : DFF_X1 port map( D => n5820, CK => CLK, Q => 
                           n10399, QN => n4540);
   REGISTERS_reg_51_29_inst : DFF_X1 port map( D => n5819, CK => CLK, Q => 
                           n10400, QN => n4539);
   REGISTERS_reg_51_28_inst : DFF_X1 port map( D => n5818, CK => CLK, Q => 
                           n10401, QN => n4538);
   REGISTERS_reg_51_27_inst : DFF_X1 port map( D => n5817, CK => CLK, Q => 
                           n10402, QN => n4537);
   REGISTERS_reg_51_26_inst : DFF_X1 port map( D => n5816, CK => CLK, Q => 
                           n10403, QN => n4536);
   REGISTERS_reg_51_25_inst : DFF_X1 port map( D => n5815, CK => CLK, Q => 
                           n10404, QN => n4535);
   REGISTERS_reg_51_24_inst : DFF_X1 port map( D => n5814, CK => CLK, Q => 
                           n10405, QN => n4534);
   REGISTERS_reg_51_23_inst : DFF_X1 port map( D => n5813, CK => CLK, Q => 
                           n10406, QN => n4533);
   REGISTERS_reg_51_22_inst : DFF_X1 port map( D => n5812, CK => CLK, Q => 
                           n10407, QN => n4532);
   REGISTERS_reg_51_21_inst : DFF_X1 port map( D => n5811, CK => CLK, Q => 
                           n10408, QN => n4531);
   REGISTERS_reg_51_20_inst : DFF_X1 port map( D => n5810, CK => CLK, Q => 
                           n10409, QN => n4530);
   REGISTERS_reg_51_19_inst : DFF_X1 port map( D => n5809, CK => CLK, Q => 
                           n10410, QN => n4529);
   REGISTERS_reg_51_18_inst : DFF_X1 port map( D => n5808, CK => CLK, Q => 
                           n10411, QN => n4528);
   REGISTERS_reg_51_17_inst : DFF_X1 port map( D => n5807, CK => CLK, Q => 
                           n10412, QN => n4527);
   REGISTERS_reg_51_16_inst : DFF_X1 port map( D => n5806, CK => CLK, Q => 
                           n10413, QN => n4526);
   REGISTERS_reg_51_15_inst : DFF_X1 port map( D => n5805, CK => CLK, Q => 
                           n10414, QN => n4525);
   REGISTERS_reg_51_14_inst : DFF_X1 port map( D => n5804, CK => CLK, Q => 
                           n10415, QN => n4524);
   REGISTERS_reg_51_13_inst : DFF_X1 port map( D => n5803, CK => CLK, Q => 
                           n10416, QN => n4523);
   REGISTERS_reg_51_12_inst : DFF_X1 port map( D => n5802, CK => CLK, Q => 
                           n10417, QN => n4522);
   REGISTERS_reg_51_11_inst : DFF_X1 port map( D => n5801, CK => CLK, Q => 
                           n10418, QN => n4521);
   REGISTERS_reg_51_10_inst : DFF_X1 port map( D => n5800, CK => CLK, Q => 
                           n10419, QN => n4520);
   REGISTERS_reg_51_9_inst : DFF_X1 port map( D => n5799, CK => CLK, Q => 
                           n10420, QN => n4519);
   REGISTERS_reg_51_8_inst : DFF_X1 port map( D => n5798, CK => CLK, Q => 
                           n10421, QN => n4518);
   REGISTERS_reg_51_7_inst : DFF_X1 port map( D => n5797, CK => CLK, Q => 
                           n10422, QN => n4517);
   REGISTERS_reg_51_6_inst : DFF_X1 port map( D => n5796, CK => CLK, Q => 
                           n10423, QN => n4516);
   REGISTERS_reg_51_5_inst : DFF_X1 port map( D => n5795, CK => CLK, Q => 
                           n10424, QN => n4515);
   REGISTERS_reg_51_4_inst : DFF_X1 port map( D => n5794, CK => CLK, Q => 
                           n10425, QN => n4514);
   REGISTERS_reg_51_3_inst : DFF_X1 port map( D => n5793, CK => CLK, Q => 
                           n10426, QN => n4513);
   REGISTERS_reg_51_2_inst : DFF_X1 port map( D => n5792, CK => CLK, Q => 
                           n10427, QN => n4512);
   REGISTERS_reg_51_1_inst : DFF_X1 port map( D => n5791, CK => CLK, Q => 
                           n10428, QN => n4511);
   REGISTERS_reg_51_0_inst : DFF_X1 port map( D => n5790, CK => CLK, Q => 
                           n10429, QN => n4510);
   REGISTERS_reg_52_31_inst : DFF_X1 port map( D => n5789, CK => CLK, Q => 
                           n10430, QN => n8449);
   REGISTERS_reg_52_30_inst : DFF_X1 port map( D => n5788, CK => CLK, Q => 
                           n10431, QN => n8417);
   REGISTERS_reg_52_29_inst : DFF_X1 port map( D => n5787, CK => CLK, Q => 
                           n10432, QN => n8385);
   REGISTERS_reg_52_28_inst : DFF_X1 port map( D => n5786, CK => CLK, Q => 
                           n10433, QN => n8353);
   REGISTERS_reg_52_27_inst : DFF_X1 port map( D => n5785, CK => CLK, Q => 
                           n10434, QN => n8321);
   REGISTERS_reg_52_26_inst : DFF_X1 port map( D => n5784, CK => CLK, Q => 
                           n10435, QN => n8289);
   REGISTERS_reg_52_25_inst : DFF_X1 port map( D => n5783, CK => CLK, Q => 
                           n10436, QN => n8257);
   REGISTERS_reg_52_24_inst : DFF_X1 port map( D => n5782, CK => CLK, Q => 
                           n10437, QN => n8225);
   REGISTERS_reg_52_23_inst : DFF_X1 port map( D => n5781, CK => CLK, Q => 
                           n10438, QN => n8193);
   REGISTERS_reg_52_22_inst : DFF_X1 port map( D => n5780, CK => CLK, Q => 
                           n10439, QN => n8161);
   REGISTERS_reg_52_21_inst : DFF_X1 port map( D => n5779, CK => CLK, Q => 
                           n10440, QN => n8129);
   REGISTERS_reg_52_20_inst : DFF_X1 port map( D => n5778, CK => CLK, Q => 
                           n10441, QN => n8097);
   REGISTERS_reg_52_19_inst : DFF_X1 port map( D => n5777, CK => CLK, Q => 
                           n10442, QN => n8065);
   REGISTERS_reg_52_18_inst : DFF_X1 port map( D => n5776, CK => CLK, Q => 
                           n10443, QN => n8033);
   REGISTERS_reg_52_17_inst : DFF_X1 port map( D => n5775, CK => CLK, Q => 
                           n10444, QN => n8001);
   REGISTERS_reg_52_16_inst : DFF_X1 port map( D => n5774, CK => CLK, Q => 
                           n10445, QN => n7969);
   REGISTERS_reg_52_15_inst : DFF_X1 port map( D => n5773, CK => CLK, Q => 
                           n10446, QN => n7937);
   REGISTERS_reg_52_14_inst : DFF_X1 port map( D => n5772, CK => CLK, Q => 
                           n10447, QN => n7905);
   REGISTERS_reg_52_13_inst : DFF_X1 port map( D => n5771, CK => CLK, Q => 
                           n10448, QN => n7873);
   REGISTERS_reg_52_12_inst : DFF_X1 port map( D => n5770, CK => CLK, Q => 
                           n10449, QN => n7841);
   REGISTERS_reg_52_11_inst : DFF_X1 port map( D => n5769, CK => CLK, Q => 
                           n10450, QN => n7809);
   REGISTERS_reg_52_10_inst : DFF_X1 port map( D => n5768, CK => CLK, Q => 
                           n10451, QN => n7777);
   REGISTERS_reg_52_9_inst : DFF_X1 port map( D => n5767, CK => CLK, Q => 
                           n10452, QN => n7745);
   REGISTERS_reg_52_8_inst : DFF_X1 port map( D => n5766, CK => CLK, Q => 
                           n10453, QN => n7713);
   REGISTERS_reg_52_7_inst : DFF_X1 port map( D => n5765, CK => CLK, Q => 
                           n10454, QN => n7681);
   REGISTERS_reg_52_6_inst : DFF_X1 port map( D => n5764, CK => CLK, Q => 
                           n10455, QN => n7649);
   REGISTERS_reg_52_5_inst : DFF_X1 port map( D => n5763, CK => CLK, Q => 
                           n10456, QN => n7617);
   REGISTERS_reg_52_4_inst : DFF_X1 port map( D => n5762, CK => CLK, Q => 
                           n10457, QN => n7585);
   REGISTERS_reg_52_3_inst : DFF_X1 port map( D => n5761, CK => CLK, Q => 
                           n10458, QN => n7553);
   REGISTERS_reg_52_2_inst : DFF_X1 port map( D => n5760, CK => CLK, Q => 
                           n10459, QN => n7521);
   REGISTERS_reg_52_1_inst : DFF_X1 port map( D => n5759, CK => CLK, Q => 
                           n10460, QN => n7489);
   REGISTERS_reg_52_0_inst : DFF_X1 port map( D => n5758, CK => CLK, Q => 
                           n10461, QN => n7457);
   REGISTERS_reg_53_31_inst : DFF_X1 port map( D => n5757, CK => CLK, Q => 
                           n10462, QN => n8448);
   REGISTERS_reg_53_30_inst : DFF_X1 port map( D => n5756, CK => CLK, Q => 
                           n10463, QN => n8416);
   REGISTERS_reg_53_29_inst : DFF_X1 port map( D => n5755, CK => CLK, Q => 
                           n10464, QN => n8384);
   REGISTERS_reg_53_28_inst : DFF_X1 port map( D => n5754, CK => CLK, Q => 
                           n10465, QN => n8352);
   REGISTERS_reg_53_27_inst : DFF_X1 port map( D => n5753, CK => CLK, Q => 
                           n10466, QN => n8320);
   REGISTERS_reg_53_26_inst : DFF_X1 port map( D => n5752, CK => CLK, Q => 
                           n10467, QN => n8288);
   REGISTERS_reg_53_25_inst : DFF_X1 port map( D => n5751, CK => CLK, Q => 
                           n10468, QN => n8256);
   REGISTERS_reg_53_24_inst : DFF_X1 port map( D => n5750, CK => CLK, Q => 
                           n10469, QN => n8224);
   REGISTERS_reg_53_23_inst : DFF_X1 port map( D => n5749, CK => CLK, Q => 
                           n10470, QN => n8192);
   REGISTERS_reg_53_22_inst : DFF_X1 port map( D => n5748, CK => CLK, Q => 
                           n10471, QN => n8160);
   REGISTERS_reg_53_21_inst : DFF_X1 port map( D => n5747, CK => CLK, Q => 
                           n10472, QN => n8128);
   REGISTERS_reg_53_20_inst : DFF_X1 port map( D => n5746, CK => CLK, Q => 
                           n10473, QN => n8096);
   REGISTERS_reg_53_19_inst : DFF_X1 port map( D => n5745, CK => CLK, Q => 
                           n10474, QN => n8064);
   REGISTERS_reg_53_18_inst : DFF_X1 port map( D => n5744, CK => CLK, Q => 
                           n10475, QN => n8032);
   REGISTERS_reg_53_17_inst : DFF_X1 port map( D => n5743, CK => CLK, Q => 
                           n10476, QN => n8000);
   REGISTERS_reg_53_16_inst : DFF_X1 port map( D => n5742, CK => CLK, Q => 
                           n10477, QN => n7968);
   REGISTERS_reg_53_15_inst : DFF_X1 port map( D => n5741, CK => CLK, Q => 
                           n10478, QN => n7936);
   REGISTERS_reg_53_14_inst : DFF_X1 port map( D => n5740, CK => CLK, Q => 
                           n10479, QN => n7904);
   REGISTERS_reg_53_13_inst : DFF_X1 port map( D => n5739, CK => CLK, Q => 
                           n10480, QN => n7872);
   REGISTERS_reg_53_12_inst : DFF_X1 port map( D => n5738, CK => CLK, Q => 
                           n10481, QN => n7840);
   REGISTERS_reg_53_11_inst : DFF_X1 port map( D => n5737, CK => CLK, Q => 
                           n10482, QN => n7808);
   REGISTERS_reg_53_10_inst : DFF_X1 port map( D => n5736, CK => CLK, Q => 
                           n10483, QN => n7776);
   REGISTERS_reg_53_9_inst : DFF_X1 port map( D => n5735, CK => CLK, Q => 
                           n10484, QN => n7744);
   REGISTERS_reg_53_8_inst : DFF_X1 port map( D => n5734, CK => CLK, Q => 
                           n10485, QN => n7712);
   REGISTERS_reg_53_7_inst : DFF_X1 port map( D => n5733, CK => CLK, Q => 
                           n10486, QN => n7680);
   REGISTERS_reg_53_6_inst : DFF_X1 port map( D => n5732, CK => CLK, Q => 
                           n10487, QN => n7648);
   REGISTERS_reg_53_5_inst : DFF_X1 port map( D => n5731, CK => CLK, Q => 
                           n10488, QN => n7616);
   REGISTERS_reg_53_4_inst : DFF_X1 port map( D => n5730, CK => CLK, Q => 
                           n10489, QN => n7584);
   REGISTERS_reg_53_3_inst : DFF_X1 port map( D => n5729, CK => CLK, Q => 
                           n10490, QN => n7552);
   REGISTERS_reg_53_2_inst : DFF_X1 port map( D => n5728, CK => CLK, Q => 
                           n10491, QN => n7520);
   REGISTERS_reg_53_1_inst : DFF_X1 port map( D => n5727, CK => CLK, Q => 
                           n10492, QN => n7488);
   REGISTERS_reg_53_0_inst : DFF_X1 port map( D => n5726, CK => CLK, Q => 
                           n10493, QN => n7456);
   REGISTERS_reg_54_31_inst : DFF_X1 port map( D => n5725, CK => CLK, Q => 
                           n10014, QN => n4509);
   REGISTERS_reg_54_30_inst : DFF_X1 port map( D => n5724, CK => CLK, Q => 
                           n10015, QN => n4508);
   REGISTERS_reg_54_29_inst : DFF_X1 port map( D => n5723, CK => CLK, Q => 
                           n10016, QN => n4507);
   REGISTERS_reg_54_28_inst : DFF_X1 port map( D => n5722, CK => CLK, Q => 
                           n10017, QN => n4506);
   REGISTERS_reg_54_27_inst : DFF_X1 port map( D => n5721, CK => CLK, Q => 
                           n10018, QN => n4505);
   REGISTERS_reg_54_26_inst : DFF_X1 port map( D => n5720, CK => CLK, Q => 
                           n10019, QN => n4504);
   REGISTERS_reg_54_25_inst : DFF_X1 port map( D => n5719, CK => CLK, Q => 
                           n10020, QN => n4503);
   REGISTERS_reg_54_24_inst : DFF_X1 port map( D => n5718, CK => CLK, Q => 
                           n10021, QN => n4502);
   REGISTERS_reg_54_23_inst : DFF_X1 port map( D => n5717, CK => CLK, Q => 
                           n10022, QN => n4501);
   REGISTERS_reg_54_22_inst : DFF_X1 port map( D => n5716, CK => CLK, Q => 
                           n10023, QN => n4500);
   REGISTERS_reg_54_21_inst : DFF_X1 port map( D => n5715, CK => CLK, Q => 
                           n10024, QN => n4499);
   REGISTERS_reg_54_20_inst : DFF_X1 port map( D => n5714, CK => CLK, Q => 
                           n10025, QN => n4498);
   REGISTERS_reg_54_19_inst : DFF_X1 port map( D => n5713, CK => CLK, Q => 
                           n10026, QN => n4497);
   REGISTERS_reg_54_18_inst : DFF_X1 port map( D => n5712, CK => CLK, Q => 
                           n10027, QN => n4496);
   REGISTERS_reg_54_17_inst : DFF_X1 port map( D => n5711, CK => CLK, Q => 
                           n10028, QN => n4495);
   REGISTERS_reg_54_16_inst : DFF_X1 port map( D => n5710, CK => CLK, Q => 
                           n10029, QN => n4494);
   REGISTERS_reg_54_15_inst : DFF_X1 port map( D => n5709, CK => CLK, Q => 
                           n10030, QN => n4493);
   REGISTERS_reg_54_14_inst : DFF_X1 port map( D => n5708, CK => CLK, Q => 
                           n10031, QN => n4492);
   REGISTERS_reg_54_13_inst : DFF_X1 port map( D => n5707, CK => CLK, Q => 
                           n10032, QN => n4491);
   REGISTERS_reg_54_12_inst : DFF_X1 port map( D => n5706, CK => CLK, Q => 
                           n10033, QN => n4490);
   REGISTERS_reg_54_11_inst : DFF_X1 port map( D => n5705, CK => CLK, Q => 
                           n10034, QN => n4489);
   REGISTERS_reg_54_10_inst : DFF_X1 port map( D => n5704, CK => CLK, Q => 
                           n10035, QN => n4488);
   REGISTERS_reg_54_9_inst : DFF_X1 port map( D => n5703, CK => CLK, Q => 
                           n10036, QN => n4487);
   REGISTERS_reg_54_8_inst : DFF_X1 port map( D => n5702, CK => CLK, Q => 
                           n10037, QN => n4486);
   REGISTERS_reg_54_7_inst : DFF_X1 port map( D => n5701, CK => CLK, Q => 
                           n10038, QN => n4485);
   REGISTERS_reg_54_6_inst : DFF_X1 port map( D => n5700, CK => CLK, Q => 
                           n10039, QN => n4484);
   REGISTERS_reg_54_5_inst : DFF_X1 port map( D => n5699, CK => CLK, Q => 
                           n10040, QN => n4483);
   REGISTERS_reg_54_4_inst : DFF_X1 port map( D => n5698, CK => CLK, Q => 
                           n10041, QN => n4482);
   REGISTERS_reg_54_3_inst : DFF_X1 port map( D => n5697, CK => CLK, Q => 
                           n10042, QN => n4481);
   REGISTERS_reg_54_2_inst : DFF_X1 port map( D => n5696, CK => CLK, Q => 
                           n10043, QN => n4480);
   REGISTERS_reg_54_1_inst : DFF_X1 port map( D => n5695, CK => CLK, Q => 
                           n10044, QN => n4479);
   REGISTERS_reg_54_0_inst : DFF_X1 port map( D => n5694, CK => CLK, Q => 
                           n10045, QN => n4478);
   REGISTERS_reg_55_23_inst : DFF_X1 port map( D => n5685, CK => CLK, Q => 
                           n8664, QN => n20119);
   REGISTERS_reg_55_22_inst : DFF_X1 port map( D => n5684, CK => CLK, Q => 
                           n8675, QN => n20118);
   REGISTERS_reg_55_21_inst : DFF_X1 port map( D => n5683, CK => CLK, Q => 
                           n8686, QN => n20117);
   REGISTERS_reg_55_20_inst : DFF_X1 port map( D => n5682, CK => CLK, Q => 
                           n8697, QN => n20116);
   REGISTERS_reg_55_19_inst : DFF_X1 port map( D => n5681, CK => CLK, Q => 
                           n8708, QN => n20115);
   REGISTERS_reg_55_18_inst : DFF_X1 port map( D => n5680, CK => CLK, Q => 
                           n8719, QN => n20114);
   REGISTERS_reg_55_17_inst : DFF_X1 port map( D => n5679, CK => CLK, Q => 
                           n8730, QN => n20113);
   REGISTERS_reg_55_16_inst : DFF_X1 port map( D => n5678, CK => CLK, Q => 
                           n8741, QN => n20112);
   REGISTERS_reg_55_15_inst : DFF_X1 port map( D => n5677, CK => CLK, Q => 
                           n8752, QN => n20111);
   REGISTERS_reg_55_14_inst : DFF_X1 port map( D => n5676, CK => CLK, Q => 
                           n8763, QN => n20110);
   REGISTERS_reg_55_13_inst : DFF_X1 port map( D => n5675, CK => CLK, Q => 
                           n8774, QN => n20109);
   REGISTERS_reg_55_12_inst : DFF_X1 port map( D => n5674, CK => CLK, Q => 
                           n8785, QN => n20108);
   REGISTERS_reg_55_11_inst : DFF_X1 port map( D => n5673, CK => CLK, Q => 
                           n8796, QN => n20107);
   REGISTERS_reg_55_10_inst : DFF_X1 port map( D => n5672, CK => CLK, Q => 
                           n8807, QN => n20106);
   REGISTERS_reg_55_9_inst : DFF_X1 port map( D => n5671, CK => CLK, Q => n8818
                           , QN => n20105);
   REGISTERS_reg_55_8_inst : DFF_X1 port map( D => n5670, CK => CLK, Q => n8829
                           , QN => n20104);
   REGISTERS_reg_55_7_inst : DFF_X1 port map( D => n5669, CK => CLK, Q => n8840
                           , QN => n20103);
   REGISTERS_reg_55_6_inst : DFF_X1 port map( D => n5668, CK => CLK, Q => n8851
                           , QN => n20102);
   REGISTERS_reg_55_5_inst : DFF_X1 port map( D => n5667, CK => CLK, Q => n8862
                           , QN => n20101);
   REGISTERS_reg_55_4_inst : DFF_X1 port map( D => n5666, CK => CLK, Q => n8873
                           , QN => n20100);
   REGISTERS_reg_55_3_inst : DFF_X1 port map( D => n5665, CK => CLK, Q => n8884
                           , QN => n20099);
   REGISTERS_reg_55_2_inst : DFF_X1 port map( D => n5664, CK => CLK, Q => n8895
                           , QN => n20098);
   REGISTERS_reg_55_1_inst : DFF_X1 port map( D => n5663, CK => CLK, Q => n8906
                           , QN => n20097);
   REGISTERS_reg_55_0_inst : DFF_X1 port map( D => n5662, CK => CLK, Q => n8917
                           , QN => n16652);
   REGISTERS_reg_56_23_inst : DFF_X1 port map( D => n5653, CK => CLK, Q => 
                           n8666, QN => n20259);
   REGISTERS_reg_56_22_inst : DFF_X1 port map( D => n5652, CK => CLK, Q => 
                           n8677, QN => n20258);
   REGISTERS_reg_56_21_inst : DFF_X1 port map( D => n5651, CK => CLK, Q => 
                           n8688, QN => n20257);
   REGISTERS_reg_56_20_inst : DFF_X1 port map( D => n5650, CK => CLK, Q => 
                           n8699, QN => n20256);
   REGISTERS_reg_56_19_inst : DFF_X1 port map( D => n5649, CK => CLK, Q => 
                           n8710, QN => n20255);
   REGISTERS_reg_56_18_inst : DFF_X1 port map( D => n5648, CK => CLK, Q => 
                           n8721, QN => n20254);
   REGISTERS_reg_56_17_inst : DFF_X1 port map( D => n5647, CK => CLK, Q => 
                           n8732, QN => n20253);
   REGISTERS_reg_56_16_inst : DFF_X1 port map( D => n5646, CK => CLK, Q => 
                           n8743, QN => n20252);
   REGISTERS_reg_56_15_inst : DFF_X1 port map( D => n5645, CK => CLK, Q => 
                           n8754, QN => n20251);
   REGISTERS_reg_56_14_inst : DFF_X1 port map( D => n5644, CK => CLK, Q => 
                           n8765, QN => n20250);
   REGISTERS_reg_56_13_inst : DFF_X1 port map( D => n5643, CK => CLK, Q => 
                           n8776, QN => n20249);
   REGISTERS_reg_56_12_inst : DFF_X1 port map( D => n5642, CK => CLK, Q => 
                           n8787, QN => n20248);
   REGISTERS_reg_56_11_inst : DFF_X1 port map( D => n5641, CK => CLK, Q => 
                           n8798, QN => n20247);
   REGISTERS_reg_56_10_inst : DFF_X1 port map( D => n5640, CK => CLK, Q => 
                           n8809, QN => n20246);
   REGISTERS_reg_56_9_inst : DFF_X1 port map( D => n5639, CK => CLK, Q => n8820
                           , QN => n20245);
   REGISTERS_reg_56_8_inst : DFF_X1 port map( D => n5638, CK => CLK, Q => n8831
                           , QN => n20244);
   REGISTERS_reg_56_7_inst : DFF_X1 port map( D => n5637, CK => CLK, Q => n8842
                           , QN => n20243);
   REGISTERS_reg_56_6_inst : DFF_X1 port map( D => n5636, CK => CLK, Q => n8853
                           , QN => n20242);
   REGISTERS_reg_56_5_inst : DFF_X1 port map( D => n5635, CK => CLK, Q => n8864
                           , QN => n20241);
   REGISTERS_reg_56_4_inst : DFF_X1 port map( D => n5634, CK => CLK, Q => n8875
                           , QN => n20240);
   REGISTERS_reg_56_3_inst : DFF_X1 port map( D => n5633, CK => CLK, Q => n8886
                           , QN => n20239);
   REGISTERS_reg_56_2_inst : DFF_X1 port map( D => n5632, CK => CLK, Q => n8897
                           , QN => n20238);
   REGISTERS_reg_56_1_inst : DFF_X1 port map( D => n5631, CK => CLK, Q => n8908
                           , QN => n20237);
   REGISTERS_reg_56_0_inst : DFF_X1 port map( D => n5630, CK => CLK, Q => n8919
                           , QN => n20236);
   REGISTERS_reg_57_23_inst : DFF_X1 port map( D => n5621, CK => CLK, Q => 
                           n8670, QN => n20235);
   REGISTERS_reg_57_22_inst : DFF_X1 port map( D => n5620, CK => CLK, Q => 
                           n8681, QN => n20234);
   REGISTERS_reg_57_21_inst : DFF_X1 port map( D => n5619, CK => CLK, Q => 
                           n8692, QN => n20233);
   REGISTERS_reg_57_20_inst : DFF_X1 port map( D => n5618, CK => CLK, Q => 
                           n8703, QN => n20232);
   REGISTERS_reg_57_19_inst : DFF_X1 port map( D => n5617, CK => CLK, Q => 
                           n8714, QN => n20231);
   REGISTERS_reg_57_18_inst : DFF_X1 port map( D => n5616, CK => CLK, Q => 
                           n8725, QN => n20230);
   REGISTERS_reg_57_17_inst : DFF_X1 port map( D => n5615, CK => CLK, Q => 
                           n8736, QN => n20229);
   REGISTERS_reg_57_16_inst : DFF_X1 port map( D => n5614, CK => CLK, Q => 
                           n8747, QN => n20228);
   REGISTERS_reg_57_15_inst : DFF_X1 port map( D => n5613, CK => CLK, Q => 
                           n8758, QN => n20227);
   REGISTERS_reg_57_14_inst : DFF_X1 port map( D => n5612, CK => CLK, Q => 
                           n8769, QN => n20226);
   REGISTERS_reg_57_13_inst : DFF_X1 port map( D => n5611, CK => CLK, Q => 
                           n8780, QN => n20225);
   REGISTERS_reg_57_12_inst : DFF_X1 port map( D => n5610, CK => CLK, Q => 
                           n8791, QN => n20224);
   REGISTERS_reg_57_11_inst : DFF_X1 port map( D => n5609, CK => CLK, Q => 
                           n8802, QN => n20223);
   REGISTERS_reg_57_10_inst : DFF_X1 port map( D => n5608, CK => CLK, Q => 
                           n8813, QN => n20222);
   REGISTERS_reg_57_9_inst : DFF_X1 port map( D => n5607, CK => CLK, Q => n8824
                           , QN => n20221);
   REGISTERS_reg_57_8_inst : DFF_X1 port map( D => n5606, CK => CLK, Q => n8835
                           , QN => n20220);
   REGISTERS_reg_57_7_inst : DFF_X1 port map( D => n5605, CK => CLK, Q => n8846
                           , QN => n20219);
   REGISTERS_reg_57_6_inst : DFF_X1 port map( D => n5604, CK => CLK, Q => n8857
                           , QN => n20218);
   REGISTERS_reg_57_5_inst : DFF_X1 port map( D => n5603, CK => CLK, Q => n8868
                           , QN => n20217);
   REGISTERS_reg_57_4_inst : DFF_X1 port map( D => n5602, CK => CLK, Q => n8879
                           , QN => n20216);
   REGISTERS_reg_57_3_inst : DFF_X1 port map( D => n5601, CK => CLK, Q => n8890
                           , QN => n20215);
   REGISTERS_reg_57_2_inst : DFF_X1 port map( D => n5600, CK => CLK, Q => n8901
                           , QN => n20214);
   REGISTERS_reg_57_1_inst : DFF_X1 port map( D => n5599, CK => CLK, Q => n8912
                           , QN => n20213);
   REGISTERS_reg_57_0_inst : DFF_X1 port map( D => n5598, CK => CLK, Q => n8923
                           , QN => n20212);
   REGISTERS_reg_58_23_inst : DFF_X1 port map( D => n5589, CK => CLK, Q => 
                           n9112, QN => n16733);
   REGISTERS_reg_58_22_inst : DFF_X1 port map( D => n5588, CK => CLK, Q => 
                           n9123, QN => n16734);
   REGISTERS_reg_58_21_inst : DFF_X1 port map( D => n5587, CK => CLK, Q => 
                           n9134, QN => n16735);
   REGISTERS_reg_58_20_inst : DFF_X1 port map( D => n5586, CK => CLK, Q => 
                           n9145, QN => n16736);
   REGISTERS_reg_58_19_inst : DFF_X1 port map( D => n5585, CK => CLK, Q => 
                           n9156, QN => n16737);
   REGISTERS_reg_58_18_inst : DFF_X1 port map( D => n5584, CK => CLK, Q => 
                           n9167, QN => n16738);
   REGISTERS_reg_58_17_inst : DFF_X1 port map( D => n5583, CK => CLK, Q => 
                           n9178, QN => n16739);
   REGISTERS_reg_58_16_inst : DFF_X1 port map( D => n5582, CK => CLK, Q => 
                           n9189, QN => n16740);
   REGISTERS_reg_58_15_inst : DFF_X1 port map( D => n5581, CK => CLK, Q => 
                           n9200, QN => n16741);
   REGISTERS_reg_58_14_inst : DFF_X1 port map( D => n5580, CK => CLK, Q => 
                           n9211, QN => n16742);
   REGISTERS_reg_58_13_inst : DFF_X1 port map( D => n5579, CK => CLK, Q => 
                           n9222, QN => n16743);
   REGISTERS_reg_58_12_inst : DFF_X1 port map( D => n5578, CK => CLK, Q => 
                           n9233, QN => n16744);
   REGISTERS_reg_58_11_inst : DFF_X1 port map( D => n5577, CK => CLK, Q => 
                           n9244, QN => n16745);
   REGISTERS_reg_58_10_inst : DFF_X1 port map( D => n5576, CK => CLK, Q => 
                           n9255, QN => n16746);
   REGISTERS_reg_58_9_inst : DFF_X1 port map( D => n5575, CK => CLK, Q => n9266
                           , QN => n16747);
   REGISTERS_reg_58_8_inst : DFF_X1 port map( D => n5574, CK => CLK, Q => n9277
                           , QN => n16748);
   REGISTERS_reg_58_7_inst : DFF_X1 port map( D => n5573, CK => CLK, Q => n9288
                           , QN => n16749);
   REGISTERS_reg_58_6_inst : DFF_X1 port map( D => n5572, CK => CLK, Q => n9299
                           , QN => n16750);
   REGISTERS_reg_58_5_inst : DFF_X1 port map( D => n5571, CK => CLK, Q => n9310
                           , QN => n16751);
   REGISTERS_reg_58_4_inst : DFF_X1 port map( D => n5570, CK => CLK, Q => n9321
                           , QN => n16752);
   REGISTERS_reg_58_3_inst : DFF_X1 port map( D => n5569, CK => CLK, Q => n9332
                           , QN => n16753);
   REGISTERS_reg_58_2_inst : DFF_X1 port map( D => n5568, CK => CLK, Q => n9343
                           , QN => n16754);
   REGISTERS_reg_58_1_inst : DFF_X1 port map( D => n5567, CK => CLK, Q => n9354
                           , QN => n16755);
   REGISTERS_reg_58_0_inst : DFF_X1 port map( D => n5566, CK => CLK, Q => n9365
                           , QN => n16756);
   REGISTERS_reg_59_31_inst : DFF_X1 port map( D => n5565, CK => CLK, Q => 
                           n19810, QN => n4413);
   REGISTERS_reg_59_30_inst : DFF_X1 port map( D => n5564, CK => CLK, Q => 
                           n19809, QN => n4412);
   REGISTERS_reg_59_29_inst : DFF_X1 port map( D => n5563, CK => CLK, Q => 
                           n19808, QN => n4411);
   REGISTERS_reg_59_28_inst : DFF_X1 port map( D => n5562, CK => CLK, Q => 
                           n19807, QN => n4410);
   REGISTERS_reg_59_27_inst : DFF_X1 port map( D => n5561, CK => CLK, Q => 
                           n19806, QN => n4409);
   REGISTERS_reg_59_26_inst : DFF_X1 port map( D => n5560, CK => CLK, Q => 
                           n19805, QN => n4408);
   REGISTERS_reg_59_25_inst : DFF_X1 port map( D => n5559, CK => CLK, Q => 
                           n19804, QN => n4407);
   REGISTERS_reg_59_24_inst : DFF_X1 port map( D => n5558, CK => CLK, Q => 
                           n19803, QN => n4406);
   REGISTERS_reg_59_23_inst : DFF_X1 port map( D => n5557, CK => CLK, Q => 
                           n19802, QN => n4405);
   REGISTERS_reg_59_22_inst : DFF_X1 port map( D => n5556, CK => CLK, Q => 
                           n19801, QN => n4404);
   REGISTERS_reg_59_21_inst : DFF_X1 port map( D => n5555, CK => CLK, Q => 
                           n19686, QN => n4403);
   REGISTERS_reg_59_20_inst : DFF_X1 port map( D => n5554, CK => CLK, Q => 
                           n19800, QN => n4402);
   REGISTERS_reg_59_19_inst : DFF_X1 port map( D => n5553, CK => CLK, Q => 
                           n19799, QN => n4401);
   REGISTERS_reg_59_18_inst : DFF_X1 port map( D => n5552, CK => CLK, Q => 
                           n19798, QN => n4400);
   REGISTERS_reg_59_17_inst : DFF_X1 port map( D => n5551, CK => CLK, Q => 
                           n19797, QN => n4399);
   REGISTERS_reg_59_16_inst : DFF_X1 port map( D => n5550, CK => CLK, Q => 
                           n19796, QN => n4398);
   REGISTERS_reg_59_15_inst : DFF_X1 port map( D => n5549, CK => CLK, Q => 
                           n19795, QN => n4397);
   REGISTERS_reg_59_14_inst : DFF_X1 port map( D => n5548, CK => CLK, Q => 
                           n19794, QN => n4396);
   REGISTERS_reg_59_13_inst : DFF_X1 port map( D => n5547, CK => CLK, Q => 
                           n19793, QN => n4395);
   REGISTERS_reg_59_12_inst : DFF_X1 port map( D => n5546, CK => CLK, Q => 
                           n19792, QN => n4394);
   REGISTERS_reg_59_11_inst : DFF_X1 port map( D => n5545, CK => CLK, Q => 
                           n19791, QN => n4393);
   REGISTERS_reg_59_10_inst : DFF_X1 port map( D => n5544, CK => CLK, Q => 
                           n19790, QN => n4392);
   REGISTERS_reg_59_9_inst : DFF_X1 port map( D => n5543, CK => CLK, Q => 
                           n19789, QN => n4391);
   REGISTERS_reg_59_8_inst : DFF_X1 port map( D => n5542, CK => CLK, Q => 
                           n19788, QN => n4390);
   REGISTERS_reg_59_7_inst : DFF_X1 port map( D => n5541, CK => CLK, Q => 
                           n19787, QN => n4389);
   REGISTERS_reg_59_6_inst : DFF_X1 port map( D => n5540, CK => CLK, Q => 
                           n19786, QN => n4388);
   REGISTERS_reg_59_5_inst : DFF_X1 port map( D => n5539, CK => CLK, Q => 
                           n19785, QN => n4387);
   REGISTERS_reg_59_4_inst : DFF_X1 port map( D => n5538, CK => CLK, Q => 
                           n19784, QN => n4386);
   REGISTERS_reg_59_3_inst : DFF_X1 port map( D => n5537, CK => CLK, Q => 
                           n19783, QN => n4385);
   REGISTERS_reg_59_2_inst : DFF_X1 port map( D => n5536, CK => CLK, Q => 
                           n19782, QN => n4384);
   REGISTERS_reg_59_1_inst : DFF_X1 port map( D => n5535, CK => CLK, Q => 
                           n19781, QN => n4383);
   REGISTERS_reg_59_0_inst : DFF_X1 port map( D => n5534, CK => CLK, Q => 
                           n19811, QN => n4382);
   REGISTERS_reg_60_0_inst : DFF_X1 port map( D => n5502, CK => CLK, Q => n9367
                           , QN => n20047);
   REGISTERS_reg_61_0_inst : DFF_X1 port map( D => n5470, CK => CLK, Q => n9371
                           , QN => n20046);
   REGISTERS_reg_62_31_inst : DFF_X1 port map( D => n5469, CK => CLK, Q => 
                           n10046, QN => n4381);
   REGISTERS_reg_62_30_inst : DFF_X1 port map( D => n5468, CK => CLK, Q => 
                           n10047, QN => n4380);
   REGISTERS_reg_62_29_inst : DFF_X1 port map( D => n5467, CK => CLK, Q => 
                           n10048, QN => n4379);
   REGISTERS_reg_62_28_inst : DFF_X1 port map( D => n5466, CK => CLK, Q => 
                           n10049, QN => n4378);
   REGISTERS_reg_62_27_inst : DFF_X1 port map( D => n5465, CK => CLK, Q => 
                           n10050, QN => n4377);
   REGISTERS_reg_62_26_inst : DFF_X1 port map( D => n5464, CK => CLK, Q => 
                           n10051, QN => n4376);
   REGISTERS_reg_62_25_inst : DFF_X1 port map( D => n5463, CK => CLK, Q => 
                           n10052, QN => n4375);
   REGISTERS_reg_62_24_inst : DFF_X1 port map( D => n5462, CK => CLK, Q => 
                           n10053, QN => n4374);
   REGISTERS_reg_62_23_inst : DFF_X1 port map( D => n5461, CK => CLK, Q => 
                           n10054, QN => n4373);
   REGISTERS_reg_62_22_inst : DFF_X1 port map( D => n5460, CK => CLK, Q => 
                           n10055, QN => n4372);
   REGISTERS_reg_62_21_inst : DFF_X1 port map( D => n5459, CK => CLK, Q => 
                           n10056, QN => n4371);
   REGISTERS_reg_62_20_inst : DFF_X1 port map( D => n5458, CK => CLK, Q => 
                           n10057, QN => n4370);
   REGISTERS_reg_62_19_inst : DFF_X1 port map( D => n5457, CK => CLK, Q => 
                           n10058, QN => n4369);
   REGISTERS_reg_62_18_inst : DFF_X1 port map( D => n5456, CK => CLK, Q => 
                           n10059, QN => n4368);
   REGISTERS_reg_62_17_inst : DFF_X1 port map( D => n5455, CK => CLK, Q => 
                           n10060, QN => n4367);
   REGISTERS_reg_62_16_inst : DFF_X1 port map( D => n5454, CK => CLK, Q => 
                           n10061, QN => n4366);
   REGISTERS_reg_62_15_inst : DFF_X1 port map( D => n5453, CK => CLK, Q => 
                           n10062, QN => n4365);
   REGISTERS_reg_62_14_inst : DFF_X1 port map( D => n5452, CK => CLK, Q => 
                           n10063, QN => n4364);
   REGISTERS_reg_62_13_inst : DFF_X1 port map( D => n5451, CK => CLK, Q => 
                           n10064, QN => n4363);
   REGISTERS_reg_62_12_inst : DFF_X1 port map( D => n5450, CK => CLK, Q => 
                           n10065, QN => n4362);
   REGISTERS_reg_62_11_inst : DFF_X1 port map( D => n5449, CK => CLK, Q => 
                           n10066, QN => n4361);
   REGISTERS_reg_62_10_inst : DFF_X1 port map( D => n5448, CK => CLK, Q => 
                           n10067, QN => n4360);
   REGISTERS_reg_62_9_inst : DFF_X1 port map( D => n5447, CK => CLK, Q => 
                           n10068, QN => n4359);
   REGISTERS_reg_62_8_inst : DFF_X1 port map( D => n5446, CK => CLK, Q => 
                           n10069, QN => n4358);
   REGISTERS_reg_62_7_inst : DFF_X1 port map( D => n5445, CK => CLK, Q => 
                           n10070, QN => n4357);
   REGISTERS_reg_62_6_inst : DFF_X1 port map( D => n5444, CK => CLK, Q => 
                           n10071, QN => n4356);
   REGISTERS_reg_62_5_inst : DFF_X1 port map( D => n5443, CK => CLK, Q => 
                           n10072, QN => n4355);
   REGISTERS_reg_62_4_inst : DFF_X1 port map( D => n5442, CK => CLK, Q => 
                           n10073, QN => n4354);
   REGISTERS_reg_62_3_inst : DFF_X1 port map( D => n5441, CK => CLK, Q => 
                           n10074, QN => n4353);
   REGISTERS_reg_62_2_inst : DFF_X1 port map( D => n5440, CK => CLK, Q => 
                           n10075, QN => n4352);
   REGISTERS_reg_62_1_inst : DFF_X1 port map( D => n5439, CK => CLK, Q => 
                           n10076, QN => n4351);
   REGISTERS_reg_62_0_inst : DFF_X1 port map( D => n5438, CK => CLK, Q => 
                           n10077, QN => n4350);
   REGISTERS_reg_63_31_inst : DFF_X1 port map( D => n5437, CK => CLK, Q => 
                           n10078, QN => n4349);
   OUT2_reg_31_inst : DFF_X1 port map( D => n5436, CK => CLK, Q => OUT2(31), QN
                           => n4348);
   REGISTERS_reg_63_30_inst : DFF_X1 port map( D => n5435, CK => CLK, Q => 
                           n10079, QN => n4347);
   OUT2_reg_30_inst : DFF_X1 port map( D => n5434, CK => CLK, Q => OUT2(30), QN
                           => n4346);
   REGISTERS_reg_63_29_inst : DFF_X1 port map( D => n5433, CK => CLK, Q => 
                           n10080, QN => n4345);
   OUT2_reg_29_inst : DFF_X1 port map( D => n5432, CK => CLK, Q => OUT2(29), QN
                           => n4344);
   REGISTERS_reg_63_28_inst : DFF_X1 port map( D => n5431, CK => CLK, Q => 
                           n10081, QN => n4343);
   OUT2_reg_28_inst : DFF_X1 port map( D => n5430, CK => CLK, Q => OUT2(28), QN
                           => n4342);
   REGISTERS_reg_63_27_inst : DFF_X1 port map( D => n5429, CK => CLK, Q => 
                           n10082, QN => n4341);
   OUT2_reg_27_inst : DFF_X1 port map( D => n5428, CK => CLK, Q => OUT2(27), QN
                           => n4340);
   REGISTERS_reg_63_26_inst : DFF_X1 port map( D => n5427, CK => CLK, Q => 
                           n10083, QN => n4339);
   OUT2_reg_26_inst : DFF_X1 port map( D => n5426, CK => CLK, Q => OUT2(26), QN
                           => n4338);
   REGISTERS_reg_63_25_inst : DFF_X1 port map( D => n5425, CK => CLK, Q => 
                           n10084, QN => n4337);
   OUT2_reg_25_inst : DFF_X1 port map( D => n5424, CK => CLK, Q => OUT2(25), QN
                           => n4336);
   REGISTERS_reg_63_24_inst : DFF_X1 port map( D => n5423, CK => CLK, Q => 
                           n10085, QN => n4335);
   OUT2_reg_24_inst : DFF_X1 port map( D => n5422, CK => CLK, Q => OUT2(24), QN
                           => n4334);
   REGISTERS_reg_63_23_inst : DFF_X1 port map( D => n5421, CK => CLK, Q => 
                           n10086, QN => n4333);
   OUT2_reg_23_inst : DFF_X1 port map( D => n5420, CK => CLK, Q => OUT2(23), QN
                           => n4332);
   REGISTERS_reg_63_22_inst : DFF_X1 port map( D => n5419, CK => CLK, Q => 
                           n10087, QN => n4331);
   OUT2_reg_22_inst : DFF_X1 port map( D => n5418, CK => CLK, Q => OUT2(22), QN
                           => n4330);
   REGISTERS_reg_63_21_inst : DFF_X1 port map( D => n5417, CK => CLK, Q => 
                           n10088, QN => n4329);
   OUT2_reg_21_inst : DFF_X1 port map( D => n5416, CK => CLK, Q => OUT2(21), QN
                           => n4328);
   REGISTERS_reg_63_20_inst : DFF_X1 port map( D => n5415, CK => CLK, Q => 
                           n10089, QN => n4327);
   OUT2_reg_20_inst : DFF_X1 port map( D => n5414, CK => CLK, Q => OUT2(20), QN
                           => n4326);
   REGISTERS_reg_63_19_inst : DFF_X1 port map( D => n5413, CK => CLK, Q => 
                           n10090, QN => n4325);
   OUT2_reg_19_inst : DFF_X1 port map( D => n5412, CK => CLK, Q => OUT2(19), QN
                           => n4324);
   REGISTERS_reg_63_18_inst : DFF_X1 port map( D => n5411, CK => CLK, Q => 
                           n10091, QN => n4323);
   OUT2_reg_18_inst : DFF_X1 port map( D => n5410, CK => CLK, Q => OUT2(18), QN
                           => n4322);
   REGISTERS_reg_63_17_inst : DFF_X1 port map( D => n5409, CK => CLK, Q => 
                           n10092, QN => n4321);
   OUT2_reg_17_inst : DFF_X1 port map( D => n5408, CK => CLK, Q => OUT2(17), QN
                           => n4320);
   REGISTERS_reg_63_16_inst : DFF_X1 port map( D => n5407, CK => CLK, Q => 
                           n10093, QN => n4319);
   OUT2_reg_16_inst : DFF_X1 port map( D => n5406, CK => CLK, Q => OUT2(16), QN
                           => n4318);
   REGISTERS_reg_63_15_inst : DFF_X1 port map( D => n5405, CK => CLK, Q => 
                           n10094, QN => n4317);
   OUT2_reg_15_inst : DFF_X1 port map( D => n5404, CK => CLK, Q => OUT2(15), QN
                           => n4316);
   REGISTERS_reg_63_14_inst : DFF_X1 port map( D => n5403, CK => CLK, Q => 
                           n10095, QN => n4315);
   OUT2_reg_14_inst : DFF_X1 port map( D => n5402, CK => CLK, Q => OUT2(14), QN
                           => n4314);
   REGISTERS_reg_63_13_inst : DFF_X1 port map( D => n5401, CK => CLK, Q => 
                           n10096, QN => n4313);
   OUT2_reg_13_inst : DFF_X1 port map( D => n5400, CK => CLK, Q => OUT2(13), QN
                           => n4312);
   REGISTERS_reg_63_12_inst : DFF_X1 port map( D => n5399, CK => CLK, Q => 
                           n10097, QN => n4311);
   OUT2_reg_12_inst : DFF_X1 port map( D => n5398, CK => CLK, Q => OUT2(12), QN
                           => n4310);
   REGISTERS_reg_63_11_inst : DFF_X1 port map( D => n5397, CK => CLK, Q => 
                           n10098, QN => n4309);
   OUT2_reg_11_inst : DFF_X1 port map( D => n5396, CK => CLK, Q => OUT2(11), QN
                           => n4308);
   REGISTERS_reg_63_10_inst : DFF_X1 port map( D => n5395, CK => CLK, Q => 
                           n10099, QN => n4307);
   OUT2_reg_10_inst : DFF_X1 port map( D => n5394, CK => CLK, Q => OUT2(10), QN
                           => n4306);
   REGISTERS_reg_63_9_inst : DFF_X1 port map( D => n5393, CK => CLK, Q => 
                           n10100, QN => n4305);
   OUT2_reg_9_inst : DFF_X1 port map( D => n5392, CK => CLK, Q => OUT2(9), QN 
                           => n4304);
   REGISTERS_reg_63_8_inst : DFF_X1 port map( D => n5391, CK => CLK, Q => 
                           n10101, QN => n4303);
   OUT2_reg_8_inst : DFF_X1 port map( D => n5390, CK => CLK, Q => OUT2(8), QN 
                           => n4302);
   REGISTERS_reg_63_7_inst : DFF_X1 port map( D => n5389, CK => CLK, Q => 
                           n10102, QN => n4301);
   OUT2_reg_7_inst : DFF_X1 port map( D => n5388, CK => CLK, Q => OUT2(7), QN 
                           => n4300);
   REGISTERS_reg_63_6_inst : DFF_X1 port map( D => n5387, CK => CLK, Q => 
                           n10103, QN => n4299);
   OUT2_reg_6_inst : DFF_X1 port map( D => n5386, CK => CLK, Q => OUT2(6), QN 
                           => n4298);
   REGISTERS_reg_63_5_inst : DFF_X1 port map( D => n5385, CK => CLK, Q => 
                           n10104, QN => n4297);
   OUT2_reg_5_inst : DFF_X1 port map( D => n5384, CK => CLK, Q => OUT2(5), QN 
                           => n4296);
   REGISTERS_reg_63_4_inst : DFF_X1 port map( D => n5383, CK => CLK, Q => 
                           n10105, QN => n4295);
   OUT2_reg_4_inst : DFF_X1 port map( D => n5382, CK => CLK, Q => OUT2(4), QN 
                           => n4294);
   REGISTERS_reg_63_3_inst : DFF_X1 port map( D => n5381, CK => CLK, Q => 
                           n10106, QN => n4293);
   OUT2_reg_3_inst : DFF_X1 port map( D => n5380, CK => CLK, Q => OUT2(3), QN 
                           => n4292);
   REGISTERS_reg_63_2_inst : DFF_X1 port map( D => n5379, CK => CLK, Q => 
                           n10107, QN => n4291);
   OUT2_reg_2_inst : DFF_X1 port map( D => n5378, CK => CLK, Q => OUT2(2), QN 
                           => n4290);
   REGISTERS_reg_63_1_inst : DFF_X1 port map( D => n5377, CK => CLK, Q => 
                           n10108, QN => n4289);
   OUT2_reg_1_inst : DFF_X1 port map( D => n5376, CK => CLK, Q => OUT2(1), QN 
                           => n4288);
   REGISTERS_reg_63_0_inst : DFF_X1 port map( D => n5375, CK => CLK, Q => 
                           n10109, QN => n4287);
   OUT2_reg_0_inst : DFF_X1 port map( D => n5374, CK => CLK, Q => OUT2(0), QN 
                           => n4286);
   OUT1_reg_31_inst : DFF_X1 port map( D => n5373, CK => CLK, Q => OUT1(31), QN
                           => n4285);
   OUT1_reg_30_inst : DFF_X1 port map( D => n5372, CK => CLK, Q => OUT1(30), QN
                           => n4284);
   OUT1_reg_29_inst : DFF_X1 port map( D => n5371, CK => CLK, Q => OUT1(29), QN
                           => n4283);
   OUT1_reg_28_inst : DFF_X1 port map( D => n5370, CK => CLK, Q => OUT1(28), QN
                           => n4282);
   OUT1_reg_27_inst : DFF_X1 port map( D => n5369, CK => CLK, Q => OUT1(27), QN
                           => n4281);
   OUT1_reg_26_inst : DFF_X1 port map( D => n5368, CK => CLK, Q => OUT1(26), QN
                           => n4280);
   OUT1_reg_25_inst : DFF_X1 port map( D => n5367, CK => CLK, Q => OUT1(25), QN
                           => n4279);
   OUT1_reg_24_inst : DFF_X1 port map( D => n5366, CK => CLK, Q => OUT1(24), QN
                           => n4278);
   OUT1_reg_23_inst : DFF_X1 port map( D => n5365, CK => CLK, Q => OUT1(23), QN
                           => n4277);
   OUT1_reg_22_inst : DFF_X1 port map( D => n5364, CK => CLK, Q => OUT1(22), QN
                           => n4276);
   OUT1_reg_21_inst : DFF_X1 port map( D => n5363, CK => CLK, Q => OUT1(21), QN
                           => n4275);
   OUT1_reg_20_inst : DFF_X1 port map( D => n5362, CK => CLK, Q => OUT1(20), QN
                           => n4274);
   OUT1_reg_19_inst : DFF_X1 port map( D => n5361, CK => CLK, Q => OUT1(19), QN
                           => n4273);
   OUT1_reg_18_inst : DFF_X1 port map( D => n5360, CK => CLK, Q => OUT1(18), QN
                           => n4272);
   OUT1_reg_17_inst : DFF_X1 port map( D => n5359, CK => CLK, Q => OUT1(17), QN
                           => n4271);
   OUT1_reg_16_inst : DFF_X1 port map( D => n5358, CK => CLK, Q => OUT1(16), QN
                           => n4270);
   OUT1_reg_15_inst : DFF_X1 port map( D => n5357, CK => CLK, Q => OUT1(15), QN
                           => n4269);
   OUT1_reg_14_inst : DFF_X1 port map( D => n5356, CK => CLK, Q => OUT1(14), QN
                           => n4268);
   OUT1_reg_13_inst : DFF_X1 port map( D => n5355, CK => CLK, Q => OUT1(13), QN
                           => n4267);
   OUT1_reg_12_inst : DFF_X1 port map( D => n5354, CK => CLK, Q => OUT1(12), QN
                           => n4266);
   OUT1_reg_11_inst : DFF_X1 port map( D => n5353, CK => CLK, Q => OUT1(11), QN
                           => n4265);
   OUT1_reg_10_inst : DFF_X1 port map( D => n5352, CK => CLK, Q => OUT1(10), QN
                           => n4264);
   OUT1_reg_9_inst : DFF_X1 port map( D => n5351, CK => CLK, Q => OUT1(9), QN 
                           => n4263);
   OUT1_reg_8_inst : DFF_X1 port map( D => n5350, CK => CLK, Q => OUT1(8), QN 
                           => n4262);
   OUT1_reg_7_inst : DFF_X1 port map( D => n5349, CK => CLK, Q => OUT1(7), QN 
                           => n4261);
   OUT1_reg_6_inst : DFF_X1 port map( D => n5348, CK => CLK, Q => OUT1(6), QN 
                           => n4260);
   OUT1_reg_5_inst : DFF_X1 port map( D => n5347, CK => CLK, Q => OUT1(5), QN 
                           => n4259);
   OUT1_reg_4_inst : DFF_X1 port map( D => n5346, CK => CLK, Q => OUT1(4), QN 
                           => n4258);
   OUT1_reg_3_inst : DFF_X1 port map( D => n5345, CK => CLK, Q => OUT1(3), QN 
                           => n4257);
   OUT1_reg_2_inst : DFF_X1 port map( D => n5344, CK => CLK, Q => OUT1(2), QN 
                           => n4256);
   OUT1_reg_1_inst : DFF_X1 port map( D => n5343, CK => CLK, Q => OUT1(1), QN 
                           => n4255);
   OUT1_reg_0_inst : DFF_X1 port map( D => n5342, CK => CLK, Q => OUT1(0), QN 
                           => n4254);
   U10604 : NOR2_X2 port map( A1 => n18374, A2 => n18375, ZN => n18350);
   U13037 : NOR2_X2 port map( A1 => n19645, A2 => n19646, ZN => n19623);
   U13040 : NAND3_X1 port map( A1 => ENABLE, A2 => n22380, A3 => RD2, ZN => 
                           n18343);
   U13041 : NAND3_X1 port map( A1 => ENABLE, A2 => n22380, A3 => RD1, ZN => 
                           n19616);
   REGISTERS_reg_60_31_inst : DFF_X1 port map( D => n5533, CK => CLK, Q => 
                           n9026, QN => n16761);
   REGISTERS_reg_60_30_inst : DFF_X1 port map( D => n5532, CK => CLK, Q => 
                           n9037, QN => n16762);
   REGISTERS_reg_60_29_inst : DFF_X1 port map( D => n5531, CK => CLK, Q => 
                           n9048, QN => n16763);
   REGISTERS_reg_60_28_inst : DFF_X1 port map( D => n5530, CK => CLK, Q => 
                           n9059, QN => n16764);
   REGISTERS_reg_60_27_inst : DFF_X1 port map( D => n5529, CK => CLK, Q => 
                           n9070, QN => n16765);
   REGISTERS_reg_60_26_inst : DFF_X1 port map( D => n5528, CK => CLK, Q => 
                           n9081, QN => n16766);
   REGISTERS_reg_60_25_inst : DFF_X1 port map( D => n5527, CK => CLK, Q => 
                           n9092, QN => n16767);
   REGISTERS_reg_60_24_inst : DFF_X1 port map( D => n5526, CK => CLK, Q => 
                           n9103, QN => n16768);
   REGISTERS_reg_61_31_inst : DFF_X1 port map( D => n5501, CK => CLK, Q => 
                           n9030, QN => n16798);
   REGISTERS_reg_61_30_inst : DFF_X1 port map( D => n5500, CK => CLK, Q => 
                           n9041, QN => n16799);
   REGISTERS_reg_61_29_inst : DFF_X1 port map( D => n5499, CK => CLK, Q => 
                           n9052, QN => n16800);
   REGISTERS_reg_61_28_inst : DFF_X1 port map( D => n5498, CK => CLK, Q => 
                           n9063, QN => n16801);
   REGISTERS_reg_61_27_inst : DFF_X1 port map( D => n5497, CK => CLK, Q => 
                           n9074, QN => n16802);
   REGISTERS_reg_61_26_inst : DFF_X1 port map( D => n5496, CK => CLK, Q => 
                           n9085, QN => n16803);
   REGISTERS_reg_61_25_inst : DFF_X1 port map( D => n5495, CK => CLK, Q => 
                           n9096, QN => n16804);
   REGISTERS_reg_61_24_inst : DFF_X1 port map( D => n5494, CK => CLK, Q => 
                           n9107, QN => n16805);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n7389, CK => CLK, Q => n8958
                           , QN => n15159);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n7388, CK => CLK, Q => n8960
                           , QN => n15160);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n7387, CK => CLK, Q => n8962
                           , QN => n15161);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n7386, CK => CLK, Q => n8964
                           , QN => n15162);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n7385, CK => CLK, Q => n8966
                           , QN => n15163);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n7384, CK => CLK, Q => n8968
                           , QN => n15164);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n7383, CK => CLK, Q => n8970
                           , QN => n15165);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n7382, CK => CLK, Q => n8972
                           , QN => n15166);
   REGISTERS_reg_56_31_inst : DFF_X1 port map( D => n5661, CK => CLK, Q => 
                           n8578, QN => n16656);
   REGISTERS_reg_56_30_inst : DFF_X1 port map( D => n5660, CK => CLK, Q => 
                           n8589, QN => n16657);
   REGISTERS_reg_56_29_inst : DFF_X1 port map( D => n5659, CK => CLK, Q => 
                           n8600, QN => n16658);
   REGISTERS_reg_56_28_inst : DFF_X1 port map( D => n5658, CK => CLK, Q => 
                           n8611, QN => n16659);
   REGISTERS_reg_56_27_inst : DFF_X1 port map( D => n5657, CK => CLK, Q => 
                           n8622, QN => n16660);
   REGISTERS_reg_56_26_inst : DFF_X1 port map( D => n5656, CK => CLK, Q => 
                           n8633, QN => n16661);
   REGISTERS_reg_56_25_inst : DFF_X1 port map( D => n5655, CK => CLK, Q => 
                           n8644, QN => n16662);
   REGISTERS_reg_56_24_inst : DFF_X1 port map( D => n5654, CK => CLK, Q => 
                           n8655, QN => n16663);
   REGISTERS_reg_58_31_inst : DFF_X1 port map( D => n5597, CK => CLK, Q => 
                           n20686, QN => n16725);
   REGISTERS_reg_58_30_inst : DFF_X1 port map( D => n5596, CK => CLK, Q => 
                           n20685, QN => n16726);
   REGISTERS_reg_58_29_inst : DFF_X1 port map( D => n5595, CK => CLK, Q => 
                           n20684, QN => n16727);
   REGISTERS_reg_58_28_inst : DFF_X1 port map( D => n5594, CK => CLK, Q => 
                           n20683, QN => n16728);
   REGISTERS_reg_58_27_inst : DFF_X1 port map( D => n5593, CK => CLK, Q => 
                           n20682, QN => n16729);
   REGISTERS_reg_58_26_inst : DFF_X1 port map( D => n5592, CK => CLK, Q => 
                           n20681, QN => n16730);
   REGISTERS_reg_58_25_inst : DFF_X1 port map( D => n5591, CK => CLK, Q => 
                           n20680, QN => n16731);
   REGISTERS_reg_58_24_inst : DFF_X1 port map( D => n5590, CK => CLK, Q => 
                           n20679, QN => n16732);
   REGISTERS_reg_55_31_inst : DFF_X1 port map( D => n5693, CK => CLK, Q => 
                           n8576, QN => n16621);
   REGISTERS_reg_55_30_inst : DFF_X1 port map( D => n5692, CK => CLK, Q => 
                           n8587, QN => n16622);
   REGISTERS_reg_55_29_inst : DFF_X1 port map( D => n5691, CK => CLK, Q => 
                           n8598, QN => n16623);
   REGISTERS_reg_55_28_inst : DFF_X1 port map( D => n5690, CK => CLK, Q => 
                           n8609, QN => n16624);
   REGISTERS_reg_55_27_inst : DFF_X1 port map( D => n5689, CK => CLK, Q => 
                           n8620, QN => n16625);
   REGISTERS_reg_55_26_inst : DFF_X1 port map( D => n5688, CK => CLK, Q => 
                           n8631, QN => n16626);
   REGISTERS_reg_55_25_inst : DFF_X1 port map( D => n5687, CK => CLK, Q => 
                           n8642, QN => n16627);
   REGISTERS_reg_55_24_inst : DFF_X1 port map( D => n5686, CK => CLK, Q => 
                           n8653, QN => n16628);
   REGISTERS_reg_47_31_inst : DFF_X1 port map( D => n5949, CK => CLK, Q => 
                           n20678, QN => n16488);
   REGISTERS_reg_47_30_inst : DFF_X1 port map( D => n5948, CK => CLK, Q => 
                           n20677, QN => n16489);
   REGISTERS_reg_47_29_inst : DFF_X1 port map( D => n5947, CK => CLK, Q => 
                           n20676, QN => n16490);
   REGISTERS_reg_47_28_inst : DFF_X1 port map( D => n5946, CK => CLK, Q => 
                           n20675, QN => n16491);
   REGISTERS_reg_47_27_inst : DFF_X1 port map( D => n5945, CK => CLK, Q => 
                           n20674, QN => n16492);
   REGISTERS_reg_47_26_inst : DFF_X1 port map( D => n5944, CK => CLK, Q => 
                           n20673, QN => n16493);
   REGISTERS_reg_47_25_inst : DFF_X1 port map( D => n5943, CK => CLK, Q => 
                           n20672, QN => n16494);
   REGISTERS_reg_47_24_inst : DFF_X1 port map( D => n5942, CK => CLK, Q => 
                           n20671, QN => n16495);
   REGISTERS_reg_43_31_inst : DFF_X1 port map( D => n6077, CK => CLK, Q => 
                           n20670, QN => n16351);
   REGISTERS_reg_43_30_inst : DFF_X1 port map( D => n6076, CK => CLK, Q => 
                           n20669, QN => n16352);
   REGISTERS_reg_43_29_inst : DFF_X1 port map( D => n6075, CK => CLK, Q => 
                           n20668, QN => n16353);
   REGISTERS_reg_43_28_inst : DFF_X1 port map( D => n6074, CK => CLK, Q => 
                           n20667, QN => n16354);
   REGISTERS_reg_43_27_inst : DFF_X1 port map( D => n6073, CK => CLK, Q => 
                           n20666, QN => n16355);
   REGISTERS_reg_43_26_inst : DFF_X1 port map( D => n6072, CK => CLK, Q => 
                           n20665, QN => n16356);
   REGISTERS_reg_43_25_inst : DFF_X1 port map( D => n6071, CK => CLK, Q => 
                           n20664, QN => n16357);
   REGISTERS_reg_43_24_inst : DFF_X1 port map( D => n6070, CK => CLK, Q => 
                           n20663, QN => n16358);
   REGISTERS_reg_57_31_inst : DFF_X1 port map( D => n5629, CK => CLK, Q => 
                           n8582, QN => n16691);
   REGISTERS_reg_57_30_inst : DFF_X1 port map( D => n5628, CK => CLK, Q => 
                           n8593, QN => n16692);
   REGISTERS_reg_57_29_inst : DFF_X1 port map( D => n5627, CK => CLK, Q => 
                           n8604, QN => n16693);
   REGISTERS_reg_57_28_inst : DFF_X1 port map( D => n5626, CK => CLK, Q => 
                           n8615, QN => n16694);
   REGISTERS_reg_57_27_inst : DFF_X1 port map( D => n5625, CK => CLK, Q => 
                           n8626, QN => n16695);
   REGISTERS_reg_57_26_inst : DFF_X1 port map( D => n5624, CK => CLK, Q => 
                           n8637, QN => n16696);
   REGISTERS_reg_57_25_inst : DFF_X1 port map( D => n5623, CK => CLK, Q => 
                           n8648, QN => n16697);
   REGISTERS_reg_57_24_inst : DFF_X1 port map( D => n5622, CK => CLK, Q => 
                           n8659, QN => n16698);
   REGISTERS_reg_50_31_inst : DFF_X1 port map( D => n5853, CK => CLK, Q => 
                           n8478, QN => n16577);
   REGISTERS_reg_50_30_inst : DFF_X1 port map( D => n5852, CK => CLK, Q => 
                           n8479, QN => n16578);
   REGISTERS_reg_50_29_inst : DFF_X1 port map( D => n5851, CK => CLK, Q => 
                           n8480, QN => n16579);
   REGISTERS_reg_50_28_inst : DFF_X1 port map( D => n5850, CK => CLK, Q => 
                           n8481, QN => n16580);
   REGISTERS_reg_50_27_inst : DFF_X1 port map( D => n5849, CK => CLK, Q => 
                           n8482, QN => n16581);
   REGISTERS_reg_50_26_inst : DFF_X1 port map( D => n5848, CK => CLK, Q => 
                           n8483, QN => n16582);
   REGISTERS_reg_50_25_inst : DFF_X1 port map( D => n5847, CK => CLK, Q => 
                           n8484, QN => n16583);
   REGISTERS_reg_50_24_inst : DFF_X1 port map( D => n5846, CK => CLK, Q => 
                           n8485, QN => n16584);
   REGISTERS_reg_49_31_inst : DFF_X1 port map( D => n5885, CK => CLK, Q => 
                           n20662, QN => n16557);
   REGISTERS_reg_49_30_inst : DFF_X1 port map( D => n5884, CK => CLK, Q => 
                           n20661, QN => n16558);
   REGISTERS_reg_49_29_inst : DFF_X1 port map( D => n5883, CK => CLK, Q => 
                           n20660, QN => n16559);
   REGISTERS_reg_49_28_inst : DFF_X1 port map( D => n5882, CK => CLK, Q => 
                           n20659, QN => n16560);
   REGISTERS_reg_49_27_inst : DFF_X1 port map( D => n5881, CK => CLK, Q => 
                           n20658, QN => n16561);
   REGISTERS_reg_49_26_inst : DFF_X1 port map( D => n5880, CK => CLK, Q => 
                           n20657, QN => n16562);
   REGISTERS_reg_49_25_inst : DFF_X1 port map( D => n5879, CK => CLK, Q => 
                           n20656, QN => n16563);
   REGISTERS_reg_49_24_inst : DFF_X1 port map( D => n5878, CK => CLK, Q => 
                           n20655, QN => n16564);
   REGISTERS_reg_48_31_inst : DFF_X1 port map( D => n5917, CK => CLK, Q => 
                           n20654, QN => n16522);
   REGISTERS_reg_48_30_inst : DFF_X1 port map( D => n5916, CK => CLK, Q => 
                           n20653, QN => n16523);
   REGISTERS_reg_48_29_inst : DFF_X1 port map( D => n5915, CK => CLK, Q => 
                           n20652, QN => n16524);
   REGISTERS_reg_48_28_inst : DFF_X1 port map( D => n5914, CK => CLK, Q => 
                           n20651, QN => n16525);
   REGISTERS_reg_48_27_inst : DFF_X1 port map( D => n5913, CK => CLK, Q => 
                           n20650, QN => n16526);
   REGISTERS_reg_48_26_inst : DFF_X1 port map( D => n5912, CK => CLK, Q => 
                           n20649, QN => n16527);
   REGISTERS_reg_48_25_inst : DFF_X1 port map( D => n5911, CK => CLK, Q => 
                           n20648, QN => n16528);
   REGISTERS_reg_48_24_inst : DFF_X1 port map( D => n5910, CK => CLK, Q => 
                           n20647, QN => n16529);
   REGISTERS_reg_46_31_inst : DFF_X1 port map( D => n5981, CK => CLK, Q => 
                           n8574, QN => n16454);
   REGISTERS_reg_46_30_inst : DFF_X1 port map( D => n5980, CK => CLK, Q => 
                           n8585, QN => n16455);
   REGISTERS_reg_46_29_inst : DFF_X1 port map( D => n5979, CK => CLK, Q => 
                           n8596, QN => n16456);
   REGISTERS_reg_46_28_inst : DFF_X1 port map( D => n5978, CK => CLK, Q => 
                           n8607, QN => n16457);
   REGISTERS_reg_46_27_inst : DFF_X1 port map( D => n5977, CK => CLK, Q => 
                           n8618, QN => n16458);
   REGISTERS_reg_46_26_inst : DFF_X1 port map( D => n5976, CK => CLK, Q => 
                           n8629, QN => n16459);
   REGISTERS_reg_46_25_inst : DFF_X1 port map( D => n5975, CK => CLK, Q => 
                           n8640, QN => n16460);
   REGISTERS_reg_46_24_inst : DFF_X1 port map( D => n5974, CK => CLK, Q => 
                           n8651, QN => n16461);
   REGISTERS_reg_44_31_inst : DFF_X1 port map( D => n6045, CK => CLK, Q => 
                           n9886, QN => n16385);
   REGISTERS_reg_44_30_inst : DFF_X1 port map( D => n6044, CK => CLK, Q => 
                           n9887, QN => n16386);
   REGISTERS_reg_44_29_inst : DFF_X1 port map( D => n6043, CK => CLK, Q => 
                           n9888, QN => n16387);
   REGISTERS_reg_44_28_inst : DFF_X1 port map( D => n6042, CK => CLK, Q => 
                           n9889, QN => n16388);
   REGISTERS_reg_44_27_inst : DFF_X1 port map( D => n6041, CK => CLK, Q => 
                           n9890, QN => n16389);
   REGISTERS_reg_44_26_inst : DFF_X1 port map( D => n6040, CK => CLK, Q => 
                           n9891, QN => n16390);
   REGISTERS_reg_44_25_inst : DFF_X1 port map( D => n6039, CK => CLK, Q => 
                           n9892, QN => n16391);
   REGISTERS_reg_44_24_inst : DFF_X1 port map( D => n6038, CK => CLK, Q => 
                           n9893, QN => n16392);
   REGISTERS_reg_39_31_inst : DFF_X1 port map( D => n6205, CK => CLK, Q => 
                           n20646, QN => n16310);
   REGISTERS_reg_39_30_inst : DFF_X1 port map( D => n6204, CK => CLK, Q => 
                           n20645, QN => n16311);
   REGISTERS_reg_39_29_inst : DFF_X1 port map( D => n6203, CK => CLK, Q => 
                           n20644, QN => n16312);
   REGISTERS_reg_39_28_inst : DFF_X1 port map( D => n6202, CK => CLK, Q => 
                           n20643, QN => n16313);
   REGISTERS_reg_39_27_inst : DFF_X1 port map( D => n6201, CK => CLK, Q => 
                           n20642, QN => n16314);
   REGISTERS_reg_39_26_inst : DFF_X1 port map( D => n6200, CK => CLK, Q => 
                           n20641, QN => n16315);
   REGISTERS_reg_39_25_inst : DFF_X1 port map( D => n6199, CK => CLK, Q => 
                           n20640, QN => n16316);
   REGISTERS_reg_39_24_inst : DFF_X1 port map( D => n6198, CK => CLK, Q => 
                           n20639, QN => n16317);
   REGISTERS_reg_35_31_inst : DFF_X1 port map( D => n6333, CK => CLK, Q => 
                           n20638, QN => n16172);
   REGISTERS_reg_35_30_inst : DFF_X1 port map( D => n6332, CK => CLK, Q => 
                           n20637, QN => n16173);
   REGISTERS_reg_35_29_inst : DFF_X1 port map( D => n6331, CK => CLK, Q => 
                           n20636, QN => n16174);
   REGISTERS_reg_35_28_inst : DFF_X1 port map( D => n6330, CK => CLK, Q => 
                           n20635, QN => n16175);
   REGISTERS_reg_35_27_inst : DFF_X1 port map( D => n6329, CK => CLK, Q => 
                           n20634, QN => n16176);
   REGISTERS_reg_35_26_inst : DFF_X1 port map( D => n6328, CK => CLK, Q => 
                           n20633, QN => n16177);
   REGISTERS_reg_35_25_inst : DFF_X1 port map( D => n6327, CK => CLK, Q => 
                           n20632, QN => n16178);
   REGISTERS_reg_35_24_inst : DFF_X1 port map( D => n6326, CK => CLK, Q => 
                           n20631, QN => n16179);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n6461, CK => CLK, Q => 
                           n20630, QN => n16067);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n6460, CK => CLK, Q => 
                           n20629, QN => n16068);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n6459, CK => CLK, Q => 
                           n20628, QN => n16069);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n6458, CK => CLK, Q => 
                           n20627, QN => n16070);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n6457, CK => CLK, Q => 
                           n20626, QN => n16071);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n6456, CK => CLK, Q => 
                           n20625, QN => n16072);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n6455, CK => CLK, Q => 
                           n20624, QN => n16073);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n6454, CK => CLK, Q => 
                           n20623, QN => n16074);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n6589, CK => CLK, Q => 
                           n9502, QN => n15930);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n6588, CK => CLK, Q => 
                           n9503, QN => n15931);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n6587, CK => CLK, Q => 
                           n9504, QN => n15932);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n6586, CK => CLK, Q => 
                           n9505, QN => n15933);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n6585, CK => CLK, Q => 
                           n9506, QN => n15934);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n6584, CK => CLK, Q => 
                           n9507, QN => n15935);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n6583, CK => CLK, Q => 
                           n9508, QN => n15936);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n6582, CK => CLK, Q => 
                           n9509, QN => n15937);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n6717, CK => CLK, Q => 
                           n9598, QN => n15857);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n6716, CK => CLK, Q => 
                           n9599, QN => n15858);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n6715, CK => CLK, Q => 
                           n9600, QN => n15859);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n6714, CK => CLK, Q => 
                           n9601, QN => n15860);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n6713, CK => CLK, Q => 
                           n9602, QN => n15861);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n6712, CK => CLK, Q => 
                           n9603, QN => n15862);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n6711, CK => CLK, Q => 
                           n9604, QN => n15863);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n6710, CK => CLK, Q => 
                           n9605, QN => n15864);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n6973, CK => CLK, Q => 
                           n8926, QN => n15610);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n6972, CK => CLK, Q => 
                           n8927, QN => n15611);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n6971, CK => CLK, Q => 
                           n8928, QN => n15612);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n6970, CK => CLK, Q => 
                           n8929, QN => n15613);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n6969, CK => CLK, Q => 
                           n8930, QN => n15614);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n6968, CK => CLK, Q => 
                           n8931, QN => n15615);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n6967, CK => CLK, Q => 
                           n8932, QN => n15616);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n6966, CK => CLK, Q => 
                           n8933, QN => n15617);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n7101, CK => CLK, Q => 
                           n20622, QN => n15472);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n7100, CK => CLK, Q => 
                           n20621, QN => n15473);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n7099, CK => CLK, Q => 
                           n20620, QN => n15474);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n7098, CK => CLK, Q => 
                           n20619, QN => n15475);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n7097, CK => CLK, Q => 
                           n20618, QN => n15476);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n7096, CK => CLK, Q => 
                           n20617, QN => n15477);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n7095, CK => CLK, Q => 
                           n20616, QN => n15478);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n7094, CK => CLK, Q => 
                           n20615, QN => n15479);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n7229, CK => CLK, Q => n8959
                           , QN => n15334);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n7228, CK => CLK, Q => n8961
                           , QN => n15335);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n7227, CK => CLK, Q => n8963
                           , QN => n15336);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n7226, CK => CLK, Q => n8965
                           , QN => n15337);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n7225, CK => CLK, Q => n8967
                           , QN => n15338);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n7224, CK => CLK, Q => n8969
                           , QN => n15339);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n7223, CK => CLK, Q => n8971
                           , QN => n15340);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n7222, CK => CLK, Q => n8973
                           , QN => n15341);
   REGISTERS_reg_45_31_inst : DFF_X1 port map( D => n6013, CK => CLK, Q => 
                           n9918, QN => n16420);
   REGISTERS_reg_45_30_inst : DFF_X1 port map( D => n6012, CK => CLK, Q => 
                           n9919, QN => n16421);
   REGISTERS_reg_45_29_inst : DFF_X1 port map( D => n6011, CK => CLK, Q => 
                           n9920, QN => n16422);
   REGISTERS_reg_45_28_inst : DFF_X1 port map( D => n6010, CK => CLK, Q => 
                           n9921, QN => n16423);
   REGISTERS_reg_45_27_inst : DFF_X1 port map( D => n6009, CK => CLK, Q => 
                           n9922, QN => n16424);
   REGISTERS_reg_45_26_inst : DFF_X1 port map( D => n6008, CK => CLK, Q => 
                           n9923, QN => n16425);
   REGISTERS_reg_45_25_inst : DFF_X1 port map( D => n6007, CK => CLK, Q => 
                           n9924, QN => n16426);
   REGISTERS_reg_45_24_inst : DFF_X1 port map( D => n6006, CK => CLK, Q => 
                           n9925, QN => n16427);
   REGISTERS_reg_38_31_inst : DFF_X1 port map( D => n6237, CK => CLK, Q => 
                           n8575, QN => n16276);
   REGISTERS_reg_38_30_inst : DFF_X1 port map( D => n6236, CK => CLK, Q => 
                           n8586, QN => n16277);
   REGISTERS_reg_38_29_inst : DFF_X1 port map( D => n6235, CK => CLK, Q => 
                           n8597, QN => n16278);
   REGISTERS_reg_38_28_inst : DFF_X1 port map( D => n6234, CK => CLK, Q => 
                           n8608, QN => n16279);
   REGISTERS_reg_38_27_inst : DFF_X1 port map( D => n6233, CK => CLK, Q => 
                           n8619, QN => n16280);
   REGISTERS_reg_38_26_inst : DFF_X1 port map( D => n6232, CK => CLK, Q => 
                           n8630, QN => n16281);
   REGISTERS_reg_38_25_inst : DFF_X1 port map( D => n6231, CK => CLK, Q => 
                           n8641, QN => n16282);
   REGISTERS_reg_38_24_inst : DFF_X1 port map( D => n6230, CK => CLK, Q => 
                           n8652, QN => n16283);
   REGISTERS_reg_37_31_inst : DFF_X1 port map( D => n6269, CK => CLK, Q => 
                           n20614, QN => n16242);
   REGISTERS_reg_37_30_inst : DFF_X1 port map( D => n6268, CK => CLK, Q => 
                           n20613, QN => n16243);
   REGISTERS_reg_37_29_inst : DFF_X1 port map( D => n6267, CK => CLK, Q => 
                           n20612, QN => n16244);
   REGISTERS_reg_37_28_inst : DFF_X1 port map( D => n6266, CK => CLK, Q => 
                           n20611, QN => n16245);
   REGISTERS_reg_37_27_inst : DFF_X1 port map( D => n6265, CK => CLK, Q => 
                           n20610, QN => n16246);
   REGISTERS_reg_37_26_inst : DFF_X1 port map( D => n6264, CK => CLK, Q => 
                           n20609, QN => n16247);
   REGISTERS_reg_37_25_inst : DFF_X1 port map( D => n6263, CK => CLK, Q => 
                           n20608, QN => n16248);
   REGISTERS_reg_37_24_inst : DFF_X1 port map( D => n6262, CK => CLK, Q => 
                           n20607, QN => n16249);
   REGISTERS_reg_36_31_inst : DFF_X1 port map( D => n6301, CK => CLK, Q => 
                           n20606, QN => n16207);
   REGISTERS_reg_36_30_inst : DFF_X1 port map( D => n6300, CK => CLK, Q => 
                           n20605, QN => n16208);
   REGISTERS_reg_36_29_inst : DFF_X1 port map( D => n6299, CK => CLK, Q => 
                           n20604, QN => n16209);
   REGISTERS_reg_36_28_inst : DFF_X1 port map( D => n6298, CK => CLK, Q => 
                           n20603, QN => n16210);
   REGISTERS_reg_36_27_inst : DFF_X1 port map( D => n6297, CK => CLK, Q => 
                           n20602, QN => n16211);
   REGISTERS_reg_36_26_inst : DFF_X1 port map( D => n6296, CK => CLK, Q => 
                           n20601, QN => n16212);
   REGISTERS_reg_36_25_inst : DFF_X1 port map( D => n6295, CK => CLK, Q => 
                           n20600, QN => n16213);
   REGISTERS_reg_36_24_inst : DFF_X1 port map( D => n6294, CK => CLK, Q => 
                           n20599, QN => n16214);
   REGISTERS_reg_33_31_inst : DFF_X1 port map( D => n6397, CK => CLK, Q => 
                           n20598, QN => n16136);
   REGISTERS_reg_33_30_inst : DFF_X1 port map( D => n6396, CK => CLK, Q => 
                           n20597, QN => n16137);
   REGISTERS_reg_33_29_inst : DFF_X1 port map( D => n6395, CK => CLK, Q => 
                           n20596, QN => n16138);
   REGISTERS_reg_33_28_inst : DFF_X1 port map( D => n6394, CK => CLK, Q => 
                           n20595, QN => n16139);
   REGISTERS_reg_33_27_inst : DFF_X1 port map( D => n6393, CK => CLK, Q => 
                           n20594, QN => n16140);
   REGISTERS_reg_33_26_inst : DFF_X1 port map( D => n6392, CK => CLK, Q => 
                           n20593, QN => n16141);
   REGISTERS_reg_33_25_inst : DFF_X1 port map( D => n6391, CK => CLK, Q => 
                           n20592, QN => n16142);
   REGISTERS_reg_33_24_inst : DFF_X1 port map( D => n6390, CK => CLK, Q => 
                           n20591, QN => n16143);
   REGISTERS_reg_32_31_inst : DFF_X1 port map( D => n6429, CK => CLK, Q => 
                           n20590, QN => n16101);
   REGISTERS_reg_32_30_inst : DFF_X1 port map( D => n6428, CK => CLK, Q => 
                           n20589, QN => n16102);
   REGISTERS_reg_32_29_inst : DFF_X1 port map( D => n6427, CK => CLK, Q => 
                           n20588, QN => n16103);
   REGISTERS_reg_32_28_inst : DFF_X1 port map( D => n6426, CK => CLK, Q => 
                           n20587, QN => n16104);
   REGISTERS_reg_32_27_inst : DFF_X1 port map( D => n6425, CK => CLK, Q => 
                           n20586, QN => n16105);
   REGISTERS_reg_32_26_inst : DFF_X1 port map( D => n6424, CK => CLK, Q => 
                           n20585, QN => n16106);
   REGISTERS_reg_32_25_inst : DFF_X1 port map( D => n6423, CK => CLK, Q => 
                           n20584, QN => n16107);
   REGISTERS_reg_32_24_inst : DFF_X1 port map( D => n6422, CK => CLK, Q => 
                           n20583, QN => n16108);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n6493, CK => CLK, Q => 
                           n20582, QN => n16033);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n6492, CK => CLK, Q => 
                           n20581, QN => n16034);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n6491, CK => CLK, Q => 
                           n20580, QN => n16035);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n6490, CK => CLK, Q => 
                           n20579, QN => n16036);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n6489, CK => CLK, Q => 
                           n20578, QN => n16037);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n6488, CK => CLK, Q => 
                           n20577, QN => n16038);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n6487, CK => CLK, Q => 
                           n20576, QN => n16039);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n6486, CK => CLK, Q => 
                           n20575, QN => n16040);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n6525, CK => CLK, Q => 
                           n9822, QN => n15999);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n6524, CK => CLK, Q => 
                           n9823, QN => n16000);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n6523, CK => CLK, Q => 
                           n9824, QN => n16001);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n6522, CK => CLK, Q => 
                           n9825, QN => n16002);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n6521, CK => CLK, Q => 
                           n9826, QN => n16003);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n6520, CK => CLK, Q => 
                           n9827, QN => n16004);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n6519, CK => CLK, Q => 
                           n9828, QN => n16005);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n6518, CK => CLK, Q => 
                           n9829, QN => n16006);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n6557, CK => CLK, Q => 
                           n9790, QN => n15964);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n6556, CK => CLK, Q => 
                           n9791, QN => n15965);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n6555, CK => CLK, Q => 
                           n9792, QN => n15966);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n6554, CK => CLK, Q => 
                           n9793, QN => n15967);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n6553, CK => CLK, Q => 
                           n9794, QN => n15968);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n6552, CK => CLK, Q => 
                           n9795, QN => n15969);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n6551, CK => CLK, Q => 
                           n9796, QN => n15970);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n6550, CK => CLK, Q => 
                           n9797, QN => n15971);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n6621, CK => CLK, Q => 
                           n20574, QN => n15896);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n6620, CK => CLK, Q => 
                           n20573, QN => n15897);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n6619, CK => CLK, Q => 
                           n20572, QN => n15898);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n6618, CK => CLK, Q => 
                           n20571, QN => n15899);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n6617, CK => CLK, Q => 
                           n20570, QN => n15900);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n6616, CK => CLK, Q => 
                           n20569, QN => n15901);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n6615, CK => CLK, Q => 
                           n20568, QN => n15902);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n6614, CK => CLK, Q => 
                           n20567, QN => n15903);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n6749, CK => CLK, Q => 
                           n20566, QN => n15823);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n6748, CK => CLK, Q => 
                           n20565, QN => n15824);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n6747, CK => CLK, Q => 
                           n20564, QN => n15825);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n6746, CK => CLK, Q => 
                           n20563, QN => n15826);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n6745, CK => CLK, Q => 
                           n20562, QN => n15827);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n6744, CK => CLK, Q => 
                           n20561, QN => n15828);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n6743, CK => CLK, Q => 
                           n20560, QN => n15829);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n6742, CK => CLK, Q => 
                           n20559, QN => n15830);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n6781, CK => CLK, Q => 
                           n20558, QN => n15789);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n6780, CK => CLK, Q => 
                           n20557, QN => n15790);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n6779, CK => CLK, Q => 
                           n20556, QN => n15791);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n6778, CK => CLK, Q => 
                           n20555, QN => n15792);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n6777, CK => CLK, Q => 
                           n20554, QN => n15793);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n6776, CK => CLK, Q => 
                           n20553, QN => n15794);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n6775, CK => CLK, Q => 
                           n20552, QN => n15795);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n6774, CK => CLK, Q => 
                           n20551, QN => n15796);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n6813, CK => CLK, Q => 
                           n20550, QN => n15754);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n6812, CK => CLK, Q => 
                           n20549, QN => n15755);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n6811, CK => CLK, Q => 
                           n20548, QN => n15756);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n6810, CK => CLK, Q => 
                           n20547, QN => n15757);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n6809, CK => CLK, Q => 
                           n20546, QN => n15758);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n6808, CK => CLK, Q => 
                           n20545, QN => n15759);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n6807, CK => CLK, Q => 
                           n20544, QN => n15760);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n6806, CK => CLK, Q => 
                           n20543, QN => n15761);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n6877, CK => CLK, Q => 
                           n9438, QN => n15717);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n6876, CK => CLK, Q => 
                           n9439, QN => n15718);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n6875, CK => CLK, Q => 
                           n9440, QN => n15719);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n6874, CK => CLK, Q => 
                           n9441, QN => n15720);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n6873, CK => CLK, Q => 
                           n9442, QN => n15721);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n6872, CK => CLK, Q => 
                           n9443, QN => n15722);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n6871, CK => CLK, Q => 
                           n9444, QN => n15723);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n6870, CK => CLK, Q => 
                           n9445, QN => n15724);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n6909, CK => CLK, Q => 
                           n20542, QN => n15683);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n6908, CK => CLK, Q => 
                           n20541, QN => n15684);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n6907, CK => CLK, Q => 
                           n20540, QN => n15685);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n6906, CK => CLK, Q => 
                           n20539, QN => n15686);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n6905, CK => CLK, Q => 
                           n20538, QN => n15687);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n6904, CK => CLK, Q => 
                           n20537, QN => n15688);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n6903, CK => CLK, Q => 
                           n20536, QN => n15689);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n6902, CK => CLK, Q => 
                           n20535, QN => n15690);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n6941, CK => CLK, Q => 
                           n20534, QN => n15648);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n6940, CK => CLK, Q => 
                           n20533, QN => n15649);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n6939, CK => CLK, Q => 
                           n20532, QN => n15650);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n6938, CK => CLK, Q => 
                           n20531, QN => n15651);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n6937, CK => CLK, Q => 
                           n20530, QN => n15652);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n6936, CK => CLK, Q => 
                           n20529, QN => n15653);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n6935, CK => CLK, Q => 
                           n20528, QN => n15654);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n6934, CK => CLK, Q => 
                           n20527, QN => n15655);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n7005, CK => CLK, Q => 
                           n20526, QN => n15576);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n7004, CK => CLK, Q => 
                           n20525, QN => n15577);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n7003, CK => CLK, Q => 
                           n20524, QN => n15578);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n7002, CK => CLK, Q => 
                           n20523, QN => n15579);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n7001, CK => CLK, Q => 
                           n20522, QN => n15580);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n7000, CK => CLK, Q => 
                           n20521, QN => n15581);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n6999, CK => CLK, Q => 
                           n20520, QN => n15582);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n6998, CK => CLK, Q => 
                           n20519, QN => n15583);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n7037, CK => CLK, Q => 
                           n8584, QN => n15542);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n7036, CK => CLK, Q => 
                           n8595, QN => n15543);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n7035, CK => CLK, Q => 
                           n8606, QN => n15544);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n7034, CK => CLK, Q => 
                           n8617, QN => n15545);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n7033, CK => CLK, Q => 
                           n8628, QN => n15546);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n7032, CK => CLK, Q => 
                           n8639, QN => n15547);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n7031, CK => CLK, Q => 
                           n8650, QN => n15548);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n7030, CK => CLK, Q => 
                           n8661, QN => n15549);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n7069, CK => CLK, Q => 
                           n8580, QN => n15507);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n7068, CK => CLK, Q => 
                           n8591, QN => n15508);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n7067, CK => CLK, Q => 
                           n8602, QN => n15509);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n7066, CK => CLK, Q => 
                           n8613, QN => n15510);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n7065, CK => CLK, Q => 
                           n8624, QN => n15511);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n7064, CK => CLK, Q => 
                           n8635, QN => n15512);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n7063, CK => CLK, Q => 
                           n8646, QN => n15513);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n7062, CK => CLK, Q => 
                           n8657, QN => n15514);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n7133, CK => CLK, Q => 
                           n20518, QN => n15438);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n7132, CK => CLK, Q => 
                           n20517, QN => n15439);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n7131, CK => CLK, Q => 
                           n20516, QN => n15440);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n7130, CK => CLK, Q => 
                           n20515, QN => n15441);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n7129, CK => CLK, Q => 
                           n20514, QN => n15442);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n7128, CK => CLK, Q => 
                           n20513, QN => n15443);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n7127, CK => CLK, Q => 
                           n20512, QN => n15444);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n7126, CK => CLK, Q => 
                           n20511, QN => n15445);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n7165, CK => CLK, Q => 
                           n20510, QN => n15404);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n7164, CK => CLK, Q => 
                           n20509, QN => n15405);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n7163, CK => CLK, Q => 
                           n20508, QN => n15406);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n7162, CK => CLK, Q => 
                           n20507, QN => n15407);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n7161, CK => CLK, Q => 
                           n20506, QN => n15408);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n7160, CK => CLK, Q => 
                           n20505, QN => n15409);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n7159, CK => CLK, Q => 
                           n20504, QN => n15410);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n7158, CK => CLK, Q => 
                           n20503, QN => n15411);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n7197, CK => CLK, Q => 
                           n20502, QN => n15369);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n7196, CK => CLK, Q => 
                           n20501, QN => n15370);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n7195, CK => CLK, Q => 
                           n20500, QN => n15371);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n7194, CK => CLK, Q => 
                           n20499, QN => n15372);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n7193, CK => CLK, Q => 
                           n20498, QN => n15373);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n7192, CK => CLK, Q => 
                           n20497, QN => n15374);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n7191, CK => CLK, Q => 
                           n20496, QN => n15375);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n7190, CK => CLK, Q => 
                           n20495, QN => n15376);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n7261, CK => CLK, Q => n8511
                           , QN => n15300);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n7260, CK => CLK, Q => n8513
                           , QN => n15301);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n7259, CK => CLK, Q => n8515
                           , QN => n15302);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n7258, CK => CLK, Q => n8517
                           , QN => n15303);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n7257, CK => CLK, Q => n8519
                           , QN => n15304);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n7256, CK => CLK, Q => n8521
                           , QN => n15305);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n7255, CK => CLK, Q => n8523
                           , QN => n15306);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n7254, CK => CLK, Q => n8525
                           , QN => n15307);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n7293, CK => CLK, Q => 
                           n20494, QN => n15266);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n7292, CK => CLK, Q => 
                           n20493, QN => n15267);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n7291, CK => CLK, Q => 
                           n20492, QN => n15268);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n7290, CK => CLK, Q => 
                           n20491, QN => n15269);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n7289, CK => CLK, Q => 
                           n20490, QN => n15270);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n7288, CK => CLK, Q => 
                           n20489, QN => n15271);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n7287, CK => CLK, Q => 
                           n20488, QN => n15272);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n7286, CK => CLK, Q => 
                           n20487, QN => n15273);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n7325, CK => CLK, Q => 
                           n20486, QN => n15231);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n7324, CK => CLK, Q => 
                           n20485, QN => n15232);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n7323, CK => CLK, Q => 
                           n20484, QN => n15233);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n7322, CK => CLK, Q => 
                           n20483, QN => n15234);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n7321, CK => CLK, Q => 
                           n20482, QN => n15235);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n7320, CK => CLK, Q => 
                           n20481, QN => n15236);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n7319, CK => CLK, Q => 
                           n20480, QN => n15237);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n7318, CK => CLK, Q => 
                           n20479, QN => n15238);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n7357, CK => CLK, Q => n8510
                           , QN => n15194);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n7356, CK => CLK, Q => n8512
                           , QN => n15195);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n7355, CK => CLK, Q => n8514
                           , QN => n15196);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n7354, CK => CLK, Q => n8516
                           , QN => n15197);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n7353, CK => CLK, Q => n8518
                           , QN => n15198);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n7352, CK => CLK, Q => n8520
                           , QN => n15199);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n7351, CK => CLK, Q => n8522
                           , QN => n15200);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n7350, CK => CLK, Q => n8524
                           , QN => n15201);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n7358, CK => CLK, Q => n9020,
                           QN => n15190);
   REGISTERS_reg_44_23_inst : DFF_X1 port map( D => n6037, CK => CLK, Q => 
                           n9894, QN => n16393);
   REGISTERS_reg_44_22_inst : DFF_X1 port map( D => n6036, CK => CLK, Q => 
                           n9895, QN => n16394);
   REGISTERS_reg_44_21_inst : DFF_X1 port map( D => n6035, CK => CLK, Q => 
                           n9896, QN => n16395);
   REGISTERS_reg_44_20_inst : DFF_X1 port map( D => n6034, CK => CLK, Q => 
                           n9897, QN => n16396);
   REGISTERS_reg_44_19_inst : DFF_X1 port map( D => n6033, CK => CLK, Q => 
                           n9898, QN => n16397);
   REGISTERS_reg_44_18_inst : DFF_X1 port map( D => n6032, CK => CLK, Q => 
                           n9899, QN => n16398);
   REGISTERS_reg_44_17_inst : DFF_X1 port map( D => n6031, CK => CLK, Q => 
                           n9900, QN => n16399);
   REGISTERS_reg_44_16_inst : DFF_X1 port map( D => n6030, CK => CLK, Q => 
                           n9901, QN => n16400);
   REGISTERS_reg_44_15_inst : DFF_X1 port map( D => n6029, CK => CLK, Q => 
                           n9902, QN => n16401);
   REGISTERS_reg_44_14_inst : DFF_X1 port map( D => n6028, CK => CLK, Q => 
                           n9903, QN => n16402);
   REGISTERS_reg_44_13_inst : DFF_X1 port map( D => n6027, CK => CLK, Q => 
                           n9904, QN => n16403);
   REGISTERS_reg_44_12_inst : DFF_X1 port map( D => n6026, CK => CLK, Q => 
                           n9905, QN => n16404);
   REGISTERS_reg_44_11_inst : DFF_X1 port map( D => n6025, CK => CLK, Q => 
                           n9906, QN => n16405);
   REGISTERS_reg_44_10_inst : DFF_X1 port map( D => n6024, CK => CLK, Q => 
                           n9907, QN => n16406);
   REGISTERS_reg_44_9_inst : DFF_X1 port map( D => n6023, CK => CLK, Q => n9908
                           , QN => n16407);
   REGISTERS_reg_44_8_inst : DFF_X1 port map( D => n6022, CK => CLK, Q => n9909
                           , QN => n16408);
   REGISTERS_reg_44_7_inst : DFF_X1 port map( D => n6021, CK => CLK, Q => n9910
                           , QN => n16409);
   REGISTERS_reg_44_6_inst : DFF_X1 port map( D => n6020, CK => CLK, Q => n9911
                           , QN => n16410);
   REGISTERS_reg_44_5_inst : DFF_X1 port map( D => n6019, CK => CLK, Q => n9912
                           , QN => n16411);
   REGISTERS_reg_44_4_inst : DFF_X1 port map( D => n6018, CK => CLK, Q => n9913
                           , QN => n16412);
   REGISTERS_reg_44_3_inst : DFF_X1 port map( D => n6017, CK => CLK, Q => n9914
                           , QN => n16413);
   REGISTERS_reg_44_2_inst : DFF_X1 port map( D => n6016, CK => CLK, Q => n9915
                           , QN => n16414);
   REGISTERS_reg_44_1_inst : DFF_X1 port map( D => n6015, CK => CLK, Q => n9916
                           , QN => n16415);
   REGISTERS_reg_44_0_inst : DFF_X1 port map( D => n6014, CK => CLK, Q => n9917
                           , QN => n16416);
   REGISTERS_reg_47_23_inst : DFF_X1 port map( D => n5941, CK => CLK, Q => 
                           n20478, QN => n16496);
   REGISTERS_reg_47_22_inst : DFF_X1 port map( D => n5940, CK => CLK, Q => 
                           n20477, QN => n16497);
   REGISTERS_reg_47_21_inst : DFF_X1 port map( D => n5939, CK => CLK, Q => 
                           n20476, QN => n16498);
   REGISTERS_reg_47_20_inst : DFF_X1 port map( D => n5938, CK => CLK, Q => 
                           n20475, QN => n16499);
   REGISTERS_reg_47_19_inst : DFF_X1 port map( D => n5937, CK => CLK, Q => 
                           n20474, QN => n16500);
   REGISTERS_reg_47_18_inst : DFF_X1 port map( D => n5936, CK => CLK, Q => 
                           n20473, QN => n16501);
   REGISTERS_reg_47_17_inst : DFF_X1 port map( D => n5935, CK => CLK, Q => 
                           n20472, QN => n16502);
   REGISTERS_reg_47_16_inst : DFF_X1 port map( D => n5934, CK => CLK, Q => 
                           n20471, QN => n16503);
   REGISTERS_reg_47_15_inst : DFF_X1 port map( D => n5933, CK => CLK, Q => 
                           n20470, QN => n16504);
   REGISTERS_reg_47_14_inst : DFF_X1 port map( D => n5932, CK => CLK, Q => 
                           n20469, QN => n16505);
   REGISTERS_reg_47_13_inst : DFF_X1 port map( D => n5931, CK => CLK, Q => 
                           n20468, QN => n16506);
   REGISTERS_reg_47_12_inst : DFF_X1 port map( D => n5930, CK => CLK, Q => 
                           n20467, QN => n16507);
   REGISTERS_reg_47_11_inst : DFF_X1 port map( D => n5929, CK => CLK, Q => 
                           n20466, QN => n16508);
   REGISTERS_reg_47_10_inst : DFF_X1 port map( D => n5928, CK => CLK, Q => 
                           n20465, QN => n16509);
   REGISTERS_reg_47_9_inst : DFF_X1 port map( D => n5927, CK => CLK, Q => 
                           n20464, QN => n16510);
   REGISTERS_reg_47_8_inst : DFF_X1 port map( D => n5926, CK => CLK, Q => 
                           n20463, QN => n16511);
   REGISTERS_reg_47_7_inst : DFF_X1 port map( D => n5925, CK => CLK, Q => 
                           n20462, QN => n16512);
   REGISTERS_reg_47_6_inst : DFF_X1 port map( D => n5924, CK => CLK, Q => 
                           n20461, QN => n16513);
   REGISTERS_reg_47_5_inst : DFF_X1 port map( D => n5923, CK => CLK, Q => 
                           n20460, QN => n16514);
   REGISTERS_reg_47_4_inst : DFF_X1 port map( D => n5922, CK => CLK, Q => 
                           n20459, QN => n16515);
   REGISTERS_reg_47_3_inst : DFF_X1 port map( D => n5921, CK => CLK, Q => 
                           n20458, QN => n16516);
   REGISTERS_reg_47_2_inst : DFF_X1 port map( D => n5920, CK => CLK, Q => 
                           n20457, QN => n16517);
   REGISTERS_reg_47_1_inst : DFF_X1 port map( D => n5919, CK => CLK, Q => 
                           n20456, QN => n16518);
   REGISTERS_reg_47_0_inst : DFF_X1 port map( D => n5918, CK => CLK, Q => 
                           n20455, QN => n16519);
   REGISTERS_reg_46_23_inst : DFF_X1 port map( D => n5973, CK => CLK, Q => 
                           n8662, QN => n16462);
   REGISTERS_reg_46_22_inst : DFF_X1 port map( D => n5972, CK => CLK, Q => 
                           n8673, QN => n16463);
   REGISTERS_reg_46_21_inst : DFF_X1 port map( D => n5971, CK => CLK, Q => 
                           n8684, QN => n16464);
   REGISTERS_reg_46_20_inst : DFF_X1 port map( D => n5970, CK => CLK, Q => 
                           n8695, QN => n16465);
   REGISTERS_reg_46_19_inst : DFF_X1 port map( D => n5969, CK => CLK, Q => 
                           n8706, QN => n16466);
   REGISTERS_reg_46_18_inst : DFF_X1 port map( D => n5968, CK => CLK, Q => 
                           n8717, QN => n16467);
   REGISTERS_reg_46_17_inst : DFF_X1 port map( D => n5967, CK => CLK, Q => 
                           n8728, QN => n16468);
   REGISTERS_reg_46_16_inst : DFF_X1 port map( D => n5966, CK => CLK, Q => 
                           n8739, QN => n16469);
   REGISTERS_reg_46_15_inst : DFF_X1 port map( D => n5965, CK => CLK, Q => 
                           n8750, QN => n16470);
   REGISTERS_reg_46_14_inst : DFF_X1 port map( D => n5964, CK => CLK, Q => 
                           n8761, QN => n16471);
   REGISTERS_reg_46_13_inst : DFF_X1 port map( D => n5963, CK => CLK, Q => 
                           n8772, QN => n16472);
   REGISTERS_reg_46_12_inst : DFF_X1 port map( D => n5962, CK => CLK, Q => 
                           n8783, QN => n16473);
   REGISTERS_reg_46_11_inst : DFF_X1 port map( D => n5961, CK => CLK, Q => 
                           n8794, QN => n16474);
   REGISTERS_reg_46_10_inst : DFF_X1 port map( D => n5960, CK => CLK, Q => 
                           n8805, QN => n16475);
   REGISTERS_reg_46_9_inst : DFF_X1 port map( D => n5959, CK => CLK, Q => n8816
                           , QN => n16476);
   REGISTERS_reg_46_8_inst : DFF_X1 port map( D => n5958, CK => CLK, Q => n8827
                           , QN => n16477);
   REGISTERS_reg_46_7_inst : DFF_X1 port map( D => n5957, CK => CLK, Q => n8838
                           , QN => n16478);
   REGISTERS_reg_46_6_inst : DFF_X1 port map( D => n5956, CK => CLK, Q => n8849
                           , QN => n16479);
   REGISTERS_reg_46_5_inst : DFF_X1 port map( D => n5955, CK => CLK, Q => n8860
                           , QN => n16480);
   REGISTERS_reg_46_4_inst : DFF_X1 port map( D => n5954, CK => CLK, Q => n8871
                           , QN => n16481);
   REGISTERS_reg_46_3_inst : DFF_X1 port map( D => n5953, CK => CLK, Q => n8882
                           , QN => n16482);
   REGISTERS_reg_46_2_inst : DFF_X1 port map( D => n5952, CK => CLK, Q => n8893
                           , QN => n16483);
   REGISTERS_reg_46_1_inst : DFF_X1 port map( D => n5951, CK => CLK, Q => n8904
                           , QN => n16484);
   REGISTERS_reg_46_0_inst : DFF_X1 port map( D => n5950, CK => CLK, Q => n8915
                           , QN => n16485);
   REGISTERS_reg_43_23_inst : DFF_X1 port map( D => n6069, CK => CLK, Q => 
                           n20454, QN => n16359);
   REGISTERS_reg_43_22_inst : DFF_X1 port map( D => n6068, CK => CLK, Q => 
                           n20453, QN => n16360);
   REGISTERS_reg_43_21_inst : DFF_X1 port map( D => n6067, CK => CLK, Q => 
                           n20452, QN => n16361);
   REGISTERS_reg_43_20_inst : DFF_X1 port map( D => n6066, CK => CLK, Q => 
                           n20451, QN => n16362);
   REGISTERS_reg_43_19_inst : DFF_X1 port map( D => n6065, CK => CLK, Q => 
                           n20450, QN => n16363);
   REGISTERS_reg_43_18_inst : DFF_X1 port map( D => n6064, CK => CLK, Q => 
                           n20449, QN => n16364);
   REGISTERS_reg_43_17_inst : DFF_X1 port map( D => n6063, CK => CLK, Q => 
                           n20448, QN => n16365);
   REGISTERS_reg_43_16_inst : DFF_X1 port map( D => n6062, CK => CLK, Q => 
                           n20447, QN => n16366);
   REGISTERS_reg_43_15_inst : DFF_X1 port map( D => n6061, CK => CLK, Q => 
                           n20446, QN => n16367);
   REGISTERS_reg_43_14_inst : DFF_X1 port map( D => n6060, CK => CLK, Q => 
                           n20445, QN => n16368);
   REGISTERS_reg_43_13_inst : DFF_X1 port map( D => n6059, CK => CLK, Q => 
                           n20444, QN => n16369);
   REGISTERS_reg_43_12_inst : DFF_X1 port map( D => n6058, CK => CLK, Q => 
                           n20443, QN => n16370);
   REGISTERS_reg_43_11_inst : DFF_X1 port map( D => n6057, CK => CLK, Q => 
                           n20442, QN => n16371);
   REGISTERS_reg_43_10_inst : DFF_X1 port map( D => n6056, CK => CLK, Q => 
                           n20441, QN => n16372);
   REGISTERS_reg_43_9_inst : DFF_X1 port map( D => n6055, CK => CLK, Q => 
                           n20440, QN => n16373);
   REGISTERS_reg_43_8_inst : DFF_X1 port map( D => n6054, CK => CLK, Q => 
                           n20439, QN => n16374);
   REGISTERS_reg_43_7_inst : DFF_X1 port map( D => n6053, CK => CLK, Q => 
                           n20438, QN => n16375);
   REGISTERS_reg_43_6_inst : DFF_X1 port map( D => n6052, CK => CLK, Q => 
                           n20437, QN => n16376);
   REGISTERS_reg_43_5_inst : DFF_X1 port map( D => n6051, CK => CLK, Q => 
                           n20436, QN => n16377);
   REGISTERS_reg_43_4_inst : DFF_X1 port map( D => n6050, CK => CLK, Q => 
                           n20435, QN => n16378);
   REGISTERS_reg_43_3_inst : DFF_X1 port map( D => n6049, CK => CLK, Q => 
                           n20434, QN => n16379);
   REGISTERS_reg_43_2_inst : DFF_X1 port map( D => n6048, CK => CLK, Q => 
                           n20433, QN => n16380);
   REGISTERS_reg_43_1_inst : DFF_X1 port map( D => n6047, CK => CLK, Q => 
                           n20432, QN => n16381);
   REGISTERS_reg_43_0_inst : DFF_X1 port map( D => n6046, CK => CLK, Q => 
                           n20431, QN => n16382);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n7381, CK => CLK, Q => n8974
                           , QN => n15167);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n7380, CK => CLK, Q => n8976
                           , QN => n15168);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n7379, CK => CLK, Q => n8978
                           , QN => n15169);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n7378, CK => CLK, Q => n8980
                           , QN => n15170);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n7377, CK => CLK, Q => n8982
                           , QN => n15171);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n7376, CK => CLK, Q => n8984
                           , QN => n15172);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n7375, CK => CLK, Q => n8986
                           , QN => n15173);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n7374, CK => CLK, Q => n8988
                           , QN => n15174);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n7373, CK => CLK, Q => n8990
                           , QN => n15175);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n7372, CK => CLK, Q => n8992
                           , QN => n15176);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n7371, CK => CLK, Q => n8994
                           , QN => n15177);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n7370, CK => CLK, Q => n8996
                           , QN => n15178);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n7369, CK => CLK, Q => n8998
                           , QN => n15179);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n7368, CK => CLK, Q => n9000
                           , QN => n15180);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n7367, CK => CLK, Q => n9002,
                           QN => n15181);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n7366, CK => CLK, Q => n9004,
                           QN => n15182);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n7365, CK => CLK, Q => n9006,
                           QN => n15183);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n7364, CK => CLK, Q => n9008,
                           QN => n15184);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n7363, CK => CLK, Q => n9010,
                           QN => n15185);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n7362, CK => CLK, Q => n9012,
                           QN => n15186);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n7361, CK => CLK, Q => n9014,
                           QN => n15187);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n7360, CK => CLK, Q => n9016,
                           QN => n15188);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n7359, CK => CLK, Q => n9018,
                           QN => n15189);
   REGISTERS_reg_60_23_inst : DFF_X1 port map( D => n5525, CK => CLK, Q => 
                           n9114, QN => n16769);
   REGISTERS_reg_60_22_inst : DFF_X1 port map( D => n5524, CK => CLK, Q => 
                           n9125, QN => n16770);
   REGISTERS_reg_60_21_inst : DFF_X1 port map( D => n5523, CK => CLK, Q => 
                           n9136, QN => n16771);
   REGISTERS_reg_60_20_inst : DFF_X1 port map( D => n5522, CK => CLK, Q => 
                           n9147, QN => n16772);
   REGISTERS_reg_60_19_inst : DFF_X1 port map( D => n5521, CK => CLK, Q => 
                           n9158, QN => n16773);
   REGISTERS_reg_60_18_inst : DFF_X1 port map( D => n5520, CK => CLK, Q => 
                           n9169, QN => n16774);
   REGISTERS_reg_60_17_inst : DFF_X1 port map( D => n5519, CK => CLK, Q => 
                           n9180, QN => n16775);
   REGISTERS_reg_60_16_inst : DFF_X1 port map( D => n5518, CK => CLK, Q => 
                           n9191, QN => n16776);
   REGISTERS_reg_60_15_inst : DFF_X1 port map( D => n5517, CK => CLK, Q => 
                           n9202, QN => n16777);
   REGISTERS_reg_60_14_inst : DFF_X1 port map( D => n5516, CK => CLK, Q => 
                           n9213, QN => n16778);
   REGISTERS_reg_60_13_inst : DFF_X1 port map( D => n5515, CK => CLK, Q => 
                           n9224, QN => n16779);
   REGISTERS_reg_60_12_inst : DFF_X1 port map( D => n5514, CK => CLK, Q => 
                           n9235, QN => n16780);
   REGISTERS_reg_60_11_inst : DFF_X1 port map( D => n5513, CK => CLK, Q => 
                           n9246, QN => n16781);
   REGISTERS_reg_60_10_inst : DFF_X1 port map( D => n5512, CK => CLK, Q => 
                           n9257, QN => n16782);
   REGISTERS_reg_60_9_inst : DFF_X1 port map( D => n5511, CK => CLK, Q => n9268
                           , QN => n16783);
   REGISTERS_reg_60_8_inst : DFF_X1 port map( D => n5510, CK => CLK, Q => n9279
                           , QN => n16784);
   REGISTERS_reg_60_7_inst : DFF_X1 port map( D => n5509, CK => CLK, Q => n9290
                           , QN => n16785);
   REGISTERS_reg_60_6_inst : DFF_X1 port map( D => n5508, CK => CLK, Q => n9301
                           , QN => n16786);
   REGISTERS_reg_60_5_inst : DFF_X1 port map( D => n5507, CK => CLK, Q => n9312
                           , QN => n16787);
   REGISTERS_reg_60_4_inst : DFF_X1 port map( D => n5506, CK => CLK, Q => n9323
                           , QN => n16788);
   REGISTERS_reg_60_3_inst : DFF_X1 port map( D => n5505, CK => CLK, Q => n9334
                           , QN => n16789);
   REGISTERS_reg_60_2_inst : DFF_X1 port map( D => n5504, CK => CLK, Q => n9345
                           , QN => n16790);
   REGISTERS_reg_60_1_inst : DFF_X1 port map( D => n5503, CK => CLK, Q => n9356
                           , QN => n16791);
   REGISTERS_reg_61_23_inst : DFF_X1 port map( D => n5493, CK => CLK, Q => 
                           n9118, QN => n16806);
   REGISTERS_reg_61_22_inst : DFF_X1 port map( D => n5492, CK => CLK, Q => 
                           n9129, QN => n16807);
   REGISTERS_reg_61_21_inst : DFF_X1 port map( D => n5491, CK => CLK, Q => 
                           n9140, QN => n16808);
   REGISTERS_reg_61_20_inst : DFF_X1 port map( D => n5490, CK => CLK, Q => 
                           n9151, QN => n16809);
   REGISTERS_reg_61_19_inst : DFF_X1 port map( D => n5489, CK => CLK, Q => 
                           n9162, QN => n16810);
   REGISTERS_reg_61_18_inst : DFF_X1 port map( D => n5488, CK => CLK, Q => 
                           n9173, QN => n16811);
   REGISTERS_reg_61_17_inst : DFF_X1 port map( D => n5487, CK => CLK, Q => 
                           n9184, QN => n16812);
   REGISTERS_reg_61_16_inst : DFF_X1 port map( D => n5486, CK => CLK, Q => 
                           n9195, QN => n16813);
   REGISTERS_reg_61_15_inst : DFF_X1 port map( D => n5485, CK => CLK, Q => 
                           n9206, QN => n16814);
   REGISTERS_reg_61_14_inst : DFF_X1 port map( D => n5484, CK => CLK, Q => 
                           n9217, QN => n16815);
   REGISTERS_reg_61_13_inst : DFF_X1 port map( D => n5483, CK => CLK, Q => 
                           n9228, QN => n16816);
   REGISTERS_reg_61_12_inst : DFF_X1 port map( D => n5482, CK => CLK, Q => 
                           n9239, QN => n16817);
   REGISTERS_reg_61_11_inst : DFF_X1 port map( D => n5481, CK => CLK, Q => 
                           n9250, QN => n16818);
   REGISTERS_reg_61_10_inst : DFF_X1 port map( D => n5480, CK => CLK, Q => 
                           n9261, QN => n16819);
   REGISTERS_reg_61_9_inst : DFF_X1 port map( D => n5479, CK => CLK, Q => n9272
                           , QN => n16820);
   REGISTERS_reg_61_8_inst : DFF_X1 port map( D => n5478, CK => CLK, Q => n9283
                           , QN => n16821);
   REGISTERS_reg_61_7_inst : DFF_X1 port map( D => n5477, CK => CLK, Q => n9294
                           , QN => n16822);
   REGISTERS_reg_61_6_inst : DFF_X1 port map( D => n5476, CK => CLK, Q => n9305
                           , QN => n16823);
   REGISTERS_reg_61_5_inst : DFF_X1 port map( D => n5475, CK => CLK, Q => n9316
                           , QN => n16824);
   REGISTERS_reg_61_4_inst : DFF_X1 port map( D => n5474, CK => CLK, Q => n9327
                           , QN => n16825);
   REGISTERS_reg_61_3_inst : DFF_X1 port map( D => n5473, CK => CLK, Q => n9338
                           , QN => n16826);
   REGISTERS_reg_61_2_inst : DFF_X1 port map( D => n5472, CK => CLK, Q => n9349
                           , QN => n16827);
   REGISTERS_reg_61_1_inst : DFF_X1 port map( D => n5471, CK => CLK, Q => n9360
                           , QN => n16828);
   REGISTERS_reg_39_23_inst : DFF_X1 port map( D => n6197, CK => CLK, Q => 
                           n20430, QN => n16318);
   REGISTERS_reg_39_22_inst : DFF_X1 port map( D => n6196, CK => CLK, Q => 
                           n20429, QN => n16319);
   REGISTERS_reg_39_21_inst : DFF_X1 port map( D => n6195, CK => CLK, Q => 
                           n20428, QN => n16320);
   REGISTERS_reg_39_20_inst : DFF_X1 port map( D => n6194, CK => CLK, Q => 
                           n20427, QN => n16321);
   REGISTERS_reg_39_19_inst : DFF_X1 port map( D => n6193, CK => CLK, Q => 
                           n20426, QN => n16322);
   REGISTERS_reg_39_18_inst : DFF_X1 port map( D => n6192, CK => CLK, Q => 
                           n20425, QN => n16323);
   REGISTERS_reg_39_17_inst : DFF_X1 port map( D => n6191, CK => CLK, Q => 
                           n20424, QN => n16324);
   REGISTERS_reg_39_16_inst : DFF_X1 port map( D => n6190, CK => CLK, Q => 
                           n20423, QN => n16325);
   REGISTERS_reg_39_15_inst : DFF_X1 port map( D => n6189, CK => CLK, Q => 
                           n20422, QN => n16326);
   REGISTERS_reg_39_14_inst : DFF_X1 port map( D => n6188, CK => CLK, Q => 
                           n20421, QN => n16327);
   REGISTERS_reg_39_13_inst : DFF_X1 port map( D => n6187, CK => CLK, Q => 
                           n20420, QN => n16328);
   REGISTERS_reg_39_12_inst : DFF_X1 port map( D => n6186, CK => CLK, Q => 
                           n20419, QN => n16329);
   REGISTERS_reg_39_11_inst : DFF_X1 port map( D => n6185, CK => CLK, Q => 
                           n20418, QN => n16330);
   REGISTERS_reg_39_10_inst : DFF_X1 port map( D => n6184, CK => CLK, Q => 
                           n20417, QN => n16331);
   REGISTERS_reg_39_9_inst : DFF_X1 port map( D => n6183, CK => CLK, Q => 
                           n20416, QN => n16332);
   REGISTERS_reg_39_8_inst : DFF_X1 port map( D => n6182, CK => CLK, Q => 
                           n20415, QN => n16333);
   REGISTERS_reg_39_7_inst : DFF_X1 port map( D => n6181, CK => CLK, Q => 
                           n20414, QN => n16334);
   REGISTERS_reg_39_6_inst : DFF_X1 port map( D => n6180, CK => CLK, Q => 
                           n20413, QN => n16335);
   REGISTERS_reg_39_5_inst : DFF_X1 port map( D => n6179, CK => CLK, Q => 
                           n20412, QN => n16336);
   REGISTERS_reg_39_4_inst : DFF_X1 port map( D => n6178, CK => CLK, Q => 
                           n20411, QN => n16337);
   REGISTERS_reg_39_3_inst : DFF_X1 port map( D => n6177, CK => CLK, Q => 
                           n20410, QN => n16338);
   REGISTERS_reg_39_2_inst : DFF_X1 port map( D => n6176, CK => CLK, Q => 
                           n20409, QN => n16339);
   REGISTERS_reg_39_1_inst : DFF_X1 port map( D => n6175, CK => CLK, Q => 
                           n20408, QN => n16340);
   REGISTERS_reg_39_0_inst : DFF_X1 port map( D => n6174, CK => CLK, Q => 
                           n20407, QN => n16341);
   REGISTERS_reg_35_23_inst : DFF_X1 port map( D => n6325, CK => CLK, Q => 
                           n20406, QN => n16180);
   REGISTERS_reg_35_22_inst : DFF_X1 port map( D => n6324, CK => CLK, Q => 
                           n20405, QN => n16181);
   REGISTERS_reg_35_21_inst : DFF_X1 port map( D => n6323, CK => CLK, Q => 
                           n20404, QN => n16182);
   REGISTERS_reg_35_20_inst : DFF_X1 port map( D => n6322, CK => CLK, Q => 
                           n20403, QN => n16183);
   REGISTERS_reg_35_19_inst : DFF_X1 port map( D => n6321, CK => CLK, Q => 
                           n20402, QN => n16184);
   REGISTERS_reg_35_18_inst : DFF_X1 port map( D => n6320, CK => CLK, Q => 
                           n20401, QN => n16185);
   REGISTERS_reg_35_17_inst : DFF_X1 port map( D => n6319, CK => CLK, Q => 
                           n20400, QN => n16186);
   REGISTERS_reg_35_16_inst : DFF_X1 port map( D => n6318, CK => CLK, Q => 
                           n20399, QN => n16187);
   REGISTERS_reg_35_15_inst : DFF_X1 port map( D => n6317, CK => CLK, Q => 
                           n20398, QN => n16188);
   REGISTERS_reg_35_14_inst : DFF_X1 port map( D => n6316, CK => CLK, Q => 
                           n20397, QN => n16189);
   REGISTERS_reg_35_13_inst : DFF_X1 port map( D => n6315, CK => CLK, Q => 
                           n20396, QN => n16190);
   REGISTERS_reg_35_12_inst : DFF_X1 port map( D => n6314, CK => CLK, Q => 
                           n20395, QN => n16191);
   REGISTERS_reg_35_11_inst : DFF_X1 port map( D => n6313, CK => CLK, Q => 
                           n20394, QN => n16192);
   REGISTERS_reg_35_10_inst : DFF_X1 port map( D => n6312, CK => CLK, Q => 
                           n20393, QN => n16193);
   REGISTERS_reg_35_9_inst : DFF_X1 port map( D => n6311, CK => CLK, Q => 
                           n20392, QN => n16194);
   REGISTERS_reg_35_8_inst : DFF_X1 port map( D => n6310, CK => CLK, Q => 
                           n20391, QN => n16195);
   REGISTERS_reg_35_7_inst : DFF_X1 port map( D => n6309, CK => CLK, Q => 
                           n20390, QN => n16196);
   REGISTERS_reg_35_6_inst : DFF_X1 port map( D => n6308, CK => CLK, Q => 
                           n20389, QN => n16197);
   REGISTERS_reg_35_5_inst : DFF_X1 port map( D => n6307, CK => CLK, Q => 
                           n20388, QN => n16198);
   REGISTERS_reg_35_4_inst : DFF_X1 port map( D => n6306, CK => CLK, Q => 
                           n20387, QN => n16199);
   REGISTERS_reg_35_3_inst : DFF_X1 port map( D => n6305, CK => CLK, Q => 
                           n20386, QN => n16200);
   REGISTERS_reg_35_2_inst : DFF_X1 port map( D => n6304, CK => CLK, Q => 
                           n20385, QN => n16201);
   REGISTERS_reg_35_1_inst : DFF_X1 port map( D => n6303, CK => CLK, Q => 
                           n20384, QN => n16202);
   REGISTERS_reg_35_0_inst : DFF_X1 port map( D => n6302, CK => CLK, Q => 
                           n20383, QN => n16203);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n6453, CK => CLK, Q => 
                           n20382, QN => n16075);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n6452, CK => CLK, Q => 
                           n20381, QN => n16076);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n6451, CK => CLK, Q => 
                           n20380, QN => n16077);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n6450, CK => CLK, Q => 
                           n20379, QN => n16078);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n6449, CK => CLK, Q => 
                           n20378, QN => n16079);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n6448, CK => CLK, Q => 
                           n20377, QN => n16080);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n6447, CK => CLK, Q => 
                           n20376, QN => n16081);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n6446, CK => CLK, Q => 
                           n20375, QN => n16082);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n6445, CK => CLK, Q => 
                           n20374, QN => n16083);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n6444, CK => CLK, Q => 
                           n20373, QN => n16084);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n6443, CK => CLK, Q => 
                           n20372, QN => n16085);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n6442, CK => CLK, Q => 
                           n20371, QN => n16086);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n6441, CK => CLK, Q => 
                           n20370, QN => n16087);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n6440, CK => CLK, Q => 
                           n20369, QN => n16088);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n6439, CK => CLK, Q => 
                           n20368, QN => n16089);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n6438, CK => CLK, Q => 
                           n20367, QN => n16090);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n6437, CK => CLK, Q => 
                           n20366, QN => n16091);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n6436, CK => CLK, Q => 
                           n20365, QN => n16092);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n6435, CK => CLK, Q => 
                           n20364, QN => n16093);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n6434, CK => CLK, Q => 
                           n20363, QN => n16094);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n6433, CK => CLK, Q => 
                           n20362, QN => n16095);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n6432, CK => CLK, Q => 
                           n20361, QN => n16096);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n6431, CK => CLK, Q => 
                           n20360, QN => n16097);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n6430, CK => CLK, Q => 
                           n20359, QN => n16098);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n6581, CK => CLK, Q => 
                           n9510, QN => n15938);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n6580, CK => CLK, Q => 
                           n9511, QN => n15939);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n6579, CK => CLK, Q => 
                           n9512, QN => n15940);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n6578, CK => CLK, Q => 
                           n9513, QN => n15941);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n6577, CK => CLK, Q => 
                           n9514, QN => n15942);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n6576, CK => CLK, Q => 
                           n9515, QN => n15943);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n6575, CK => CLK, Q => 
                           n9516, QN => n15944);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n6574, CK => CLK, Q => 
                           n9517, QN => n15945);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n6573, CK => CLK, Q => 
                           n9518, QN => n15946);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n6572, CK => CLK, Q => 
                           n9519, QN => n15947);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n6571, CK => CLK, Q => 
                           n9520, QN => n15948);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n6570, CK => CLK, Q => 
                           n9521, QN => n15949);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n6569, CK => CLK, Q => 
                           n9522, QN => n15950);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n6568, CK => CLK, Q => 
                           n9523, QN => n15951);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n6567, CK => CLK, Q => n9524
                           , QN => n15952);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n6566, CK => CLK, Q => n9525
                           , QN => n15953);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n6565, CK => CLK, Q => n9526
                           , QN => n15954);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n6564, CK => CLK, Q => n9527
                           , QN => n15955);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n6563, CK => CLK, Q => n9528
                           , QN => n15956);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n6562, CK => CLK, Q => n9529
                           , QN => n15957);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n6561, CK => CLK, Q => n9530
                           , QN => n15958);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n6560, CK => CLK, Q => n9531
                           , QN => n15959);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n6559, CK => CLK, Q => n9532
                           , QN => n15960);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n6558, CK => CLK, Q => n9533
                           , QN => n15961);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n6709, CK => CLK, Q => 
                           n9606, QN => n15865);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n6708, CK => CLK, Q => 
                           n9607, QN => n15866);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n6707, CK => CLK, Q => 
                           n9608, QN => n15867);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n6706, CK => CLK, Q => 
                           n9609, QN => n15868);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n6705, CK => CLK, Q => 
                           n9610, QN => n15869);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n6704, CK => CLK, Q => 
                           n9611, QN => n15870);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n6703, CK => CLK, Q => 
                           n9612, QN => n15871);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n6702, CK => CLK, Q => 
                           n9613, QN => n15872);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n6701, CK => CLK, Q => 
                           n9614, QN => n15873);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n6700, CK => CLK, Q => 
                           n9615, QN => n15874);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n6699, CK => CLK, Q => 
                           n9616, QN => n15875);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n6698, CK => CLK, Q => 
                           n9617, QN => n15876);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n6697, CK => CLK, Q => 
                           n9618, QN => n15877);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n6696, CK => CLK, Q => 
                           n9619, QN => n15878);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n6695, CK => CLK, Q => n9620
                           , QN => n15879);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n6694, CK => CLK, Q => n9621
                           , QN => n15880);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n6693, CK => CLK, Q => n9622
                           , QN => n15881);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n6692, CK => CLK, Q => n9623
                           , QN => n15882);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n6691, CK => CLK, Q => n9624
                           , QN => n15883);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n6690, CK => CLK, Q => n9625
                           , QN => n15884);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n6689, CK => CLK, Q => n9626
                           , QN => n15885);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n6688, CK => CLK, Q => n9627
                           , QN => n15886);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n6687, CK => CLK, Q => n9628
                           , QN => n15887);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n6686, CK => CLK, Q => n9629
                           , QN => n15888);
   REGISTERS_reg_45_23_inst : DFF_X1 port map( D => n6005, CK => CLK, Q => 
                           n9926, QN => n16428);
   REGISTERS_reg_45_22_inst : DFF_X1 port map( D => n6004, CK => CLK, Q => 
                           n9927, QN => n16429);
   REGISTERS_reg_45_21_inst : DFF_X1 port map( D => n6003, CK => CLK, Q => 
                           n9928, QN => n16430);
   REGISTERS_reg_45_20_inst : DFF_X1 port map( D => n6002, CK => CLK, Q => 
                           n9929, QN => n16431);
   REGISTERS_reg_45_19_inst : DFF_X1 port map( D => n6001, CK => CLK, Q => 
                           n9930, QN => n16432);
   REGISTERS_reg_45_18_inst : DFF_X1 port map( D => n6000, CK => CLK, Q => 
                           n9931, QN => n16433);
   REGISTERS_reg_45_17_inst : DFF_X1 port map( D => n5999, CK => CLK, Q => 
                           n9932, QN => n16434);
   REGISTERS_reg_45_16_inst : DFF_X1 port map( D => n5998, CK => CLK, Q => 
                           n9933, QN => n16435);
   REGISTERS_reg_45_15_inst : DFF_X1 port map( D => n5997, CK => CLK, Q => 
                           n9934, QN => n16436);
   REGISTERS_reg_45_14_inst : DFF_X1 port map( D => n5996, CK => CLK, Q => 
                           n9935, QN => n16437);
   REGISTERS_reg_45_13_inst : DFF_X1 port map( D => n5995, CK => CLK, Q => 
                           n9936, QN => n16438);
   REGISTERS_reg_45_12_inst : DFF_X1 port map( D => n5994, CK => CLK, Q => 
                           n9937, QN => n16439);
   REGISTERS_reg_45_11_inst : DFF_X1 port map( D => n5993, CK => CLK, Q => 
                           n9938, QN => n16440);
   REGISTERS_reg_45_10_inst : DFF_X1 port map( D => n5992, CK => CLK, Q => 
                           n9939, QN => n16441);
   REGISTERS_reg_45_9_inst : DFF_X1 port map( D => n5991, CK => CLK, Q => n9940
                           , QN => n16442);
   REGISTERS_reg_45_8_inst : DFF_X1 port map( D => n5990, CK => CLK, Q => n9941
                           , QN => n16443);
   REGISTERS_reg_45_7_inst : DFF_X1 port map( D => n5989, CK => CLK, Q => n9942
                           , QN => n16444);
   REGISTERS_reg_45_6_inst : DFF_X1 port map( D => n5988, CK => CLK, Q => n9943
                           , QN => n16445);
   REGISTERS_reg_45_5_inst : DFF_X1 port map( D => n5987, CK => CLK, Q => n9944
                           , QN => n16446);
   REGISTERS_reg_45_4_inst : DFF_X1 port map( D => n5986, CK => CLK, Q => n9945
                           , QN => n16447);
   REGISTERS_reg_45_3_inst : DFF_X1 port map( D => n5985, CK => CLK, Q => n9946
                           , QN => n16448);
   REGISTERS_reg_45_2_inst : DFF_X1 port map( D => n5984, CK => CLK, Q => n9947
                           , QN => n16449);
   REGISTERS_reg_45_1_inst : DFF_X1 port map( D => n5983, CK => CLK, Q => n9948
                           , QN => n16450);
   REGISTERS_reg_45_0_inst : DFF_X1 port map( D => n5982, CK => CLK, Q => n9949
                           , QN => n16451);
   REGISTERS_reg_38_23_inst : DFF_X1 port map( D => n6229, CK => CLK, Q => 
                           n8663, QN => n16284);
   REGISTERS_reg_38_22_inst : DFF_X1 port map( D => n6228, CK => CLK, Q => 
                           n8674, QN => n16285);
   REGISTERS_reg_38_21_inst : DFF_X1 port map( D => n6227, CK => CLK, Q => 
                           n8685, QN => n16286);
   REGISTERS_reg_38_20_inst : DFF_X1 port map( D => n6226, CK => CLK, Q => 
                           n8696, QN => n16287);
   REGISTERS_reg_38_19_inst : DFF_X1 port map( D => n6225, CK => CLK, Q => 
                           n8707, QN => n16288);
   REGISTERS_reg_38_18_inst : DFF_X1 port map( D => n6224, CK => CLK, Q => 
                           n8718, QN => n16289);
   REGISTERS_reg_38_17_inst : DFF_X1 port map( D => n6223, CK => CLK, Q => 
                           n8729, QN => n16290);
   REGISTERS_reg_38_16_inst : DFF_X1 port map( D => n6222, CK => CLK, Q => 
                           n8740, QN => n16291);
   REGISTERS_reg_38_15_inst : DFF_X1 port map( D => n6221, CK => CLK, Q => 
                           n8751, QN => n16292);
   REGISTERS_reg_38_14_inst : DFF_X1 port map( D => n6220, CK => CLK, Q => 
                           n8762, QN => n16293);
   REGISTERS_reg_38_13_inst : DFF_X1 port map( D => n6219, CK => CLK, Q => 
                           n8773, QN => n16294);
   REGISTERS_reg_38_12_inst : DFF_X1 port map( D => n6218, CK => CLK, Q => 
                           n8784, QN => n16295);
   REGISTERS_reg_38_11_inst : DFF_X1 port map( D => n6217, CK => CLK, Q => 
                           n8795, QN => n16296);
   REGISTERS_reg_38_10_inst : DFF_X1 port map( D => n6216, CK => CLK, Q => 
                           n8806, QN => n16297);
   REGISTERS_reg_38_9_inst : DFF_X1 port map( D => n6215, CK => CLK, Q => n8817
                           , QN => n16298);
   REGISTERS_reg_38_8_inst : DFF_X1 port map( D => n6214, CK => CLK, Q => n8828
                           , QN => n16299);
   REGISTERS_reg_38_7_inst : DFF_X1 port map( D => n6213, CK => CLK, Q => n8839
                           , QN => n16300);
   REGISTERS_reg_38_6_inst : DFF_X1 port map( D => n6212, CK => CLK, Q => n8850
                           , QN => n16301);
   REGISTERS_reg_38_5_inst : DFF_X1 port map( D => n6211, CK => CLK, Q => n8861
                           , QN => n16302);
   REGISTERS_reg_38_4_inst : DFF_X1 port map( D => n6210, CK => CLK, Q => n8872
                           , QN => n16303);
   REGISTERS_reg_38_3_inst : DFF_X1 port map( D => n6209, CK => CLK, Q => n8883
                           , QN => n16304);
   REGISTERS_reg_38_2_inst : DFF_X1 port map( D => n6208, CK => CLK, Q => n8894
                           , QN => n16305);
   REGISTERS_reg_38_1_inst : DFF_X1 port map( D => n6207, CK => CLK, Q => n8905
                           , QN => n16306);
   REGISTERS_reg_38_0_inst : DFF_X1 port map( D => n6206, CK => CLK, Q => n8916
                           , QN => n16307);
   REGISTERS_reg_37_23_inst : DFF_X1 port map( D => n6261, CK => CLK, Q => 
                           n20358, QN => n16250);
   REGISTERS_reg_37_22_inst : DFF_X1 port map( D => n6260, CK => CLK, Q => 
                           n20357, QN => n16251);
   REGISTERS_reg_37_21_inst : DFF_X1 port map( D => n6259, CK => CLK, Q => 
                           n20356, QN => n16252);
   REGISTERS_reg_37_20_inst : DFF_X1 port map( D => n6258, CK => CLK, Q => 
                           n20355, QN => n16253);
   REGISTERS_reg_37_19_inst : DFF_X1 port map( D => n6257, CK => CLK, Q => 
                           n20354, QN => n16254);
   REGISTERS_reg_37_18_inst : DFF_X1 port map( D => n6256, CK => CLK, Q => 
                           n20353, QN => n16255);
   REGISTERS_reg_37_17_inst : DFF_X1 port map( D => n6255, CK => CLK, Q => 
                           n20352, QN => n16256);
   REGISTERS_reg_37_16_inst : DFF_X1 port map( D => n6254, CK => CLK, Q => 
                           n20351, QN => n16257);
   REGISTERS_reg_37_15_inst : DFF_X1 port map( D => n6253, CK => CLK, Q => 
                           n20350, QN => n16258);
   REGISTERS_reg_37_14_inst : DFF_X1 port map( D => n6252, CK => CLK, Q => 
                           n20349, QN => n16259);
   REGISTERS_reg_37_13_inst : DFF_X1 port map( D => n6251, CK => CLK, Q => 
                           n20348, QN => n16260);
   REGISTERS_reg_37_12_inst : DFF_X1 port map( D => n6250, CK => CLK, Q => 
                           n20347, QN => n16261);
   REGISTERS_reg_37_11_inst : DFF_X1 port map( D => n6249, CK => CLK, Q => 
                           n20346, QN => n16262);
   REGISTERS_reg_37_10_inst : DFF_X1 port map( D => n6248, CK => CLK, Q => 
                           n20345, QN => n16263);
   REGISTERS_reg_37_9_inst : DFF_X1 port map( D => n6247, CK => CLK, Q => 
                           n20344, QN => n16264);
   REGISTERS_reg_37_8_inst : DFF_X1 port map( D => n6246, CK => CLK, Q => 
                           n20343, QN => n16265);
   REGISTERS_reg_37_7_inst : DFF_X1 port map( D => n6245, CK => CLK, Q => 
                           n20342, QN => n16266);
   REGISTERS_reg_37_6_inst : DFF_X1 port map( D => n6244, CK => CLK, Q => 
                           n20341, QN => n16267);
   REGISTERS_reg_37_5_inst : DFF_X1 port map( D => n6243, CK => CLK, Q => 
                           n20340, QN => n16268);
   REGISTERS_reg_37_4_inst : DFF_X1 port map( D => n6242, CK => CLK, Q => 
                           n20339, QN => n16269);
   REGISTERS_reg_37_3_inst : DFF_X1 port map( D => n6241, CK => CLK, Q => 
                           n20338, QN => n16270);
   REGISTERS_reg_37_2_inst : DFF_X1 port map( D => n6240, CK => CLK, Q => 
                           n20337, QN => n16271);
   REGISTERS_reg_37_1_inst : DFF_X1 port map( D => n6239, CK => CLK, Q => 
                           n20336, QN => n16272);
   REGISTERS_reg_37_0_inst : DFF_X1 port map( D => n6238, CK => CLK, Q => 
                           n20335, QN => n16273);
   REGISTERS_reg_36_23_inst : DFF_X1 port map( D => n6293, CK => CLK, Q => 
                           n20334, QN => n16215);
   REGISTERS_reg_36_22_inst : DFF_X1 port map( D => n6292, CK => CLK, Q => 
                           n20333, QN => n16216);
   REGISTERS_reg_36_21_inst : DFF_X1 port map( D => n6291, CK => CLK, Q => 
                           n20332, QN => n16217);
   REGISTERS_reg_36_20_inst : DFF_X1 port map( D => n6290, CK => CLK, Q => 
                           n20331, QN => n16218);
   REGISTERS_reg_36_19_inst : DFF_X1 port map( D => n6289, CK => CLK, Q => 
                           n20330, QN => n16219);
   REGISTERS_reg_36_18_inst : DFF_X1 port map( D => n6288, CK => CLK, Q => 
                           n20329, QN => n16220);
   REGISTERS_reg_36_17_inst : DFF_X1 port map( D => n6287, CK => CLK, Q => 
                           n20328, QN => n16221);
   REGISTERS_reg_36_16_inst : DFF_X1 port map( D => n6286, CK => CLK, Q => 
                           n20327, QN => n16222);
   REGISTERS_reg_36_15_inst : DFF_X1 port map( D => n6285, CK => CLK, Q => 
                           n20326, QN => n16223);
   REGISTERS_reg_36_14_inst : DFF_X1 port map( D => n6284, CK => CLK, Q => 
                           n20325, QN => n16224);
   REGISTERS_reg_36_13_inst : DFF_X1 port map( D => n6283, CK => CLK, Q => 
                           n20324, QN => n16225);
   REGISTERS_reg_36_12_inst : DFF_X1 port map( D => n6282, CK => CLK, Q => 
                           n20323, QN => n16226);
   REGISTERS_reg_36_11_inst : DFF_X1 port map( D => n6281, CK => CLK, Q => 
                           n20322, QN => n16227);
   REGISTERS_reg_36_10_inst : DFF_X1 port map( D => n6280, CK => CLK, Q => 
                           n20321, QN => n16228);
   REGISTERS_reg_36_9_inst : DFF_X1 port map( D => n6279, CK => CLK, Q => 
                           n20320, QN => n16229);
   REGISTERS_reg_36_8_inst : DFF_X1 port map( D => n6278, CK => CLK, Q => 
                           n20319, QN => n16230);
   REGISTERS_reg_36_7_inst : DFF_X1 port map( D => n6277, CK => CLK, Q => 
                           n20318, QN => n16231);
   REGISTERS_reg_36_6_inst : DFF_X1 port map( D => n6276, CK => CLK, Q => 
                           n20317, QN => n16232);
   REGISTERS_reg_36_5_inst : DFF_X1 port map( D => n6275, CK => CLK, Q => 
                           n20316, QN => n16233);
   REGISTERS_reg_36_4_inst : DFF_X1 port map( D => n6274, CK => CLK, Q => 
                           n20315, QN => n16234);
   REGISTERS_reg_36_3_inst : DFF_X1 port map( D => n6273, CK => CLK, Q => 
                           n20314, QN => n16235);
   REGISTERS_reg_36_2_inst : DFF_X1 port map( D => n6272, CK => CLK, Q => 
                           n20313, QN => n16236);
   REGISTERS_reg_36_1_inst : DFF_X1 port map( D => n6271, CK => CLK, Q => 
                           n20312, QN => n16237);
   REGISTERS_reg_36_0_inst : DFF_X1 port map( D => n6270, CK => CLK, Q => 
                           n20311, QN => n16238);
   REGISTERS_reg_33_23_inst : DFF_X1 port map( D => n6389, CK => CLK, Q => 
                           n20310, QN => n16144);
   REGISTERS_reg_33_22_inst : DFF_X1 port map( D => n6388, CK => CLK, Q => 
                           n20309, QN => n16145);
   REGISTERS_reg_33_21_inst : DFF_X1 port map( D => n6387, CK => CLK, Q => 
                           n20308, QN => n16146);
   U13042 : INV_X1 port map( A => ADD_RD1(2), ZN => n19661);
   U13043 : INV_X1 port map( A => ADD_RD2(2), ZN => n18394);
   U13044 : INV_X1 port map( A => n21909, ZN => n21902);
   U13045 : INV_X1 port map( A => n22017, ZN => n22010);
   U13046 : INV_X1 port map( A => n22161, ZN => n22154);
   U13047 : INV_X1 port map( A => n22574, ZN => n22567);
   U13048 : INV_X1 port map( A => n21837, ZN => n21830);
   U13049 : INV_X1 port map( A => n21873, ZN => n21866);
   U13050 : INV_X1 port map( A => n21945, ZN => n21938);
   U13051 : INV_X1 port map( A => n21981, ZN => n21974);
   U13052 : INV_X1 port map( A => n22053, ZN => n22046);
   U13053 : INV_X1 port map( A => n22089, ZN => n22082);
   U13054 : INV_X1 port map( A => n22125, ZN => n22118);
   U13055 : INV_X1 port map( A => n22197, ZN => n22190);
   U13056 : INV_X1 port map( A => n22233, ZN => n22226);
   U13057 : INV_X1 port map( A => n22269, ZN => n22262);
   U13058 : INV_X1 port map( A => n22305, ZN => n22298);
   U13059 : INV_X1 port map( A => n22341, ZN => n22334);
   U13060 : INV_X1 port map( A => n21810, ZN => n21801);
   U13061 : INV_X1 port map( A => n21819, ZN => n21812);
   U13062 : INV_X1 port map( A => n21846, ZN => n21839);
   U13063 : INV_X1 port map( A => n21891, ZN => n21884);
   U13064 : INV_X1 port map( A => n21900, ZN => n21893);
   U13065 : INV_X1 port map( A => n21918, ZN => n21911);
   U13066 : INV_X1 port map( A => n21999, ZN => n21992);
   U13067 : INV_X1 port map( A => n22008, ZN => n22001);
   U13068 : INV_X1 port map( A => n22071, ZN => n22064);
   U13069 : INV_X1 port map( A => n22152, ZN => n22145);
   U13070 : INV_X1 port map( A => n22206, ZN => n22199);
   U13071 : INV_X1 port map( A => n22368, ZN => n22361);
   U13072 : INV_X1 port map( A => n21936, ZN => n21929);
   U13073 : INV_X1 port map( A => n21828, ZN => n21821);
   U13074 : INV_X1 port map( A => n21855, ZN => n21848);
   U13075 : INV_X1 port map( A => n21864, ZN => n21857);
   U13076 : INV_X1 port map( A => n21882, ZN => n21875);
   U13077 : INV_X1 port map( A => n21927, ZN => n21920);
   U13078 : INV_X1 port map( A => n21954, ZN => n21947);
   U13079 : INV_X1 port map( A => n21963, ZN => n21956);
   U13080 : INV_X1 port map( A => n21972, ZN => n21965);
   U13081 : INV_X1 port map( A => n21990, ZN => n21983);
   U13082 : INV_X1 port map( A => n22026, ZN => n22019);
   U13083 : INV_X1 port map( A => n22035, ZN => n22028);
   U13084 : INV_X1 port map( A => n22044, ZN => n22037);
   U13085 : INV_X1 port map( A => n22062, ZN => n22055);
   U13086 : INV_X1 port map( A => n22080, ZN => n22073);
   U13087 : INV_X1 port map( A => n22098, ZN => n22091);
   U13088 : INV_X1 port map( A => n22107, ZN => n22100);
   U13089 : INV_X1 port map( A => n22116, ZN => n22109);
   U13090 : INV_X1 port map( A => n22134, ZN => n22127);
   U13091 : INV_X1 port map( A => n22143, ZN => n22136);
   U13092 : INV_X1 port map( A => n22170, ZN => n22163);
   U13093 : INV_X1 port map( A => n22179, ZN => n22172);
   U13094 : INV_X1 port map( A => n22188, ZN => n22181);
   U13095 : INV_X1 port map( A => n22215, ZN => n22208);
   U13096 : INV_X1 port map( A => n22224, ZN => n22217);
   U13097 : INV_X1 port map( A => n22242, ZN => n22235);
   U13098 : INV_X1 port map( A => n22251, ZN => n22244);
   U13099 : INV_X1 port map( A => n22260, ZN => n22253);
   U13100 : INV_X1 port map( A => n22278, ZN => n22271);
   U13101 : INV_X1 port map( A => n22287, ZN => n22280);
   U13102 : INV_X1 port map( A => n22296, ZN => n22289);
   U13103 : INV_X1 port map( A => n22314, ZN => n22307);
   U13104 : INV_X1 port map( A => n22323, ZN => n22316);
   U13105 : INV_X1 port map( A => n22332, ZN => n22325);
   U13106 : INV_X1 port map( A => n22350, ZN => n22343);
   U13107 : INV_X1 port map( A => n22359, ZN => n22352);
   U13108 : BUF_X1 port map( A => n18496, Z => n20839);
   U13109 : BUF_X1 port map( A => n18496, Z => n20840);
   U13110 : BUF_X1 port map( A => n16922, Z => n21396);
   U13111 : BUF_X1 port map( A => n16922, Z => n21397);
   U13112 : BUF_X1 port map( A => n18457, Z => n21107);
   U13113 : BUF_X1 port map( A => n18457, Z => n21108);
   U13114 : BUF_X1 port map( A => n16876, Z => n21664);
   U13115 : BUF_X1 port map( A => n16876, Z => n21665);
   U13116 : BUF_X1 port map( A => n18496, Z => n20841);
   U13117 : BUF_X1 port map( A => n16922, Z => n21398);
   U13118 : BUF_X1 port map( A => n18457, Z => n21109);
   U13119 : BUF_X1 port map( A => n16876, Z => n21666);
   U13120 : INV_X1 port map( A => n18494, ZN => n20895);
   U13121 : INV_X1 port map( A => n18429, ZN => n21168);
   U13122 : INV_X1 port map( A => n16920, ZN => n21452);
   U13123 : INV_X1 port map( A => n16846, ZN => n21725);
   U13124 : INV_X1 port map( A => n18499, ZN => n20850);
   U13125 : INV_X1 port map( A => n18444, ZN => n21236);
   U13126 : INV_X1 port map( A => n18440, ZN => n21184);
   U13127 : INV_X1 port map( A => n18493, ZN => n20887);
   U13128 : INV_X1 port map( A => n18434, ZN => n21134);
   U13129 : INV_X1 port map( A => n18440, ZN => n21185);
   U13130 : INV_X1 port map( A => n18499, ZN => n20851);
   U13131 : INV_X1 port map( A => n16926, ZN => n21407);
   U13132 : INV_X1 port map( A => n16862, ZN => n21793);
   U13133 : INV_X1 port map( A => n16858, ZN => n21741);
   U13134 : INV_X1 port map( A => n16919, ZN => n21444);
   U13135 : INV_X1 port map( A => n16852, ZN => n21691);
   U13136 : INV_X1 port map( A => n16858, ZN => n21742);
   U13137 : INV_X1 port map( A => n16926, ZN => n21408);
   U13138 : BUF_X1 port map( A => n21838, Z => n21831);
   U13139 : BUF_X1 port map( A => n21838, Z => n21832);
   U13140 : BUF_X1 port map( A => n21838, Z => n21833);
   U13141 : BUF_X1 port map( A => n21838, Z => n21834);
   U13142 : BUF_X1 port map( A => n21838, Z => n21835);
   U13143 : BUF_X1 port map( A => n21838, Z => n21836);
   U13144 : BUF_X1 port map( A => n21874, Z => n21867);
   U13145 : BUF_X1 port map( A => n21874, Z => n21868);
   U13146 : BUF_X1 port map( A => n21874, Z => n21869);
   U13147 : BUF_X1 port map( A => n21874, Z => n21870);
   U13148 : BUF_X1 port map( A => n21874, Z => n21871);
   U13149 : BUF_X1 port map( A => n21874, Z => n21872);
   U13150 : BUF_X1 port map( A => n21910, Z => n21903);
   U13151 : BUF_X1 port map( A => n21910, Z => n21904);
   U13152 : BUF_X1 port map( A => n21910, Z => n21905);
   U13153 : BUF_X1 port map( A => n21910, Z => n21906);
   U13154 : BUF_X1 port map( A => n21910, Z => n21907);
   U13155 : BUF_X1 port map( A => n21910, Z => n21908);
   U13156 : BUF_X1 port map( A => n21946, Z => n21939);
   U13157 : BUF_X1 port map( A => n21946, Z => n21940);
   U13158 : BUF_X1 port map( A => n21946, Z => n21941);
   U13159 : BUF_X1 port map( A => n21946, Z => n21942);
   U13160 : BUF_X1 port map( A => n21946, Z => n21943);
   U13161 : BUF_X1 port map( A => n21946, Z => n21944);
   U13162 : BUF_X1 port map( A => n21982, Z => n21975);
   U13163 : BUF_X1 port map( A => n21982, Z => n21976);
   U13164 : BUF_X1 port map( A => n21982, Z => n21977);
   U13165 : BUF_X1 port map( A => n21982, Z => n21978);
   U13166 : BUF_X1 port map( A => n21982, Z => n21979);
   U13167 : BUF_X1 port map( A => n21982, Z => n21980);
   U13168 : BUF_X1 port map( A => n22018, Z => n22011);
   U13169 : BUF_X1 port map( A => n22018, Z => n22012);
   U13170 : BUF_X1 port map( A => n22018, Z => n22013);
   U13171 : BUF_X1 port map( A => n22018, Z => n22014);
   U13172 : BUF_X1 port map( A => n22018, Z => n22015);
   U13173 : BUF_X1 port map( A => n22018, Z => n22016);
   U13174 : BUF_X1 port map( A => n22054, Z => n22047);
   U13175 : BUF_X1 port map( A => n22054, Z => n22048);
   U13176 : BUF_X1 port map( A => n22054, Z => n22049);
   U13177 : BUF_X1 port map( A => n22054, Z => n22050);
   U13178 : BUF_X1 port map( A => n22054, Z => n22051);
   U13179 : BUF_X1 port map( A => n22054, Z => n22052);
   U13180 : BUF_X1 port map( A => n22090, Z => n22083);
   U13181 : BUF_X1 port map( A => n22090, Z => n22084);
   U13182 : BUF_X1 port map( A => n22090, Z => n22085);
   U13183 : BUF_X1 port map( A => n22090, Z => n22086);
   U13184 : BUF_X1 port map( A => n22090, Z => n22087);
   U13185 : BUF_X1 port map( A => n22090, Z => n22088);
   U13186 : BUF_X1 port map( A => n22126, Z => n22119);
   U13187 : BUF_X1 port map( A => n22126, Z => n22120);
   U13188 : BUF_X1 port map( A => n22126, Z => n22121);
   U13189 : BUF_X1 port map( A => n22126, Z => n22122);
   U13190 : BUF_X1 port map( A => n22126, Z => n22123);
   U13191 : BUF_X1 port map( A => n22126, Z => n22124);
   U13192 : BUF_X1 port map( A => n22162, Z => n22155);
   U13193 : BUF_X1 port map( A => n22162, Z => n22156);
   U13194 : BUF_X1 port map( A => n22162, Z => n22157);
   U13195 : BUF_X1 port map( A => n22162, Z => n22158);
   U13196 : BUF_X1 port map( A => n22162, Z => n22159);
   U13197 : BUF_X1 port map( A => n22162, Z => n22160);
   U13198 : BUF_X1 port map( A => n22198, Z => n22191);
   U13199 : BUF_X1 port map( A => n22198, Z => n22192);
   U13200 : BUF_X1 port map( A => n22198, Z => n22193);
   U13201 : BUF_X1 port map( A => n22198, Z => n22194);
   U13202 : BUF_X1 port map( A => n22198, Z => n22195);
   U13203 : BUF_X1 port map( A => n22198, Z => n22196);
   U13204 : BUF_X1 port map( A => n22234, Z => n22227);
   U13205 : BUF_X1 port map( A => n22234, Z => n22228);
   U13206 : BUF_X1 port map( A => n22234, Z => n22229);
   U13207 : BUF_X1 port map( A => n22234, Z => n22230);
   U13208 : BUF_X1 port map( A => n22234, Z => n22231);
   U13209 : BUF_X1 port map( A => n22234, Z => n22232);
   U13210 : BUF_X1 port map( A => n22270, Z => n22263);
   U13211 : BUF_X1 port map( A => n22270, Z => n22264);
   U13212 : BUF_X1 port map( A => n22270, Z => n22265);
   U13213 : BUF_X1 port map( A => n22270, Z => n22266);
   U13214 : BUF_X1 port map( A => n22270, Z => n22267);
   U13215 : BUF_X1 port map( A => n22270, Z => n22268);
   U13216 : BUF_X1 port map( A => n22306, Z => n22299);
   U13217 : BUF_X1 port map( A => n22306, Z => n22300);
   U13218 : BUF_X1 port map( A => n22306, Z => n22301);
   U13219 : BUF_X1 port map( A => n22306, Z => n22302);
   U13220 : BUF_X1 port map( A => n22306, Z => n22303);
   U13221 : BUF_X1 port map( A => n22306, Z => n22304);
   U13222 : BUF_X1 port map( A => n22342, Z => n22335);
   U13223 : BUF_X1 port map( A => n22342, Z => n22336);
   U13224 : BUF_X1 port map( A => n22342, Z => n22337);
   U13225 : BUF_X1 port map( A => n22342, Z => n22338);
   U13226 : BUF_X1 port map( A => n22342, Z => n22339);
   U13227 : BUF_X1 port map( A => n22342, Z => n22340);
   U13228 : BUF_X1 port map( A => n22575, Z => n22568);
   U13229 : BUF_X1 port map( A => n22575, Z => n22569);
   U13230 : BUF_X1 port map( A => n22575, Z => n22570);
   U13231 : BUF_X1 port map( A => n22575, Z => n22571);
   U13232 : BUF_X1 port map( A => n22575, Z => n22572);
   U13233 : BUF_X1 port map( A => n22575, Z => n22573);
   U13234 : BUF_X1 port map( A => n22575, Z => n22574);
   U13235 : BUF_X1 port map( A => n21838, Z => n21837);
   U13236 : BUF_X1 port map( A => n21874, Z => n21873);
   U13237 : BUF_X1 port map( A => n21910, Z => n21909);
   U13238 : BUF_X1 port map( A => n21946, Z => n21945);
   U13239 : BUF_X1 port map( A => n21982, Z => n21981);
   U13240 : BUF_X1 port map( A => n22018, Z => n22017);
   U13241 : BUF_X1 port map( A => n22054, Z => n22053);
   U13242 : BUF_X1 port map( A => n22090, Z => n22089);
   U13243 : BUF_X1 port map( A => n22126, Z => n22125);
   U13244 : BUF_X1 port map( A => n22162, Z => n22161);
   U13245 : BUF_X1 port map( A => n22198, Z => n22197);
   U13246 : BUF_X1 port map( A => n22234, Z => n22233);
   U13247 : BUF_X1 port map( A => n22270, Z => n22269);
   U13248 : BUF_X1 port map( A => n22306, Z => n22305);
   U13249 : BUF_X1 port map( A => n22342, Z => n22341);
   U13250 : BUF_X1 port map( A => n21811, Z => n21810);
   U13251 : BUF_X1 port map( A => n21807, Z => n21808);
   U13252 : BUF_X1 port map( A => n21811, Z => n21807);
   U13253 : BUF_X1 port map( A => n21811, Z => n21806);
   U13254 : BUF_X1 port map( A => n21811, Z => n21805);
   U13255 : BUF_X1 port map( A => n21811, Z => n21804);
   U13256 : BUF_X1 port map( A => n21811, Z => n21803);
   U13257 : BUF_X1 port map( A => n21811, Z => n21802);
   U13258 : BUF_X1 port map( A => n21806, Z => n21809);
   U13259 : INV_X1 port map( A => n21030, ZN => n19624);
   U13260 : INV_X1 port map( A => n21587, ZN => n18351);
   U13261 : INV_X1 port map( A => n20877, ZN => n19674);
   U13262 : INV_X1 port map( A => n21434, ZN => n18410);
   U13263 : INV_X1 port map( A => n20733, ZN => n19634);
   U13264 : INV_X1 port map( A => n21290, ZN => n18361);
   U13265 : INV_X1 port map( A => n20985, ZN => n19637);
   U13266 : INV_X1 port map( A => n21542, ZN => n18365);
   U13267 : INV_X1 port map( A => n16760, ZN => n21838);
   U13268 : OAI21_X1 port map( B1 => n15152, B2 => n16793, A => n22380, ZN => 
                           n16760);
   U13269 : INV_X1 port map( A => n16655, ZN => n21874);
   U13270 : OAI21_X1 port map( B1 => n15152, B2 => n16688, A => n22380, ZN => 
                           n16655);
   U13271 : INV_X1 port map( A => n16613, ZN => n21910);
   U13272 : OAI21_X1 port map( B1 => n15152, B2 => n16614, A => n22379, ZN => 
                           n16613);
   U13273 : INV_X1 port map( A => n16521, ZN => n21946);
   U13274 : OAI21_X1 port map( B1 => n15152, B2 => n16554, A => n22379, ZN => 
                           n16521);
   U13275 : INV_X1 port map( A => n16384, ZN => n21982);
   U13276 : OAI21_X1 port map( B1 => n15152, B2 => n16417, A => n22379, ZN => 
                           n16384);
   U13277 : INV_X1 port map( A => n16343, ZN => n22018);
   U13278 : OAI21_X1 port map( B1 => n15152, B2 => n16344, A => n22378, ZN => 
                           n16343);
   U13279 : INV_X1 port map( A => n16206, ZN => n22054);
   U13280 : OAI21_X1 port map( B1 => n15152, B2 => n16239, A => n22378, ZN => 
                           n16206);
   U13281 : INV_X1 port map( A => n16100, ZN => n22090);
   U13282 : OAI21_X1 port map( B1 => n15152, B2 => n16133, A => n22378, ZN => 
                           n16100);
   U13283 : INV_X1 port map( A => n15963, ZN => n22126);
   U13284 : OAI21_X1 port map( B1 => n15152, B2 => n15996, A => n22377, ZN => 
                           n15963);
   U13285 : INV_X1 port map( A => n15890, ZN => n22162);
   U13286 : OAI21_X1 port map( B1 => n15152, B2 => n15891, A => n22377, ZN => 
                           n15890);
   U13287 : INV_X1 port map( A => n15753, ZN => n22198);
   U13288 : OAI21_X1 port map( B1 => n15152, B2 => n15786, A => n22377, ZN => 
                           n15753);
   U13289 : INV_X1 port map( A => n15647, ZN => n22234);
   U13290 : OAI21_X1 port map( B1 => n15152, B2 => n15680, A => n22377, ZN => 
                           n15647);
   U13291 : INV_X1 port map( A => n15506, ZN => n22270);
   U13292 : OAI21_X1 port map( B1 => n15152, B2 => n15539, A => n22376, ZN => 
                           n15506);
   U13293 : INV_X1 port map( A => n15368, ZN => n22306);
   U13294 : OAI21_X1 port map( B1 => n15152, B2 => n15401, A => n22376, ZN => 
                           n15368);
   U13295 : INV_X1 port map( A => n15230, ZN => n22342);
   U13296 : OAI21_X1 port map( B1 => n15152, B2 => n15263, A => n22376, ZN => 
                           n15230);
   U13297 : INV_X1 port map( A => n15119, ZN => n22575);
   U13298 : OAI21_X1 port map( B1 => n15151, B2 => n15152, A => n22375, ZN => 
                           n15119);
   U13299 : NAND2_X1 port map( A1 => n19623, A2 => n19634, ZN => n18429);
   U13300 : NAND2_X1 port map( A1 => n18350, A2 => n18361, ZN => n16846);
   U13301 : NAND2_X1 port map( A1 => n19623, A2 => n19673, ZN => n18494);
   U13302 : NAND2_X1 port map( A1 => n18350, A2 => n18409, ZN => n16920);
   U13303 : NAND2_X1 port map( A1 => n19623, A2 => n19674, ZN => n18493);
   U13304 : NAND2_X1 port map( A1 => n19623, A2 => n19624, ZN => n18444);
   U13305 : NAND2_X1 port map( A1 => n18350, A2 => n18410, ZN => n16919);
   U13306 : NAND2_X1 port map( A1 => n18350, A2 => n18351, ZN => n16862);
   U13307 : NAND2_X1 port map( A1 => n19623, A2 => n20782, ZN => n18499);
   U13308 : NAND2_X1 port map( A1 => n19623, A2 => n20909, ZN => n18434);
   U13309 : NAND2_X1 port map( A1 => n19623, A2 => n21069, ZN => n18440);
   U13310 : NAND2_X1 port map( A1 => n18350, A2 => n21339, ZN => n16926);
   U13311 : NAND2_X1 port map( A1 => n18350, A2 => n21466, ZN => n16852);
   U13312 : NAND2_X1 port map( A1 => n18350, A2 => n21626, ZN => n16858);
   U13313 : NAND2_X1 port map( A1 => n19623, A2 => n20972, ZN => n18457);
   U13314 : NAND2_X1 port map( A1 => n18350, A2 => n21529, ZN => n16876);
   U13315 : BUF_X1 port map( A => n22371, Z => n22378);
   U13316 : BUF_X1 port map( A => n22371, Z => n22377);
   U13317 : BUF_X1 port map( A => n22371, Z => n22376);
   U13318 : BUF_X1 port map( A => n22372, Z => n22379);
   U13319 : BUF_X1 port map( A => n22370, Z => n22373);
   U13320 : BUF_X1 port map( A => n22370, Z => n22374);
   U13321 : BUF_X1 port map( A => n22370, Z => n22375);
   U13322 : BUF_X1 port map( A => n18473, Z => n20733);
   U13323 : BUF_X1 port map( A => n16894, Z => n21290);
   U13324 : BUF_X1 port map( A => n18478, Z => n20877);
   U13325 : BUF_X1 port map( A => n16899, Z => n21434);
   U13326 : BUF_X1 port map( A => n18473, Z => n20729);
   U13327 : BUF_X1 port map( A => n16894, Z => n21286);
   U13328 : BUF_X1 port map( A => n18478, Z => n20873);
   U13329 : BUF_X1 port map( A => n18473, Z => n20731);
   U13330 : BUF_X1 port map( A => n18478, Z => n20875);
   U13331 : BUF_X1 port map( A => n18473, Z => n20730);
   U13332 : BUF_X1 port map( A => n18478, Z => n20874);
   U13333 : BUF_X1 port map( A => n18473, Z => n20732);
   U13334 : BUF_X1 port map( A => n18478, Z => n20876);
   U13335 : BUF_X1 port map( A => n16899, Z => n21430);
   U13336 : BUF_X1 port map( A => n16894, Z => n21288);
   U13337 : BUF_X1 port map( A => n16899, Z => n21432);
   U13338 : BUF_X1 port map( A => n16894, Z => n21287);
   U13339 : BUF_X1 port map( A => n16899, Z => n21431);
   U13340 : BUF_X1 port map( A => n16894, Z => n21289);
   U13341 : BUF_X1 port map( A => n16899, Z => n21433);
   U13342 : BUF_X1 port map( A => n18462, Z => n21030);
   U13343 : BUF_X1 port map( A => n16881, Z => n21587);
   U13344 : BUF_X1 port map( A => n18467, Z => n20985);
   U13345 : BUF_X1 port map( A => n16887, Z => n21542);
   U13346 : BUF_X1 port map( A => n18451, Z => n20978);
   U13347 : BUF_X1 port map( A => n18437, Z => n21209);
   U13348 : BUF_X1 port map( A => n18451, Z => n20979);
   U13349 : BUF_X1 port map( A => n16869, Z => n21535);
   U13350 : BUF_X1 port map( A => n16855, Z => n21766);
   U13351 : BUF_X1 port map( A => n16869, Z => n21536);
   U13352 : BUF_X1 port map( A => n18462, Z => n21026);
   U13353 : BUF_X1 port map( A => n18462, Z => n21028);
   U13354 : BUF_X1 port map( A => n18462, Z => n21027);
   U13355 : BUF_X1 port map( A => n18467, Z => n20984);
   U13356 : BUF_X1 port map( A => n18462, Z => n21029);
   U13357 : BUF_X1 port map( A => n16881, Z => n21583);
   U13358 : BUF_X1 port map( A => n16881, Z => n21585);
   U13359 : BUF_X1 port map( A => n16881, Z => n21584);
   U13360 : BUF_X1 port map( A => n16887, Z => n21541);
   U13361 : BUF_X1 port map( A => n16881, Z => n21586);
   U13362 : BUF_X1 port map( A => n18467, Z => n20981);
   U13363 : BUF_X1 port map( A => n18467, Z => n20983);
   U13364 : BUF_X1 port map( A => n18467, Z => n20982);
   U13365 : BUF_X1 port map( A => n16887, Z => n21538);
   U13366 : BUF_X1 port map( A => n16887, Z => n21540);
   U13367 : BUF_X1 port map( A => n16887, Z => n21539);
   U13368 : BUF_X1 port map( A => n18437, Z => n21210);
   U13369 : BUF_X1 port map( A => n16855, Z => n21767);
   U13370 : BUF_X1 port map( A => n18473, Z => n20734);
   U13371 : BUF_X1 port map( A => n16894, Z => n21291);
   U13372 : BUF_X1 port map( A => n18478, Z => n20878);
   U13373 : BUF_X1 port map( A => n16899, Z => n21435);
   U13374 : BUF_X1 port map( A => n18451, Z => n20980);
   U13375 : BUF_X1 port map( A => n18437, Z => n21211);
   U13376 : BUF_X1 port map( A => n16869, Z => n21537);
   U13377 : BUF_X1 port map( A => n16855, Z => n21768);
   U13378 : BUF_X1 port map( A => n18462, Z => n21031);
   U13379 : BUF_X1 port map( A => n16881, Z => n21588);
   U13380 : BUF_X1 port map( A => n18467, Z => n20986);
   U13381 : BUF_X1 port map( A => n16887, Z => n21543);
   U13382 : BUF_X1 port map( A => n22372, Z => n22380);
   U13383 : AND2_X1 port map( A1 => n19623, A2 => n19633, ZN => n18495);
   U13384 : AND2_X1 port map( A1 => n19623, A2 => n20716, ZN => n18500);
   U13385 : AND2_X1 port map( A1 => n19623, A2 => n19635, ZN => n18426);
   U13386 : AND2_X1 port map( A1 => n19623, A2 => n21023, ZN => n18425);
   U13387 : AND2_X1 port map( A1 => n19623, A2 => n19637, ZN => n18432);
   U13388 : AND2_X1 port map( A1 => n19623, A2 => n19626, ZN => n18442);
   U13389 : AND2_X1 port map( A1 => n19623, A2 => n21101, ZN => n18436);
   U13390 : AND2_X1 port map( A1 => n18350, A2 => n18360, ZN => n16921);
   U13391 : AND2_X1 port map( A1 => n18350, A2 => n21273, ZN => n16927);
   U13392 : AND2_X1 port map( A1 => n18350, A2 => n18362, ZN => n16843);
   U13393 : AND2_X1 port map( A1 => n18350, A2 => n21580, ZN => n16842);
   U13394 : AND2_X1 port map( A1 => n18350, A2 => n18365, ZN => n16849);
   U13395 : AND2_X1 port map( A1 => n18350, A2 => n18353, ZN => n16860);
   U13396 : AND2_X1 port map( A1 => n18350, A2 => n21658, ZN => n16854);
   U13397 : AND2_X1 port map( A1 => n19623, A2 => n20835, ZN => n18496);
   U13398 : AND2_X1 port map( A1 => n18350, A2 => n21392, ZN => n16922);
   U13399 : BUF_X1 port map( A => n21820, Z => n21813);
   U13400 : BUF_X1 port map( A => n21820, Z => n21814);
   U13401 : BUF_X1 port map( A => n21820, Z => n21815);
   U13402 : BUF_X1 port map( A => n21820, Z => n21816);
   U13403 : BUF_X1 port map( A => n21820, Z => n21817);
   U13404 : BUF_X1 port map( A => n21820, Z => n21818);
   U13405 : BUF_X1 port map( A => n21829, Z => n21822);
   U13406 : BUF_X1 port map( A => n21829, Z => n21823);
   U13407 : BUF_X1 port map( A => n21829, Z => n21824);
   U13408 : BUF_X1 port map( A => n21829, Z => n21825);
   U13409 : BUF_X1 port map( A => n21829, Z => n21826);
   U13410 : BUF_X1 port map( A => n21829, Z => n21827);
   U13411 : BUF_X1 port map( A => n21847, Z => n21840);
   U13412 : BUF_X1 port map( A => n21847, Z => n21841);
   U13413 : BUF_X1 port map( A => n21847, Z => n21842);
   U13414 : BUF_X1 port map( A => n21847, Z => n21843);
   U13415 : BUF_X1 port map( A => n21847, Z => n21844);
   U13416 : BUF_X1 port map( A => n21847, Z => n21845);
   U13417 : BUF_X1 port map( A => n21856, Z => n21849);
   U13418 : BUF_X1 port map( A => n21856, Z => n21850);
   U13419 : BUF_X1 port map( A => n21856, Z => n21851);
   U13420 : BUF_X1 port map( A => n21856, Z => n21852);
   U13421 : BUF_X1 port map( A => n21856, Z => n21853);
   U13422 : BUF_X1 port map( A => n21856, Z => n21854);
   U13423 : BUF_X1 port map( A => n21865, Z => n21858);
   U13424 : BUF_X1 port map( A => n21865, Z => n21859);
   U13425 : BUF_X1 port map( A => n21865, Z => n21860);
   U13426 : BUF_X1 port map( A => n21865, Z => n21861);
   U13427 : BUF_X1 port map( A => n21865, Z => n21862);
   U13428 : BUF_X1 port map( A => n21865, Z => n21863);
   U13429 : BUF_X1 port map( A => n21883, Z => n21876);
   U13430 : BUF_X1 port map( A => n21883, Z => n21877);
   U13431 : BUF_X1 port map( A => n21883, Z => n21878);
   U13432 : BUF_X1 port map( A => n21883, Z => n21879);
   U13433 : BUF_X1 port map( A => n21883, Z => n21880);
   U13434 : BUF_X1 port map( A => n21883, Z => n21881);
   U13435 : BUF_X1 port map( A => n21892, Z => n21885);
   U13436 : BUF_X1 port map( A => n21892, Z => n21886);
   U13437 : BUF_X1 port map( A => n21892, Z => n21887);
   U13438 : BUF_X1 port map( A => n21892, Z => n21888);
   U13439 : BUF_X1 port map( A => n21892, Z => n21889);
   U13440 : BUF_X1 port map( A => n21892, Z => n21890);
   U13441 : BUF_X1 port map( A => n21901, Z => n21894);
   U13442 : BUF_X1 port map( A => n21901, Z => n21895);
   U13443 : BUF_X1 port map( A => n21901, Z => n21896);
   U13444 : BUF_X1 port map( A => n21901, Z => n21897);
   U13445 : BUF_X1 port map( A => n21901, Z => n21898);
   U13446 : BUF_X1 port map( A => n21901, Z => n21899);
   U13447 : BUF_X1 port map( A => n21919, Z => n21912);
   U13448 : BUF_X1 port map( A => n21919, Z => n21913);
   U13449 : BUF_X1 port map( A => n21919, Z => n21914);
   U13450 : BUF_X1 port map( A => n21919, Z => n21915);
   U13451 : BUF_X1 port map( A => n21919, Z => n21916);
   U13452 : BUF_X1 port map( A => n21919, Z => n21917);
   U13453 : BUF_X1 port map( A => n21928, Z => n21921);
   U13454 : BUF_X1 port map( A => n21928, Z => n21922);
   U13455 : BUF_X1 port map( A => n21928, Z => n21923);
   U13456 : BUF_X1 port map( A => n21928, Z => n21924);
   U13457 : BUF_X1 port map( A => n21928, Z => n21925);
   U13458 : BUF_X1 port map( A => n21928, Z => n21926);
   U13459 : BUF_X1 port map( A => n21937, Z => n21930);
   U13460 : BUF_X1 port map( A => n21937, Z => n21931);
   U13461 : BUF_X1 port map( A => n21937, Z => n21932);
   U13462 : BUF_X1 port map( A => n21937, Z => n21933);
   U13463 : BUF_X1 port map( A => n21937, Z => n21934);
   U13464 : BUF_X1 port map( A => n21937, Z => n21935);
   U13465 : BUF_X1 port map( A => n21955, Z => n21948);
   U13466 : BUF_X1 port map( A => n21955, Z => n21949);
   U13467 : BUF_X1 port map( A => n21955, Z => n21950);
   U13468 : BUF_X1 port map( A => n21955, Z => n21951);
   U13469 : BUF_X1 port map( A => n21955, Z => n21952);
   U13470 : BUF_X1 port map( A => n21955, Z => n21953);
   U13471 : BUF_X1 port map( A => n21964, Z => n21957);
   U13472 : BUF_X1 port map( A => n21964, Z => n21958);
   U13473 : BUF_X1 port map( A => n21964, Z => n21959);
   U13474 : BUF_X1 port map( A => n21964, Z => n21960);
   U13475 : BUF_X1 port map( A => n21964, Z => n21961);
   U13476 : BUF_X1 port map( A => n21964, Z => n21962);
   U13477 : BUF_X1 port map( A => n21973, Z => n21966);
   U13478 : BUF_X1 port map( A => n21973, Z => n21967);
   U13479 : BUF_X1 port map( A => n21973, Z => n21968);
   U13480 : BUF_X1 port map( A => n21973, Z => n21969);
   U13481 : BUF_X1 port map( A => n21973, Z => n21970);
   U13482 : BUF_X1 port map( A => n21973, Z => n21971);
   U13483 : BUF_X1 port map( A => n21991, Z => n21984);
   U13484 : BUF_X1 port map( A => n21991, Z => n21985);
   U13485 : BUF_X1 port map( A => n21991, Z => n21986);
   U13486 : BUF_X1 port map( A => n21991, Z => n21987);
   U13487 : BUF_X1 port map( A => n21991, Z => n21988);
   U13488 : BUF_X1 port map( A => n21991, Z => n21989);
   U13489 : BUF_X1 port map( A => n22000, Z => n21993);
   U13490 : BUF_X1 port map( A => n22000, Z => n21994);
   U13491 : BUF_X1 port map( A => n22000, Z => n21995);
   U13492 : BUF_X1 port map( A => n22000, Z => n21996);
   U13493 : BUF_X1 port map( A => n22000, Z => n21997);
   U13494 : BUF_X1 port map( A => n22000, Z => n21998);
   U13495 : BUF_X1 port map( A => n22009, Z => n22002);
   U13496 : BUF_X1 port map( A => n22009, Z => n22003);
   U13497 : BUF_X1 port map( A => n22009, Z => n22004);
   U13498 : BUF_X1 port map( A => n22009, Z => n22005);
   U13499 : BUF_X1 port map( A => n22009, Z => n22006);
   U13500 : BUF_X1 port map( A => n22009, Z => n22007);
   U13501 : BUF_X1 port map( A => n22027, Z => n22020);
   U13502 : BUF_X1 port map( A => n22027, Z => n22021);
   U13503 : BUF_X1 port map( A => n22027, Z => n22022);
   U13504 : BUF_X1 port map( A => n22027, Z => n22023);
   U13505 : BUF_X1 port map( A => n22027, Z => n22024);
   U13506 : BUF_X1 port map( A => n22027, Z => n22025);
   U13507 : BUF_X1 port map( A => n22036, Z => n22029);
   U13508 : BUF_X1 port map( A => n22036, Z => n22030);
   U13509 : BUF_X1 port map( A => n22036, Z => n22031);
   U13510 : BUF_X1 port map( A => n22036, Z => n22032);
   U13511 : BUF_X1 port map( A => n22036, Z => n22033);
   U13512 : BUF_X1 port map( A => n22036, Z => n22034);
   U13513 : BUF_X1 port map( A => n22045, Z => n22038);
   U13514 : BUF_X1 port map( A => n22045, Z => n22039);
   U13515 : BUF_X1 port map( A => n22045, Z => n22040);
   U13516 : BUF_X1 port map( A => n22045, Z => n22041);
   U13517 : BUF_X1 port map( A => n22045, Z => n22042);
   U13518 : BUF_X1 port map( A => n22045, Z => n22043);
   U13519 : BUF_X1 port map( A => n22063, Z => n22056);
   U13520 : BUF_X1 port map( A => n22063, Z => n22057);
   U13521 : BUF_X1 port map( A => n22063, Z => n22058);
   U13522 : BUF_X1 port map( A => n22063, Z => n22059);
   U13523 : BUF_X1 port map( A => n22063, Z => n22060);
   U13524 : BUF_X1 port map( A => n22063, Z => n22061);
   U13525 : BUF_X1 port map( A => n22072, Z => n22065);
   U13526 : BUF_X1 port map( A => n22072, Z => n22066);
   U13527 : BUF_X1 port map( A => n22072, Z => n22067);
   U13528 : BUF_X1 port map( A => n22072, Z => n22068);
   U13529 : BUF_X1 port map( A => n22072, Z => n22069);
   U13530 : BUF_X1 port map( A => n22072, Z => n22070);
   U13531 : BUF_X1 port map( A => n22081, Z => n22074);
   U13532 : BUF_X1 port map( A => n22081, Z => n22075);
   U13533 : BUF_X1 port map( A => n22081, Z => n22076);
   U13534 : BUF_X1 port map( A => n22081, Z => n22077);
   U13535 : BUF_X1 port map( A => n22081, Z => n22078);
   U13536 : BUF_X1 port map( A => n22081, Z => n22079);
   U13537 : BUF_X1 port map( A => n22099, Z => n22092);
   U13538 : BUF_X1 port map( A => n22099, Z => n22093);
   U13539 : BUF_X1 port map( A => n22099, Z => n22094);
   U13540 : BUF_X1 port map( A => n22099, Z => n22095);
   U13541 : BUF_X1 port map( A => n22099, Z => n22096);
   U13542 : BUF_X1 port map( A => n22099, Z => n22097);
   U13543 : BUF_X1 port map( A => n22108, Z => n22101);
   U13544 : BUF_X1 port map( A => n22108, Z => n22102);
   U13545 : BUF_X1 port map( A => n22108, Z => n22103);
   U13546 : BUF_X1 port map( A => n22108, Z => n22104);
   U13547 : BUF_X1 port map( A => n22108, Z => n22105);
   U13548 : BUF_X1 port map( A => n22108, Z => n22106);
   U13549 : BUF_X1 port map( A => n22117, Z => n22110);
   U13550 : BUF_X1 port map( A => n22117, Z => n22111);
   U13551 : BUF_X1 port map( A => n22117, Z => n22112);
   U13552 : BUF_X1 port map( A => n22117, Z => n22113);
   U13553 : BUF_X1 port map( A => n22117, Z => n22114);
   U13554 : BUF_X1 port map( A => n22117, Z => n22115);
   U13555 : BUF_X1 port map( A => n22135, Z => n22128);
   U13556 : BUF_X1 port map( A => n22135, Z => n22129);
   U13557 : BUF_X1 port map( A => n22135, Z => n22130);
   U13558 : BUF_X1 port map( A => n22135, Z => n22131);
   U13559 : BUF_X1 port map( A => n22135, Z => n22132);
   U13560 : BUF_X1 port map( A => n22135, Z => n22133);
   U13561 : BUF_X1 port map( A => n22144, Z => n22137);
   U13562 : BUF_X1 port map( A => n22144, Z => n22138);
   U13563 : BUF_X1 port map( A => n22144, Z => n22139);
   U13564 : BUF_X1 port map( A => n22144, Z => n22140);
   U13565 : BUF_X1 port map( A => n22144, Z => n22141);
   U13566 : BUF_X1 port map( A => n22144, Z => n22142);
   U13567 : BUF_X1 port map( A => n22153, Z => n22146);
   U13568 : BUF_X1 port map( A => n22153, Z => n22147);
   U13569 : BUF_X1 port map( A => n22153, Z => n22148);
   U13570 : BUF_X1 port map( A => n22153, Z => n22149);
   U13571 : BUF_X1 port map( A => n22153, Z => n22150);
   U13572 : BUF_X1 port map( A => n22153, Z => n22151);
   U13573 : BUF_X1 port map( A => n22171, Z => n22164);
   U13574 : BUF_X1 port map( A => n22171, Z => n22165);
   U13575 : BUF_X1 port map( A => n22171, Z => n22166);
   U13576 : BUF_X1 port map( A => n22171, Z => n22167);
   U13577 : BUF_X1 port map( A => n22171, Z => n22168);
   U13578 : BUF_X1 port map( A => n22171, Z => n22169);
   U13579 : BUF_X1 port map( A => n22180, Z => n22173);
   U13580 : BUF_X1 port map( A => n22180, Z => n22174);
   U13581 : BUF_X1 port map( A => n22180, Z => n22175);
   U13582 : BUF_X1 port map( A => n22180, Z => n22176);
   U13583 : BUF_X1 port map( A => n22180, Z => n22177);
   U13584 : BUF_X1 port map( A => n22180, Z => n22178);
   U13585 : BUF_X1 port map( A => n22189, Z => n22182);
   U13586 : BUF_X1 port map( A => n22189, Z => n22183);
   U13587 : BUF_X1 port map( A => n22189, Z => n22184);
   U13588 : BUF_X1 port map( A => n22189, Z => n22185);
   U13589 : BUF_X1 port map( A => n22189, Z => n22186);
   U13590 : BUF_X1 port map( A => n22189, Z => n22187);
   U13591 : BUF_X1 port map( A => n22207, Z => n22200);
   U13592 : BUF_X1 port map( A => n22207, Z => n22201);
   U13593 : BUF_X1 port map( A => n22207, Z => n22202);
   U13594 : BUF_X1 port map( A => n22207, Z => n22203);
   U13595 : BUF_X1 port map( A => n22207, Z => n22204);
   U13596 : BUF_X1 port map( A => n22207, Z => n22205);
   U13597 : BUF_X1 port map( A => n22216, Z => n22209);
   U13598 : BUF_X1 port map( A => n22216, Z => n22210);
   U13599 : BUF_X1 port map( A => n22216, Z => n22211);
   U13600 : BUF_X1 port map( A => n22216, Z => n22212);
   U13601 : BUF_X1 port map( A => n22216, Z => n22213);
   U13602 : BUF_X1 port map( A => n22216, Z => n22214);
   U13603 : BUF_X1 port map( A => n22225, Z => n22218);
   U13604 : BUF_X1 port map( A => n22225, Z => n22219);
   U13605 : BUF_X1 port map( A => n22225, Z => n22220);
   U13606 : BUF_X1 port map( A => n22225, Z => n22221);
   U13607 : BUF_X1 port map( A => n22225, Z => n22222);
   U13608 : BUF_X1 port map( A => n22225, Z => n22223);
   U13609 : BUF_X1 port map( A => n22243, Z => n22236);
   U13610 : BUF_X1 port map( A => n22243, Z => n22237);
   U13611 : BUF_X1 port map( A => n22243, Z => n22238);
   U13612 : BUF_X1 port map( A => n22243, Z => n22239);
   U13613 : BUF_X1 port map( A => n22243, Z => n22240);
   U13614 : BUF_X1 port map( A => n22243, Z => n22241);
   U13615 : BUF_X1 port map( A => n22252, Z => n22245);
   U13616 : BUF_X1 port map( A => n22252, Z => n22246);
   U13617 : BUF_X1 port map( A => n22252, Z => n22247);
   U13618 : BUF_X1 port map( A => n22252, Z => n22248);
   U13619 : BUF_X1 port map( A => n22252, Z => n22249);
   U13620 : BUF_X1 port map( A => n22252, Z => n22250);
   U13621 : BUF_X1 port map( A => n22261, Z => n22254);
   U13622 : BUF_X1 port map( A => n22261, Z => n22255);
   U13623 : BUF_X1 port map( A => n22261, Z => n22256);
   U13624 : BUF_X1 port map( A => n22261, Z => n22257);
   U13625 : BUF_X1 port map( A => n22261, Z => n22258);
   U13626 : BUF_X1 port map( A => n22261, Z => n22259);
   U13627 : BUF_X1 port map( A => n22279, Z => n22272);
   U13628 : BUF_X1 port map( A => n22279, Z => n22273);
   U13629 : BUF_X1 port map( A => n22279, Z => n22274);
   U13630 : BUF_X1 port map( A => n22279, Z => n22275);
   U13631 : BUF_X1 port map( A => n22279, Z => n22276);
   U13632 : BUF_X1 port map( A => n22279, Z => n22277);
   U13633 : BUF_X1 port map( A => n22288, Z => n22281);
   U13634 : BUF_X1 port map( A => n22288, Z => n22282);
   U13635 : BUF_X1 port map( A => n22288, Z => n22283);
   U13636 : BUF_X1 port map( A => n22288, Z => n22284);
   U13637 : BUF_X1 port map( A => n22288, Z => n22285);
   U13638 : BUF_X1 port map( A => n22288, Z => n22286);
   U13639 : BUF_X1 port map( A => n22297, Z => n22290);
   U13640 : BUF_X1 port map( A => n22297, Z => n22291);
   U13641 : BUF_X1 port map( A => n22297, Z => n22292);
   U13642 : BUF_X1 port map( A => n22297, Z => n22293);
   U13643 : BUF_X1 port map( A => n22297, Z => n22294);
   U13644 : BUF_X1 port map( A => n22297, Z => n22295);
   U13645 : BUF_X1 port map( A => n22315, Z => n22308);
   U13646 : BUF_X1 port map( A => n22315, Z => n22309);
   U13647 : BUF_X1 port map( A => n22315, Z => n22310);
   U13648 : BUF_X1 port map( A => n22315, Z => n22311);
   U13649 : BUF_X1 port map( A => n22315, Z => n22312);
   U13650 : BUF_X1 port map( A => n22315, Z => n22313);
   U13651 : BUF_X1 port map( A => n22324, Z => n22317);
   U13652 : BUF_X1 port map( A => n22324, Z => n22318);
   U13653 : BUF_X1 port map( A => n22324, Z => n22319);
   U13654 : BUF_X1 port map( A => n22324, Z => n22320);
   U13655 : BUF_X1 port map( A => n22324, Z => n22321);
   U13656 : BUF_X1 port map( A => n22324, Z => n22322);
   U13657 : BUF_X1 port map( A => n22333, Z => n22326);
   U13658 : BUF_X1 port map( A => n22333, Z => n22327);
   U13659 : BUF_X1 port map( A => n22333, Z => n22328);
   U13660 : BUF_X1 port map( A => n22333, Z => n22329);
   U13661 : BUF_X1 port map( A => n22333, Z => n22330);
   U13662 : BUF_X1 port map( A => n22333, Z => n22331);
   U13663 : BUF_X1 port map( A => n22351, Z => n22344);
   U13664 : BUF_X1 port map( A => n22351, Z => n22345);
   U13665 : BUF_X1 port map( A => n22351, Z => n22346);
   U13666 : BUF_X1 port map( A => n22351, Z => n22347);
   U13667 : BUF_X1 port map( A => n22351, Z => n22348);
   U13668 : BUF_X1 port map( A => n22351, Z => n22349);
   U13669 : BUF_X1 port map( A => n22360, Z => n22353);
   U13670 : BUF_X1 port map( A => n22360, Z => n22354);
   U13671 : BUF_X1 port map( A => n22360, Z => n22355);
   U13672 : BUF_X1 port map( A => n22360, Z => n22356);
   U13673 : BUF_X1 port map( A => n22360, Z => n22357);
   U13674 : BUF_X1 port map( A => n22360, Z => n22358);
   U13675 : BUF_X1 port map( A => n22369, Z => n22362);
   U13676 : BUF_X1 port map( A => n22369, Z => n22363);
   U13677 : BUF_X1 port map( A => n22369, Z => n22364);
   U13678 : BUF_X1 port map( A => n22369, Z => n22365);
   U13679 : BUF_X1 port map( A => n22369, Z => n22366);
   U13680 : BUF_X1 port map( A => n22369, Z => n22367);
   U13681 : INV_X1 port map( A => n18445, ZN => n21228);
   U13682 : INV_X1 port map( A => n18435, ZN => n21126);
   U13683 : INV_X1 port map( A => n16863, ZN => n21785);
   U13684 : INV_X1 port map( A => n16853, ZN => n21683);
   U13685 : INV_X1 port map( A => n18428, ZN => n21176);
   U13686 : INV_X1 port map( A => n16845, ZN => n21733);
   U13687 : INV_X1 port map( A => n18439, ZN => n21193);
   U13688 : INV_X1 port map( A => n18430, ZN => n21159);
   U13689 : INV_X1 port map( A => n18498, ZN => n20842);
   U13690 : INV_X1 port map( A => n18504, ZN => n20784);
   U13691 : INV_X1 port map( A => n18503, ZN => n20743);
   U13692 : INV_X1 port map( A => n18430, ZN => n21160);
   U13693 : INV_X1 port map( A => n16857, ZN => n21750);
   U13694 : INV_X1 port map( A => n16847, ZN => n21716);
   U13695 : INV_X1 port map( A => n16925, ZN => n21399);
   U13696 : INV_X1 port map( A => n16931, ZN => n21341);
   U13697 : INV_X1 port map( A => n16930, ZN => n21300);
   U13698 : INV_X1 port map( A => n16847, ZN => n21717);
   U13699 : BUF_X1 port map( A => n22351, Z => n22350);
   U13700 : BUF_X1 port map( A => n22360, Z => n22359);
   U13701 : BUF_X1 port map( A => n22369, Z => n22368);
   U13702 : BUF_X1 port map( A => n21820, Z => n21819);
   U13703 : BUF_X1 port map( A => n21829, Z => n21828);
   U13704 : BUF_X1 port map( A => n21847, Z => n21846);
   U13705 : BUF_X1 port map( A => n21856, Z => n21855);
   U13706 : BUF_X1 port map( A => n21865, Z => n21864);
   U13707 : BUF_X1 port map( A => n21883, Z => n21882);
   U13708 : BUF_X1 port map( A => n21892, Z => n21891);
   U13709 : BUF_X1 port map( A => n21901, Z => n21900);
   U13710 : BUF_X1 port map( A => n21919, Z => n21918);
   U13711 : BUF_X1 port map( A => n21928, Z => n21927);
   U13712 : BUF_X1 port map( A => n21937, Z => n21936);
   U13713 : BUF_X1 port map( A => n21955, Z => n21954);
   U13714 : BUF_X1 port map( A => n21964, Z => n21963);
   U13715 : BUF_X1 port map( A => n21973, Z => n21972);
   U13716 : BUF_X1 port map( A => n21991, Z => n21990);
   U13717 : BUF_X1 port map( A => n22000, Z => n21999);
   U13718 : BUF_X1 port map( A => n22009, Z => n22008);
   U13719 : BUF_X1 port map( A => n22027, Z => n22026);
   U13720 : BUF_X1 port map( A => n22036, Z => n22035);
   U13721 : BUF_X1 port map( A => n22045, Z => n22044);
   U13722 : BUF_X1 port map( A => n22063, Z => n22062);
   U13723 : BUF_X1 port map( A => n22072, Z => n22071);
   U13724 : BUF_X1 port map( A => n22081, Z => n22080);
   U13725 : BUF_X1 port map( A => n22099, Z => n22098);
   U13726 : BUF_X1 port map( A => n22108, Z => n22107);
   U13727 : BUF_X1 port map( A => n22117, Z => n22116);
   U13728 : BUF_X1 port map( A => n22135, Z => n22134);
   U13729 : BUF_X1 port map( A => n22144, Z => n22143);
   U13730 : BUF_X1 port map( A => n22153, Z => n22152);
   U13731 : BUF_X1 port map( A => n22171, Z => n22170);
   U13732 : BUF_X1 port map( A => n22180, Z => n22179);
   U13733 : BUF_X1 port map( A => n22189, Z => n22188);
   U13734 : BUF_X1 port map( A => n22207, Z => n22206);
   U13735 : BUF_X1 port map( A => n22216, Z => n22215);
   U13736 : BUF_X1 port map( A => n22225, Z => n22224);
   U13737 : BUF_X1 port map( A => n22243, Z => n22242);
   U13738 : BUF_X1 port map( A => n22252, Z => n22251);
   U13739 : BUF_X1 port map( A => n22261, Z => n22260);
   U13740 : BUF_X1 port map( A => n22279, Z => n22278);
   U13741 : BUF_X1 port map( A => n22288, Z => n22287);
   U13742 : BUF_X1 port map( A => n22297, Z => n22296);
   U13743 : BUF_X1 port map( A => n22315, Z => n22314);
   U13744 : BUF_X1 port map( A => n22324, Z => n22323);
   U13745 : BUF_X1 port map( A => n22333, Z => n22332);
   U13746 : INV_X1 port map( A => n20991, ZN => n19635);
   U13747 : INV_X1 port map( A => n21548, ZN => n18362);
   U13748 : INV_X1 port map( A => n20796, ZN => n19633);
   U13749 : INV_X1 port map( A => n21353, ZN => n18360);
   U13750 : INV_X1 port map( A => n20863, ZN => n19673);
   U13751 : INV_X1 port map( A => n21420, ZN => n18409);
   U13752 : INV_X1 port map( A => n21036, ZN => n19626);
   U13753 : INV_X1 port map( A => n21593, ZN => n18353);
   U13754 : INV_X1 port map( A => n16832, ZN => n21811);
   U13755 : INV_X4 port map( A => n19616, ZN => n18417);
   U13756 : INV_X4 port map( A => n18343, ZN => n16834);
   U13757 : NAND2_X1 port map( A1 => n19645, A2 => n19646, ZN => n21105);
   U13758 : NAND2_X1 port map( A1 => n19645, A2 => n19646, ZN => n21106);
   U13759 : NAND2_X1 port map( A1 => n18374, A2 => n18375, ZN => n21662);
   U13760 : NAND2_X1 port map( A1 => n18374, A2 => n18375, ZN => n21663);
   U13761 : NAND2_X1 port map( A1 => n19645, A2 => n19646, ZN => n18456);
   U13762 : NAND2_X1 port map( A1 => n18374, A2 => n18375, ZN => n16875);
   U13763 : NOR3_X1 port map( A1 => n19665, A2 => n19671, A3 => n19666, ZN => 
                           n19677);
   U13764 : NOR3_X1 port map( A1 => n18399, A2 => n18406, A3 => n18400, ZN => 
                           n18414);
   U13765 : NAND2_X1 port map( A1 => n16794, A2 => n16795, ZN => n15152);
   U13766 : INV_X1 port map( A => n16831, ZN => n21820);
   U13767 : OAI21_X1 port map( B1 => n15191, B2 => n16793, A => n22380, ZN => 
                           n16831);
   U13768 : INV_X1 port map( A => n16724, ZN => n21856);
   U13769 : OAI21_X1 port map( B1 => n15191, B2 => n16688, A => n22380, ZN => 
                           n16724);
   U13770 : INV_X1 port map( A => n16618, ZN => n21892);
   U13771 : OAI21_X1 port map( B1 => n15191, B2 => n16614, A => n22380, ZN => 
                           n16618);
   U13772 : INV_X1 port map( A => n16576, ZN => n21928);
   U13773 : OAI21_X1 port map( B1 => n15191, B2 => n16554, A => n22379, ZN => 
                           n16576);
   U13774 : INV_X1 port map( A => n16453, ZN => n21964);
   U13775 : OAI21_X1 port map( B1 => n15191, B2 => n16417, A => n22379, ZN => 
                           n16453);
   U13776 : INV_X1 port map( A => n16348, ZN => n22000);
   U13777 : OAI21_X1 port map( B1 => n15191, B2 => n16344, A => n22379, ZN => 
                           n16348);
   U13778 : INV_X1 port map( A => n16275, ZN => n22036);
   U13779 : OAI21_X1 port map( B1 => n15191, B2 => n16239, A => n22378, ZN => 
                           n16275);
   U13780 : INV_X1 port map( A => n16169, ZN => n22072);
   U13781 : OAI21_X1 port map( B1 => n15191, B2 => n16133, A => n22378, ZN => 
                           n16169);
   U13782 : INV_X1 port map( A => n16032, ZN => n22108);
   U13783 : OAI21_X1 port map( B1 => n15191, B2 => n15996, A => n22378, ZN => 
                           n16032);
   U13784 : INV_X1 port map( A => n15895, ZN => n22144);
   U13785 : OAI21_X1 port map( B1 => n15191, B2 => n15891, A => n22377, ZN => 
                           n15895);
   U13786 : INV_X1 port map( A => n15822, ZN => n22180);
   U13787 : OAI21_X1 port map( B1 => n15191, B2 => n15786, A => n22378, ZN => 
                           n15822);
   U13788 : INV_X1 port map( A => n15716, ZN => n22216);
   U13789 : OAI21_X1 port map( B1 => n15191, B2 => n15680, A => n22377, ZN => 
                           n15716);
   U13790 : INV_X1 port map( A => n15575, ZN => n22252);
   U13791 : OAI21_X1 port map( B1 => n15191, B2 => n15539, A => n22376, ZN => 
                           n15575);
   U13792 : INV_X1 port map( A => n15437, ZN => n22288);
   U13793 : OAI21_X1 port map( B1 => n15191, B2 => n15401, A => n22376, ZN => 
                           n15437);
   U13794 : INV_X1 port map( A => n15299, ZN => n22324);
   U13795 : OAI21_X1 port map( B1 => n15191, B2 => n15263, A => n22376, ZN => 
                           n15299);
   U13796 : INV_X1 port map( A => n15193, ZN => n22351);
   U13797 : OAI21_X1 port map( B1 => n15151, B2 => n15226, A => n22376, ZN => 
                           n15193);
   U13798 : INV_X1 port map( A => n15158, ZN => n22360);
   U13799 : OAI21_X1 port map( B1 => n15151, B2 => n15191, A => n22375, ZN => 
                           n15158);
   U13800 : INV_X1 port map( A => n15155, ZN => n22369);
   U13801 : OAI21_X1 port map( B1 => n15151, B2 => n15156, A => n22375, ZN => 
                           n15155);
   U13802 : NAND2_X1 port map( A1 => n19663, A2 => n19661, ZN => n18462);
   U13803 : NAND2_X1 port map( A1 => n18396, A2 => n18394, ZN => n16881);
   U13804 : NAND2_X1 port map( A1 => n19678, A2 => n19661, ZN => n18473);
   U13805 : NAND2_X1 port map( A1 => n18415, A2 => n18394, ZN => n16894);
   U13806 : NAND2_X1 port map( A1 => n19667, A2 => n19661, ZN => n18467);
   U13807 : NAND2_X1 port map( A1 => n18401, A2 => n18394, ZN => n16887);
   U13808 : NAND2_X1 port map( A1 => n19675, A2 => n19661, ZN => n18478);
   U13809 : NAND2_X1 port map( A1 => n18411, A2 => n18394, ZN => n16899);
   U13810 : OAI22_X1 port map( A1 => n16203, A2 => n18493, B1 => n16341, B2 => 
                           n18494, ZN => n19672);
   U13811 : OAI22_X1 port map( A1 => n16203, A2 => n16919, B1 => n16341, B2 => 
                           n16920, ZN => n18408);
   U13812 : INV_X1 port map( A => n19636, ZN => n19629);
   U13813 : OAI22_X1 port map( A1 => n21128, A2 => n15854, B1 => n21141, B2 => 
                           n16519, ZN => n19636);
   U13814 : INV_X1 port map( A => n18363, ZN => n18356);
   U13815 : OAI22_X1 port map( A1 => n21685, A2 => n15854, B1 => n21698, B2 => 
                           n16519, ZN => n18363);
   U13816 : BUF_X1 port map( A => n15150, Z => n22381);
   U13817 : BUF_X1 port map( A => n15149, Z => n22391);
   U13818 : BUF_X1 port map( A => n15148, Z => n22397);
   U13819 : BUF_X1 port map( A => n15147, Z => n22403);
   U13820 : BUF_X1 port map( A => n15146, Z => n22409);
   U13821 : BUF_X1 port map( A => n15145, Z => n22415);
   U13822 : BUF_X1 port map( A => n15144, Z => n22421);
   U13823 : BUF_X1 port map( A => n15143, Z => n22427);
   U13824 : BUF_X1 port map( A => n15142, Z => n22433);
   U13825 : BUF_X1 port map( A => n15141, Z => n22439);
   U13826 : BUF_X1 port map( A => n15140, Z => n22445);
   U13827 : BUF_X1 port map( A => n15139, Z => n22451);
   U13828 : BUF_X1 port map( A => n15138, Z => n22457);
   U13829 : BUF_X1 port map( A => n15137, Z => n22463);
   U13830 : BUF_X1 port map( A => n15136, Z => n22469);
   U13831 : BUF_X1 port map( A => n15135, Z => n22475);
   U13832 : BUF_X1 port map( A => n15134, Z => n22481);
   U13833 : BUF_X1 port map( A => n15133, Z => n22487);
   U13834 : BUF_X1 port map( A => n15132, Z => n22493);
   U13835 : BUF_X1 port map( A => n15131, Z => n22499);
   U13836 : BUF_X1 port map( A => n15130, Z => n22505);
   U13837 : BUF_X1 port map( A => n15129, Z => n22511);
   U13838 : BUF_X1 port map( A => n15128, Z => n22517);
   U13839 : BUF_X1 port map( A => n15127, Z => n22523);
   U13840 : BUF_X1 port map( A => n15126, Z => n22529);
   U13841 : BUF_X1 port map( A => n15125, Z => n22535);
   U13842 : BUF_X1 port map( A => n15124, Z => n22541);
   U13843 : BUF_X1 port map( A => n15123, Z => n22547);
   U13844 : BUF_X1 port map( A => n15122, Z => n22553);
   U13845 : BUF_X1 port map( A => n15121, Z => n22559);
   U13846 : BUF_X1 port map( A => n15120, Z => n22565);
   U13847 : BUF_X1 port map( A => n15118, Z => n22580);
   U13848 : BUF_X1 port map( A => n15150, Z => n22382);
   U13849 : BUF_X1 port map( A => n15149, Z => n22390);
   U13850 : BUF_X1 port map( A => n15148, Z => n22396);
   U13851 : BUF_X1 port map( A => n15147, Z => n22402);
   U13852 : BUF_X1 port map( A => n15146, Z => n22408);
   U13853 : BUF_X1 port map( A => n15145, Z => n22414);
   U13854 : BUF_X1 port map( A => n15144, Z => n22420);
   U13855 : BUF_X1 port map( A => n15143, Z => n22426);
   U13856 : BUF_X1 port map( A => n15142, Z => n22432);
   U13857 : BUF_X1 port map( A => n15141, Z => n22438);
   U13858 : BUF_X1 port map( A => n15140, Z => n22444);
   U13859 : BUF_X1 port map( A => n15139, Z => n22450);
   U13860 : BUF_X1 port map( A => n15138, Z => n22456);
   U13861 : BUF_X1 port map( A => n15137, Z => n22462);
   U13862 : BUF_X1 port map( A => n15136, Z => n22468);
   U13863 : BUF_X1 port map( A => n15135, Z => n22474);
   U13864 : BUF_X1 port map( A => n15134, Z => n22480);
   U13865 : BUF_X1 port map( A => n15133, Z => n22486);
   U13866 : BUF_X1 port map( A => n15132, Z => n22492);
   U13867 : BUF_X1 port map( A => n15131, Z => n22498);
   U13868 : BUF_X1 port map( A => n15130, Z => n22504);
   U13869 : BUF_X1 port map( A => n15129, Z => n22510);
   U13870 : BUF_X1 port map( A => n15128, Z => n22516);
   U13871 : BUF_X1 port map( A => n15127, Z => n22522);
   U13872 : BUF_X1 port map( A => n15126, Z => n22528);
   U13873 : BUF_X1 port map( A => n15125, Z => n22534);
   U13874 : BUF_X1 port map( A => n15124, Z => n22540);
   U13875 : BUF_X1 port map( A => n15123, Z => n22546);
   U13876 : BUF_X1 port map( A => n15122, Z => n22552);
   U13877 : BUF_X1 port map( A => n15121, Z => n22558);
   U13878 : BUF_X1 port map( A => n15120, Z => n22564);
   U13879 : BUF_X1 port map( A => n15118, Z => n22579);
   U13880 : BUF_X1 port map( A => n15150, Z => n22383);
   U13881 : BUF_X1 port map( A => n15149, Z => n22389);
   U13882 : BUF_X1 port map( A => n15148, Z => n22395);
   U13883 : BUF_X1 port map( A => n15147, Z => n22401);
   U13884 : BUF_X1 port map( A => n15146, Z => n22407);
   U13885 : BUF_X1 port map( A => n15145, Z => n22413);
   U13886 : BUF_X1 port map( A => n15144, Z => n22419);
   U13887 : BUF_X1 port map( A => n15143, Z => n22425);
   U13888 : BUF_X1 port map( A => n15142, Z => n22431);
   U13889 : BUF_X1 port map( A => n15141, Z => n22437);
   U13890 : BUF_X1 port map( A => n15140, Z => n22443);
   U13891 : BUF_X1 port map( A => n15139, Z => n22449);
   U13892 : BUF_X1 port map( A => n15138, Z => n22455);
   U13893 : BUF_X1 port map( A => n15137, Z => n22461);
   U13894 : BUF_X1 port map( A => n15136, Z => n22467);
   U13895 : BUF_X1 port map( A => n15135, Z => n22473);
   U13896 : BUF_X1 port map( A => n15134, Z => n22479);
   U13897 : BUF_X1 port map( A => n15133, Z => n22485);
   U13898 : BUF_X1 port map( A => n15132, Z => n22491);
   U13899 : BUF_X1 port map( A => n15131, Z => n22497);
   U13900 : BUF_X1 port map( A => n15130, Z => n22503);
   U13901 : BUF_X1 port map( A => n15129, Z => n22509);
   U13902 : BUF_X1 port map( A => n15128, Z => n22515);
   U13903 : BUF_X1 port map( A => n15127, Z => n22521);
   U13904 : BUF_X1 port map( A => n15126, Z => n22527);
   U13905 : BUF_X1 port map( A => n15125, Z => n22533);
   U13906 : BUF_X1 port map( A => n15124, Z => n22539);
   U13907 : BUF_X1 port map( A => n15123, Z => n22545);
   U13908 : BUF_X1 port map( A => n15122, Z => n22551);
   U13909 : BUF_X1 port map( A => n15121, Z => n22557);
   U13910 : BUF_X1 port map( A => n15120, Z => n22563);
   U13911 : BUF_X1 port map( A => n15118, Z => n22578);
   U13912 : BUF_X1 port map( A => n15150, Z => n22384);
   U13913 : BUF_X1 port map( A => n15149, Z => n22388);
   U13914 : BUF_X1 port map( A => n15148, Z => n22394);
   U13915 : BUF_X1 port map( A => n15147, Z => n22400);
   U13916 : BUF_X1 port map( A => n15146, Z => n22406);
   U13917 : BUF_X1 port map( A => n15145, Z => n22412);
   U13918 : BUF_X1 port map( A => n15144, Z => n22418);
   U13919 : BUF_X1 port map( A => n15143, Z => n22424);
   U13920 : BUF_X1 port map( A => n15142, Z => n22430);
   U13921 : BUF_X1 port map( A => n15141, Z => n22436);
   U13922 : BUF_X1 port map( A => n15140, Z => n22442);
   U13923 : BUF_X1 port map( A => n15139, Z => n22448);
   U13924 : BUF_X1 port map( A => n15138, Z => n22454);
   U13925 : BUF_X1 port map( A => n15137, Z => n22460);
   U13926 : BUF_X1 port map( A => n15136, Z => n22466);
   U13927 : BUF_X1 port map( A => n15135, Z => n22472);
   U13928 : BUF_X1 port map( A => n15134, Z => n22478);
   U13929 : BUF_X1 port map( A => n15133, Z => n22484);
   U13930 : BUF_X1 port map( A => n15132, Z => n22490);
   U13931 : BUF_X1 port map( A => n15131, Z => n22496);
   U13932 : BUF_X1 port map( A => n15130, Z => n22502);
   U13933 : BUF_X1 port map( A => n15129, Z => n22508);
   U13934 : BUF_X1 port map( A => n15128, Z => n22514);
   U13935 : BUF_X1 port map( A => n15127, Z => n22520);
   U13936 : BUF_X1 port map( A => n15126, Z => n22526);
   U13937 : BUF_X1 port map( A => n15125, Z => n22532);
   U13938 : BUF_X1 port map( A => n15124, Z => n22538);
   U13939 : BUF_X1 port map( A => n15123, Z => n22544);
   U13940 : BUF_X1 port map( A => n15122, Z => n22550);
   U13941 : BUF_X1 port map( A => n15121, Z => n22556);
   U13942 : BUF_X1 port map( A => n15120, Z => n22562);
   U13943 : BUF_X1 port map( A => n15118, Z => n22577);
   U13944 : BUF_X1 port map( A => n15150, Z => n22385);
   U13945 : BUF_X1 port map( A => n15149, Z => n22387);
   U13946 : BUF_X1 port map( A => n15148, Z => n22393);
   U13947 : BUF_X1 port map( A => n15147, Z => n22399);
   U13948 : BUF_X1 port map( A => n15146, Z => n22405);
   U13949 : BUF_X1 port map( A => n15145, Z => n22411);
   U13950 : BUF_X1 port map( A => n15144, Z => n22417);
   U13951 : BUF_X1 port map( A => n15143, Z => n22423);
   U13952 : BUF_X1 port map( A => n15142, Z => n22429);
   U13953 : BUF_X1 port map( A => n15141, Z => n22435);
   U13954 : BUF_X1 port map( A => n15140, Z => n22441);
   U13955 : BUF_X1 port map( A => n15139, Z => n22447);
   U13956 : BUF_X1 port map( A => n15138, Z => n22453);
   U13957 : BUF_X1 port map( A => n15137, Z => n22459);
   U13958 : BUF_X1 port map( A => n15136, Z => n22465);
   U13959 : BUF_X1 port map( A => n15135, Z => n22471);
   U13960 : BUF_X1 port map( A => n15134, Z => n22477);
   U13961 : BUF_X1 port map( A => n15133, Z => n22483);
   U13962 : BUF_X1 port map( A => n15132, Z => n22489);
   U13963 : BUF_X1 port map( A => n15131, Z => n22495);
   U13964 : BUF_X1 port map( A => n15130, Z => n22501);
   U13965 : BUF_X1 port map( A => n15129, Z => n22507);
   U13966 : BUF_X1 port map( A => n15128, Z => n22513);
   U13967 : BUF_X1 port map( A => n15127, Z => n22519);
   U13968 : BUF_X1 port map( A => n15126, Z => n22525);
   U13969 : BUF_X1 port map( A => n15125, Z => n22531);
   U13970 : BUF_X1 port map( A => n15124, Z => n22537);
   U13971 : BUF_X1 port map( A => n15123, Z => n22543);
   U13972 : BUF_X1 port map( A => n15122, Z => n22549);
   U13973 : BUF_X1 port map( A => n15121, Z => n22555);
   U13974 : BUF_X1 port map( A => n15120, Z => n22561);
   U13975 : BUF_X1 port map( A => n15118, Z => n22576);
   U13976 : OAI22_X1 port map( A1 => n21853, A2 => n22529, B1 => n16724, B2 => 
                           n16732, ZN => n5590);
   U13977 : OAI22_X1 port map( A1 => n21854, A2 => n22535, B1 => n16724, B2 => 
                           n16731, ZN => n5591);
   U13978 : OAI22_X1 port map( A1 => n21854, A2 => n22541, B1 => n16724, B2 => 
                           n16730, ZN => n5592);
   U13979 : OAI22_X1 port map( A1 => n21854, A2 => n22547, B1 => n21848, B2 => 
                           n16729, ZN => n5593);
   U13980 : OAI22_X1 port map( A1 => n21854, A2 => n22553, B1 => n21848, B2 => 
                           n16728, ZN => n5594);
   U13981 : OAI22_X1 port map( A1 => n21854, A2 => n22559, B1 => n21848, B2 => 
                           n16727, ZN => n5595);
   U13982 : OAI22_X1 port map( A1 => n21855, A2 => n22565, B1 => n21848, B2 => 
                           n16726, ZN => n5596);
   U13983 : OAI22_X1 port map( A1 => n21855, A2 => n22580, B1 => n16724, B2 => 
                           n16725, ZN => n5597);
   U13984 : OAI22_X1 port map( A1 => n21934, A2 => n22529, B1 => n16556, B2 => 
                           n16564, ZN => n5878);
   U13985 : OAI22_X1 port map( A1 => n21935, A2 => n22535, B1 => n16556, B2 => 
                           n16563, ZN => n5879);
   U13986 : OAI22_X1 port map( A1 => n21935, A2 => n22541, B1 => n16556, B2 => 
                           n16562, ZN => n5880);
   U13987 : OAI22_X1 port map( A1 => n21935, A2 => n22547, B1 => n21929, B2 => 
                           n16561, ZN => n5881);
   U13988 : OAI22_X1 port map( A1 => n21935, A2 => n22553, B1 => n21929, B2 => 
                           n16560, ZN => n5882);
   U13989 : OAI22_X1 port map( A1 => n21935, A2 => n22559, B1 => n21929, B2 => 
                           n16559, ZN => n5883);
   U13990 : OAI22_X1 port map( A1 => n21936, A2 => n22565, B1 => n21929, B2 => 
                           n16558, ZN => n5884);
   U13991 : OAI22_X1 port map( A1 => n21936, A2 => n22580, B1 => n16556, B2 => 
                           n16557, ZN => n5885);
   U13992 : OAI22_X1 port map( A1 => n21943, A2 => n22529, B1 => n16521, B2 => 
                           n16529, ZN => n5910);
   U13993 : OAI22_X1 port map( A1 => n21944, A2 => n22535, B1 => n16521, B2 => 
                           n16528, ZN => n5911);
   U13994 : OAI22_X1 port map( A1 => n21944, A2 => n22541, B1 => n16521, B2 => 
                           n16527, ZN => n5912);
   U13995 : OAI22_X1 port map( A1 => n21944, A2 => n22547, B1 => n21938, B2 => 
                           n16526, ZN => n5913);
   U13996 : OAI22_X1 port map( A1 => n21944, A2 => n22553, B1 => n21938, B2 => 
                           n16525, ZN => n5914);
   U13997 : OAI22_X1 port map( A1 => n21944, A2 => n22559, B1 => n21938, B2 => 
                           n16524, ZN => n5915);
   U13998 : OAI22_X1 port map( A1 => n21945, A2 => n22565, B1 => n21938, B2 => 
                           n16523, ZN => n5916);
   U13999 : OAI22_X1 port map( A1 => n21945, A2 => n22580, B1 => n16521, B2 => 
                           n16522, ZN => n5917);
   U14000 : OAI22_X1 port map( A1 => n21952, A2 => n22528, B1 => n16487, B2 => 
                           n16495, ZN => n5942);
   U14001 : OAI22_X1 port map( A1 => n21953, A2 => n22534, B1 => n16487, B2 => 
                           n16494, ZN => n5943);
   U14002 : OAI22_X1 port map( A1 => n21953, A2 => n22540, B1 => n16487, B2 => 
                           n16493, ZN => n5944);
   U14003 : OAI22_X1 port map( A1 => n21953, A2 => n22546, B1 => n21947, B2 => 
                           n16492, ZN => n5945);
   U14004 : OAI22_X1 port map( A1 => n21953, A2 => n22552, B1 => n21947, B2 => 
                           n16491, ZN => n5946);
   U14005 : OAI22_X1 port map( A1 => n21953, A2 => n22558, B1 => n21947, B2 => 
                           n16490, ZN => n5947);
   U14006 : OAI22_X1 port map( A1 => n21954, A2 => n22564, B1 => n21947, B2 => 
                           n16489, ZN => n5948);
   U14007 : OAI22_X1 port map( A1 => n21954, A2 => n22579, B1 => n16487, B2 => 
                           n16488, ZN => n5949);
   U14008 : OAI22_X1 port map( A1 => n21988, A2 => n22528, B1 => n16350, B2 => 
                           n16358, ZN => n6070);
   U14009 : OAI22_X1 port map( A1 => n21989, A2 => n22534, B1 => n16350, B2 => 
                           n16357, ZN => n6071);
   U14010 : OAI22_X1 port map( A1 => n21989, A2 => n22540, B1 => n16350, B2 => 
                           n16356, ZN => n6072);
   U14011 : OAI22_X1 port map( A1 => n21989, A2 => n22546, B1 => n21983, B2 => 
                           n16355, ZN => n6073);
   U14012 : OAI22_X1 port map( A1 => n21989, A2 => n22552, B1 => n21983, B2 => 
                           n16354, ZN => n6074);
   U14013 : OAI22_X1 port map( A1 => n21989, A2 => n22558, B1 => n21983, B2 => 
                           n16353, ZN => n6075);
   U14014 : OAI22_X1 port map( A1 => n21990, A2 => n22564, B1 => n21983, B2 => 
                           n16352, ZN => n6076);
   U14015 : OAI22_X1 port map( A1 => n21990, A2 => n22579, B1 => n16350, B2 => 
                           n16351, ZN => n6077);
   U14016 : OAI22_X1 port map( A1 => n22024, A2 => n22528, B1 => n16309, B2 => 
                           n16317, ZN => n6198);
   U14017 : OAI22_X1 port map( A1 => n22025, A2 => n22534, B1 => n16309, B2 => 
                           n16316, ZN => n6199);
   U14018 : OAI22_X1 port map( A1 => n22025, A2 => n22540, B1 => n16309, B2 => 
                           n16315, ZN => n6200);
   U14019 : OAI22_X1 port map( A1 => n22025, A2 => n22546, B1 => n22019, B2 => 
                           n16314, ZN => n6201);
   U14020 : OAI22_X1 port map( A1 => n22025, A2 => n22552, B1 => n22019, B2 => 
                           n16313, ZN => n6202);
   U14021 : OAI22_X1 port map( A1 => n22025, A2 => n22558, B1 => n22019, B2 => 
                           n16312, ZN => n6203);
   U14022 : OAI22_X1 port map( A1 => n22026, A2 => n22564, B1 => n22019, B2 => 
                           n16311, ZN => n6204);
   U14023 : OAI22_X1 port map( A1 => n22026, A2 => n22579, B1 => n16309, B2 => 
                           n16310, ZN => n6205);
   U14024 : OAI22_X1 port map( A1 => n22042, A2 => n22528, B1 => n16241, B2 => 
                           n16249, ZN => n6262);
   U14025 : OAI22_X1 port map( A1 => n22043, A2 => n22534, B1 => n16241, B2 => 
                           n16248, ZN => n6263);
   U14026 : OAI22_X1 port map( A1 => n22043, A2 => n22540, B1 => n16241, B2 => 
                           n16247, ZN => n6264);
   U14027 : OAI22_X1 port map( A1 => n22043, A2 => n22546, B1 => n22037, B2 => 
                           n16246, ZN => n6265);
   U14028 : OAI22_X1 port map( A1 => n22043, A2 => n22552, B1 => n22037, B2 => 
                           n16245, ZN => n6266);
   U14029 : OAI22_X1 port map( A1 => n22043, A2 => n22558, B1 => n22037, B2 => 
                           n16244, ZN => n6267);
   U14030 : OAI22_X1 port map( A1 => n22044, A2 => n22564, B1 => n22037, B2 => 
                           n16243, ZN => n6268);
   U14031 : OAI22_X1 port map( A1 => n22044, A2 => n22579, B1 => n16241, B2 => 
                           n16242, ZN => n6269);
   U14032 : OAI22_X1 port map( A1 => n22051, A2 => n22528, B1 => n16206, B2 => 
                           n16214, ZN => n6294);
   U14033 : OAI22_X1 port map( A1 => n22052, A2 => n22534, B1 => n16206, B2 => 
                           n16213, ZN => n6295);
   U14034 : OAI22_X1 port map( A1 => n22052, A2 => n22540, B1 => n16206, B2 => 
                           n16212, ZN => n6296);
   U14035 : OAI22_X1 port map( A1 => n22052, A2 => n22546, B1 => n22046, B2 => 
                           n16211, ZN => n6297);
   U14036 : OAI22_X1 port map( A1 => n22052, A2 => n22552, B1 => n22046, B2 => 
                           n16210, ZN => n6298);
   U14037 : OAI22_X1 port map( A1 => n22052, A2 => n22558, B1 => n22046, B2 => 
                           n16209, ZN => n6299);
   U14038 : OAI22_X1 port map( A1 => n22053, A2 => n22564, B1 => n22046, B2 => 
                           n16208, ZN => n6300);
   U14039 : OAI22_X1 port map( A1 => n22053, A2 => n22579, B1 => n16206, B2 => 
                           n16207, ZN => n6301);
   U14040 : OAI22_X1 port map( A1 => n22060, A2 => n22527, B1 => n16171, B2 => 
                           n16179, ZN => n6326);
   U14041 : OAI22_X1 port map( A1 => n22061, A2 => n22533, B1 => n16171, B2 => 
                           n16178, ZN => n6327);
   U14042 : OAI22_X1 port map( A1 => n22061, A2 => n22539, B1 => n16171, B2 => 
                           n16177, ZN => n6328);
   U14043 : OAI22_X1 port map( A1 => n22061, A2 => n22545, B1 => n22055, B2 => 
                           n16176, ZN => n6329);
   U14044 : OAI22_X1 port map( A1 => n22061, A2 => n22551, B1 => n22055, B2 => 
                           n16175, ZN => n6330);
   U14045 : OAI22_X1 port map( A1 => n22061, A2 => n22557, B1 => n22055, B2 => 
                           n16174, ZN => n6331);
   U14046 : OAI22_X1 port map( A1 => n22062, A2 => n22563, B1 => n22055, B2 => 
                           n16173, ZN => n6332);
   U14047 : OAI22_X1 port map( A1 => n22062, A2 => n22578, B1 => n16171, B2 => 
                           n16172, ZN => n6333);
   U14048 : OAI22_X1 port map( A1 => n22078, A2 => n22527, B1 => n16135, B2 => 
                           n16143, ZN => n6390);
   U14049 : OAI22_X1 port map( A1 => n22079, A2 => n22533, B1 => n16135, B2 => 
                           n16142, ZN => n6391);
   U14050 : OAI22_X1 port map( A1 => n22079, A2 => n22539, B1 => n16135, B2 => 
                           n16141, ZN => n6392);
   U14051 : OAI22_X1 port map( A1 => n22079, A2 => n22545, B1 => n22073, B2 => 
                           n16140, ZN => n6393);
   U14052 : OAI22_X1 port map( A1 => n22079, A2 => n22551, B1 => n22073, B2 => 
                           n16139, ZN => n6394);
   U14053 : OAI22_X1 port map( A1 => n22079, A2 => n22557, B1 => n22073, B2 => 
                           n16138, ZN => n6395);
   U14054 : OAI22_X1 port map( A1 => n22080, A2 => n22563, B1 => n22073, B2 => 
                           n16137, ZN => n6396);
   U14055 : OAI22_X1 port map( A1 => n22080, A2 => n22578, B1 => n16135, B2 => 
                           n16136, ZN => n6397);
   U14056 : OAI22_X1 port map( A1 => n22087, A2 => n22527, B1 => n16100, B2 => 
                           n16108, ZN => n6422);
   U14057 : OAI22_X1 port map( A1 => n22088, A2 => n22533, B1 => n16100, B2 => 
                           n16107, ZN => n6423);
   U14058 : OAI22_X1 port map( A1 => n22088, A2 => n22539, B1 => n16100, B2 => 
                           n16106, ZN => n6424);
   U14059 : OAI22_X1 port map( A1 => n22088, A2 => n22545, B1 => n22082, B2 => 
                           n16105, ZN => n6425);
   U14060 : OAI22_X1 port map( A1 => n22088, A2 => n22551, B1 => n22082, B2 => 
                           n16104, ZN => n6426);
   U14061 : OAI22_X1 port map( A1 => n22088, A2 => n22557, B1 => n22082, B2 => 
                           n16103, ZN => n6427);
   U14062 : OAI22_X1 port map( A1 => n22089, A2 => n22563, B1 => n22082, B2 => 
                           n16102, ZN => n6428);
   U14063 : OAI22_X1 port map( A1 => n22089, A2 => n22578, B1 => n16100, B2 => 
                           n16101, ZN => n6429);
   U14064 : OAI22_X1 port map( A1 => n22096, A2 => n22527, B1 => n16066, B2 => 
                           n16074, ZN => n6454);
   U14065 : OAI22_X1 port map( A1 => n22097, A2 => n22533, B1 => n16066, B2 => 
                           n16073, ZN => n6455);
   U14066 : OAI22_X1 port map( A1 => n22097, A2 => n22539, B1 => n16066, B2 => 
                           n16072, ZN => n6456);
   U14067 : OAI22_X1 port map( A1 => n22097, A2 => n22545, B1 => n22091, B2 => 
                           n16071, ZN => n6457);
   U14068 : OAI22_X1 port map( A1 => n22097, A2 => n22551, B1 => n22091, B2 => 
                           n16070, ZN => n6458);
   U14069 : OAI22_X1 port map( A1 => n22097, A2 => n22557, B1 => n22091, B2 => 
                           n16069, ZN => n6459);
   U14070 : OAI22_X1 port map( A1 => n22098, A2 => n22563, B1 => n22091, B2 => 
                           n16068, ZN => n6460);
   U14071 : OAI22_X1 port map( A1 => n22098, A2 => n22578, B1 => n16066, B2 => 
                           n16067, ZN => n6461);
   U14072 : OAI22_X1 port map( A1 => n22105, A2 => n22527, B1 => n16032, B2 => 
                           n16040, ZN => n6486);
   U14073 : OAI22_X1 port map( A1 => n22106, A2 => n22533, B1 => n16032, B2 => 
                           n16039, ZN => n6487);
   U14074 : OAI22_X1 port map( A1 => n22106, A2 => n22539, B1 => n16032, B2 => 
                           n16038, ZN => n6488);
   U14075 : OAI22_X1 port map( A1 => n22106, A2 => n22545, B1 => n22100, B2 => 
                           n16037, ZN => n6489);
   U14076 : OAI22_X1 port map( A1 => n22106, A2 => n22551, B1 => n22100, B2 => 
                           n16036, ZN => n6490);
   U14077 : OAI22_X1 port map( A1 => n22106, A2 => n22557, B1 => n22100, B2 => 
                           n16035, ZN => n6491);
   U14078 : OAI22_X1 port map( A1 => n22107, A2 => n22563, B1 => n22100, B2 => 
                           n16034, ZN => n6492);
   U14079 : OAI22_X1 port map( A1 => n22107, A2 => n22578, B1 => n16032, B2 => 
                           n16033, ZN => n6493);
   U14080 : OAI22_X1 port map( A1 => n22141, A2 => n22527, B1 => n15895, B2 => 
                           n15903, ZN => n6614);
   U14081 : OAI22_X1 port map( A1 => n22142, A2 => n22533, B1 => n15895, B2 => 
                           n15902, ZN => n6615);
   U14082 : OAI22_X1 port map( A1 => n22142, A2 => n22539, B1 => n15895, B2 => 
                           n15901, ZN => n6616);
   U14083 : OAI22_X1 port map( A1 => n22142, A2 => n22545, B1 => n22136, B2 => 
                           n15900, ZN => n6617);
   U14084 : OAI22_X1 port map( A1 => n22142, A2 => n22551, B1 => n22136, B2 => 
                           n15899, ZN => n6618);
   U14085 : OAI22_X1 port map( A1 => n22142, A2 => n22557, B1 => n22136, B2 => 
                           n15898, ZN => n6619);
   U14086 : OAI22_X1 port map( A1 => n22143, A2 => n22563, B1 => n22136, B2 => 
                           n15897, ZN => n6620);
   U14087 : OAI22_X1 port map( A1 => n22143, A2 => n22578, B1 => n15895, B2 => 
                           n15896, ZN => n6621);
   U14088 : OAI22_X1 port map( A1 => n22177, A2 => n22526, B1 => n15822, B2 => 
                           n15830, ZN => n6742);
   U14089 : OAI22_X1 port map( A1 => n22178, A2 => n22532, B1 => n15822, B2 => 
                           n15829, ZN => n6743);
   U14090 : OAI22_X1 port map( A1 => n22178, A2 => n22538, B1 => n15822, B2 => 
                           n15828, ZN => n6744);
   U14091 : OAI22_X1 port map( A1 => n22178, A2 => n22544, B1 => n22172, B2 => 
                           n15827, ZN => n6745);
   U14092 : OAI22_X1 port map( A1 => n22178, A2 => n22550, B1 => n22172, B2 => 
                           n15826, ZN => n6746);
   U14093 : OAI22_X1 port map( A1 => n22178, A2 => n22556, B1 => n22172, B2 => 
                           n15825, ZN => n6747);
   U14094 : OAI22_X1 port map( A1 => n22179, A2 => n22562, B1 => n22172, B2 => 
                           n15824, ZN => n6748);
   U14095 : OAI22_X1 port map( A1 => n22179, A2 => n22577, B1 => n15822, B2 => 
                           n15823, ZN => n6749);
   U14096 : OAI22_X1 port map( A1 => n22186, A2 => n22526, B1 => n15788, B2 => 
                           n15796, ZN => n6774);
   U14097 : OAI22_X1 port map( A1 => n22187, A2 => n22532, B1 => n15788, B2 => 
                           n15795, ZN => n6775);
   U14098 : OAI22_X1 port map( A1 => n22187, A2 => n22538, B1 => n15788, B2 => 
                           n15794, ZN => n6776);
   U14099 : OAI22_X1 port map( A1 => n22187, A2 => n22544, B1 => n22181, B2 => 
                           n15793, ZN => n6777);
   U14100 : OAI22_X1 port map( A1 => n22187, A2 => n22550, B1 => n22181, B2 => 
                           n15792, ZN => n6778);
   U14101 : OAI22_X1 port map( A1 => n22187, A2 => n22556, B1 => n22181, B2 => 
                           n15791, ZN => n6779);
   U14102 : OAI22_X1 port map( A1 => n22188, A2 => n22562, B1 => n22181, B2 => 
                           n15790, ZN => n6780);
   U14103 : OAI22_X1 port map( A1 => n22188, A2 => n22577, B1 => n15788, B2 => 
                           n15789, ZN => n6781);
   U14104 : OAI22_X1 port map( A1 => n22195, A2 => n22526, B1 => n15753, B2 => 
                           n15761, ZN => n6806);
   U14105 : OAI22_X1 port map( A1 => n22196, A2 => n22532, B1 => n15753, B2 => 
                           n15760, ZN => n6807);
   U14106 : OAI22_X1 port map( A1 => n22196, A2 => n22538, B1 => n15753, B2 => 
                           n15759, ZN => n6808);
   U14107 : OAI22_X1 port map( A1 => n22196, A2 => n22544, B1 => n22190, B2 => 
                           n15758, ZN => n6809);
   U14108 : OAI22_X1 port map( A1 => n22196, A2 => n22550, B1 => n22190, B2 => 
                           n15757, ZN => n6810);
   U14109 : OAI22_X1 port map( A1 => n22196, A2 => n22556, B1 => n22190, B2 => 
                           n15756, ZN => n6811);
   U14110 : OAI22_X1 port map( A1 => n22197, A2 => n22562, B1 => n22190, B2 => 
                           n15755, ZN => n6812);
   U14111 : OAI22_X1 port map( A1 => n22197, A2 => n22577, B1 => n15753, B2 => 
                           n15754, ZN => n6813);
   U14112 : OAI22_X1 port map( A1 => n22222, A2 => n22526, B1 => n15682, B2 => 
                           n15690, ZN => n6902);
   U14113 : OAI22_X1 port map( A1 => n22223, A2 => n22532, B1 => n15682, B2 => 
                           n15689, ZN => n6903);
   U14114 : OAI22_X1 port map( A1 => n22223, A2 => n22538, B1 => n15682, B2 => 
                           n15688, ZN => n6904);
   U14115 : OAI22_X1 port map( A1 => n22223, A2 => n22544, B1 => n22217, B2 => 
                           n15687, ZN => n6905);
   U14116 : OAI22_X1 port map( A1 => n22223, A2 => n22550, B1 => n22217, B2 => 
                           n15686, ZN => n6906);
   U14117 : OAI22_X1 port map( A1 => n22223, A2 => n22556, B1 => n22217, B2 => 
                           n15685, ZN => n6907);
   U14118 : OAI22_X1 port map( A1 => n22224, A2 => n22562, B1 => n22217, B2 => 
                           n15684, ZN => n6908);
   U14119 : OAI22_X1 port map( A1 => n22224, A2 => n22577, B1 => n15682, B2 => 
                           n15683, ZN => n6909);
   U14120 : OAI22_X1 port map( A1 => n22231, A2 => n22526, B1 => n15647, B2 => 
                           n15655, ZN => n6934);
   U14121 : OAI22_X1 port map( A1 => n22232, A2 => n22532, B1 => n15647, B2 => 
                           n15654, ZN => n6935);
   U14122 : OAI22_X1 port map( A1 => n22232, A2 => n22538, B1 => n15647, B2 => 
                           n15653, ZN => n6936);
   U14123 : OAI22_X1 port map( A1 => n22232, A2 => n22544, B1 => n22226, B2 => 
                           n15652, ZN => n6937);
   U14124 : OAI22_X1 port map( A1 => n22232, A2 => n22550, B1 => n22226, B2 => 
                           n15651, ZN => n6938);
   U14125 : OAI22_X1 port map( A1 => n22232, A2 => n22556, B1 => n22226, B2 => 
                           n15650, ZN => n6939);
   U14126 : OAI22_X1 port map( A1 => n22233, A2 => n22562, B1 => n22226, B2 => 
                           n15649, ZN => n6940);
   U14127 : OAI22_X1 port map( A1 => n22233, A2 => n22577, B1 => n15647, B2 => 
                           n15648, ZN => n6941);
   U14128 : OAI22_X1 port map( A1 => n22249, A2 => n22526, B1 => n15575, B2 => 
                           n15583, ZN => n6998);
   U14129 : OAI22_X1 port map( A1 => n22250, A2 => n22532, B1 => n15575, B2 => 
                           n15582, ZN => n6999);
   U14130 : OAI22_X1 port map( A1 => n22250, A2 => n22538, B1 => n15575, B2 => 
                           n15581, ZN => n7000);
   U14131 : OAI22_X1 port map( A1 => n22250, A2 => n22544, B1 => n22244, B2 => 
                           n15580, ZN => n7001);
   U14132 : OAI22_X1 port map( A1 => n22250, A2 => n22550, B1 => n22244, B2 => 
                           n15579, ZN => n7002);
   U14133 : OAI22_X1 port map( A1 => n22250, A2 => n22556, B1 => n22244, B2 => 
                           n15578, ZN => n7003);
   U14134 : OAI22_X1 port map( A1 => n22251, A2 => n22562, B1 => n22244, B2 => 
                           n15577, ZN => n7004);
   U14135 : OAI22_X1 port map( A1 => n22251, A2 => n22577, B1 => n15575, B2 => 
                           n15576, ZN => n7005);
   U14136 : OAI22_X1 port map( A1 => n22276, A2 => n22525, B1 => n15471, B2 => 
                           n15479, ZN => n7094);
   U14137 : OAI22_X1 port map( A1 => n22277, A2 => n22531, B1 => n15471, B2 => 
                           n15478, ZN => n7095);
   U14138 : OAI22_X1 port map( A1 => n22277, A2 => n22537, B1 => n15471, B2 => 
                           n15477, ZN => n7096);
   U14139 : OAI22_X1 port map( A1 => n22277, A2 => n22543, B1 => n22271, B2 => 
                           n15476, ZN => n7097);
   U14140 : OAI22_X1 port map( A1 => n22277, A2 => n22549, B1 => n22271, B2 => 
                           n15475, ZN => n7098);
   U14141 : OAI22_X1 port map( A1 => n22277, A2 => n22555, B1 => n22271, B2 => 
                           n15474, ZN => n7099);
   U14142 : OAI22_X1 port map( A1 => n22278, A2 => n22561, B1 => n22271, B2 => 
                           n15473, ZN => n7100);
   U14143 : OAI22_X1 port map( A1 => n22278, A2 => n22576, B1 => n15471, B2 => 
                           n15472, ZN => n7101);
   U14144 : OAI22_X1 port map( A1 => n22285, A2 => n22525, B1 => n15437, B2 => 
                           n15445, ZN => n7126);
   U14145 : OAI22_X1 port map( A1 => n22286, A2 => n22531, B1 => n15437, B2 => 
                           n15444, ZN => n7127);
   U14146 : OAI22_X1 port map( A1 => n22286, A2 => n22537, B1 => n15437, B2 => 
                           n15443, ZN => n7128);
   U14147 : OAI22_X1 port map( A1 => n22286, A2 => n22543, B1 => n22280, B2 => 
                           n15442, ZN => n7129);
   U14148 : OAI22_X1 port map( A1 => n22286, A2 => n22549, B1 => n22280, B2 => 
                           n15441, ZN => n7130);
   U14149 : OAI22_X1 port map( A1 => n22286, A2 => n22555, B1 => n22280, B2 => 
                           n15440, ZN => n7131);
   U14150 : OAI22_X1 port map( A1 => n22287, A2 => n22561, B1 => n22280, B2 => 
                           n15439, ZN => n7132);
   U14151 : OAI22_X1 port map( A1 => n22287, A2 => n22576, B1 => n15437, B2 => 
                           n15438, ZN => n7133);
   U14152 : OAI22_X1 port map( A1 => n22294, A2 => n22525, B1 => n15403, B2 => 
                           n15411, ZN => n7158);
   U14153 : OAI22_X1 port map( A1 => n22295, A2 => n22531, B1 => n15403, B2 => 
                           n15410, ZN => n7159);
   U14154 : OAI22_X1 port map( A1 => n22295, A2 => n22537, B1 => n15403, B2 => 
                           n15409, ZN => n7160);
   U14155 : OAI22_X1 port map( A1 => n22295, A2 => n22543, B1 => n22289, B2 => 
                           n15408, ZN => n7161);
   U14156 : OAI22_X1 port map( A1 => n22295, A2 => n22549, B1 => n22289, B2 => 
                           n15407, ZN => n7162);
   U14157 : OAI22_X1 port map( A1 => n22295, A2 => n22555, B1 => n22289, B2 => 
                           n15406, ZN => n7163);
   U14158 : OAI22_X1 port map( A1 => n22296, A2 => n22561, B1 => n22289, B2 => 
                           n15405, ZN => n7164);
   U14159 : OAI22_X1 port map( A1 => n22296, A2 => n22576, B1 => n15403, B2 => 
                           n15404, ZN => n7165);
   U14160 : OAI22_X1 port map( A1 => n22303, A2 => n22525, B1 => n15368, B2 => 
                           n15376, ZN => n7190);
   U14161 : OAI22_X1 port map( A1 => n22304, A2 => n22531, B1 => n15368, B2 => 
                           n15375, ZN => n7191);
   U14162 : OAI22_X1 port map( A1 => n22304, A2 => n22537, B1 => n15368, B2 => 
                           n15374, ZN => n7192);
   U14163 : OAI22_X1 port map( A1 => n22304, A2 => n22543, B1 => n22298, B2 => 
                           n15373, ZN => n7193);
   U14164 : OAI22_X1 port map( A1 => n22304, A2 => n22549, B1 => n22298, B2 => 
                           n15372, ZN => n7194);
   U14165 : OAI22_X1 port map( A1 => n22304, A2 => n22555, B1 => n22298, B2 => 
                           n15371, ZN => n7195);
   U14166 : OAI22_X1 port map( A1 => n22305, A2 => n22561, B1 => n22298, B2 => 
                           n15370, ZN => n7196);
   U14167 : OAI22_X1 port map( A1 => n22305, A2 => n22576, B1 => n15368, B2 => 
                           n15369, ZN => n7197);
   U14168 : OAI22_X1 port map( A1 => n22330, A2 => n22525, B1 => n15265, B2 => 
                           n15273, ZN => n7286);
   U14169 : OAI22_X1 port map( A1 => n22331, A2 => n22531, B1 => n15265, B2 => 
                           n15272, ZN => n7287);
   U14170 : OAI22_X1 port map( A1 => n22331, A2 => n22537, B1 => n15265, B2 => 
                           n15271, ZN => n7288);
   U14171 : OAI22_X1 port map( A1 => n22331, A2 => n22543, B1 => n22325, B2 => 
                           n15270, ZN => n7289);
   U14172 : OAI22_X1 port map( A1 => n22331, A2 => n22549, B1 => n22325, B2 => 
                           n15269, ZN => n7290);
   U14173 : OAI22_X1 port map( A1 => n22331, A2 => n22555, B1 => n22325, B2 => 
                           n15268, ZN => n7291);
   U14174 : OAI22_X1 port map( A1 => n22332, A2 => n22561, B1 => n22325, B2 => 
                           n15267, ZN => n7292);
   U14175 : OAI22_X1 port map( A1 => n22332, A2 => n22576, B1 => n15265, B2 => 
                           n15266, ZN => n7293);
   U14176 : OAI22_X1 port map( A1 => n22339, A2 => n22525, B1 => n15230, B2 => 
                           n15238, ZN => n7318);
   U14177 : OAI22_X1 port map( A1 => n22340, A2 => n22531, B1 => n15230, B2 => 
                           n15237, ZN => n7319);
   U14178 : OAI22_X1 port map( A1 => n22340, A2 => n22537, B1 => n15230, B2 => 
                           n15236, ZN => n7320);
   U14179 : OAI22_X1 port map( A1 => n22340, A2 => n22543, B1 => n22334, B2 => 
                           n15235, ZN => n7321);
   U14180 : OAI22_X1 port map( A1 => n22340, A2 => n22549, B1 => n22334, B2 => 
                           n15234, ZN => n7322);
   U14181 : OAI22_X1 port map( A1 => n22340, A2 => n22555, B1 => n22334, B2 => 
                           n15233, ZN => n7323);
   U14182 : OAI22_X1 port map( A1 => n22341, A2 => n22561, B1 => n22334, B2 => 
                           n15232, ZN => n7324);
   U14183 : OAI22_X1 port map( A1 => n22341, A2 => n22576, B1 => n15230, B2 => 
                           n15231, ZN => n7325);
   U14184 : NAND2_X1 port map( A1 => n19625, A2 => n19633, ZN => n18428);
   U14185 : NAND2_X1 port map( A1 => n18352, A2 => n18360, ZN => n16845);
   U14186 : NAND2_X1 port map( A1 => n19625, A2 => n19635, ZN => n18435);
   U14187 : NAND2_X1 port map( A1 => n19625, A2 => n19624, ZN => n18445);
   U14188 : NAND2_X1 port map( A1 => n18352, A2 => n18362, ZN => n16853);
   U14189 : NAND2_X1 port map( A1 => n18352, A2 => n18351, ZN => n16863);
   U14190 : NAND2_X1 port map( A1 => n19625, A2 => n20812, ZN => n18498);
   U14191 : NAND2_X1 port map( A1 => n19625, A2 => n20757, ZN => n18504);
   U14192 : NAND2_X1 port map( A1 => n19625, A2 => n20693, ZN => n18503);
   U14193 : NAND2_X1 port map( A1 => n19625, A2 => n20999, ZN => n18430);
   U14194 : NAND2_X1 port map( A1 => n19625, A2 => n21044, ZN => n18439);
   U14195 : NAND2_X1 port map( A1 => n18352, A2 => n21369, ZN => n16925);
   U14196 : NAND2_X1 port map( A1 => n18352, A2 => n21314, ZN => n16931);
   U14197 : NAND2_X1 port map( A1 => n18352, A2 => n21250, ZN => n16930);
   U14198 : NAND2_X1 port map( A1 => n18352, A2 => n21556, ZN => n16847);
   U14199 : NAND2_X1 port map( A1 => n18352, A2 => n21601, ZN => n16857);
   U14200 : BUF_X1 port map( A => n18468, Z => n20991);
   U14201 : BUF_X1 port map( A => n16888, Z => n21548);
   U14202 : BUF_X1 port map( A => n18463, Z => n21036);
   U14203 : BUF_X1 port map( A => n16882, Z => n21593);
   U14204 : BUF_X1 port map( A => n18468, Z => n20987);
   U14205 : BUF_X1 port map( A => n16888, Z => n21544);
   U14206 : BUF_X1 port map( A => n18463, Z => n21032);
   U14207 : BUF_X1 port map( A => n18468, Z => n20989);
   U14208 : BUF_X1 port map( A => n18463, Z => n21034);
   U14209 : BUF_X1 port map( A => n18468, Z => n20988);
   U14210 : BUF_X1 port map( A => n18463, Z => n21033);
   U14211 : BUF_X1 port map( A => n18468, Z => n20990);
   U14212 : BUF_X1 port map( A => n18463, Z => n21035);
   U14213 : BUF_X1 port map( A => n16882, Z => n21589);
   U14214 : BUF_X1 port map( A => n16888, Z => n21546);
   U14215 : BUF_X1 port map( A => n16882, Z => n21591);
   U14216 : BUF_X1 port map( A => n16888, Z => n21545);
   U14217 : BUF_X1 port map( A => n16882, Z => n21590);
   U14218 : BUF_X1 port map( A => n16888, Z => n21547);
   U14219 : BUF_X1 port map( A => n16882, Z => n21592);
   U14220 : OAI22_X1 port map( A1 => n21932, A2 => n22469, B1 => n21929, B2 => 
                           n16574, ZN => n5868);
   U14221 : OAI22_X1 port map( A1 => n21933, A2 => n22475, B1 => n21929, B2 => 
                           n16573, ZN => n5869);
   U14222 : OAI22_X1 port map( A1 => n21933, A2 => n22481, B1 => n21929, B2 => 
                           n16572, ZN => n5870);
   U14223 : OAI22_X1 port map( A1 => n21933, A2 => n22487, B1 => n21929, B2 => 
                           n16571, ZN => n5871);
   U14224 : OAI22_X1 port map( A1 => n21933, A2 => n22493, B1 => n21929, B2 => 
                           n16570, ZN => n5872);
   U14225 : OAI22_X1 port map( A1 => n21933, A2 => n22499, B1 => n21929, B2 => 
                           n16569, ZN => n5873);
   U14226 : OAI22_X1 port map( A1 => n21934, A2 => n22505, B1 => n21929, B2 => 
                           n16568, ZN => n5874);
   U14227 : OAI22_X1 port map( A1 => n21934, A2 => n22511, B1 => n21929, B2 => 
                           n16567, ZN => n5875);
   U14228 : OAI22_X1 port map( A1 => n21934, A2 => n22517, B1 => n21929, B2 => 
                           n16566, ZN => n5876);
   U14229 : OAI22_X1 port map( A1 => n21934, A2 => n22523, B1 => n21929, B2 => 
                           n16565, ZN => n5877);
   U14230 : OAI22_X1 port map( A1 => n21849, A2 => n22381, B1 => n21848, B2 => 
                           n16756, ZN => n5566);
   U14231 : OAI22_X1 port map( A1 => n21849, A2 => n22391, B1 => n21848, B2 => 
                           n16755, ZN => n5567);
   U14232 : OAI22_X1 port map( A1 => n21849, A2 => n22397, B1 => n21848, B2 => 
                           n16754, ZN => n5568);
   U14233 : OAI22_X1 port map( A1 => n21849, A2 => n22403, B1 => n21848, B2 => 
                           n16753, ZN => n5569);
   U14234 : OAI22_X1 port map( A1 => n21849, A2 => n22409, B1 => n21848, B2 => 
                           n16752, ZN => n5570);
   U14235 : OAI22_X1 port map( A1 => n21850, A2 => n22415, B1 => n21848, B2 => 
                           n16751, ZN => n5571);
   U14236 : OAI22_X1 port map( A1 => n21850, A2 => n22421, B1 => n21848, B2 => 
                           n16750, ZN => n5572);
   U14237 : OAI22_X1 port map( A1 => n21850, A2 => n22427, B1 => n21848, B2 => 
                           n16749, ZN => n5573);
   U14238 : OAI22_X1 port map( A1 => n21850, A2 => n22433, B1 => n21848, B2 => 
                           n16748, ZN => n5574);
   U14239 : OAI22_X1 port map( A1 => n21850, A2 => n22439, B1 => n21848, B2 => 
                           n16747, ZN => n5575);
   U14240 : OAI22_X1 port map( A1 => n21851, A2 => n22445, B1 => n21848, B2 => 
                           n16746, ZN => n5576);
   U14241 : OAI22_X1 port map( A1 => n21851, A2 => n22451, B1 => n21848, B2 => 
                           n16745, ZN => n5577);
   U14242 : OAI22_X1 port map( A1 => n21851, A2 => n22457, B1 => n21848, B2 => 
                           n16744, ZN => n5578);
   U14243 : OAI22_X1 port map( A1 => n21851, A2 => n22463, B1 => n21848, B2 => 
                           n16743, ZN => n5579);
   U14244 : OAI22_X1 port map( A1 => n21851, A2 => n22469, B1 => n16724, B2 => 
                           n16742, ZN => n5580);
   U14245 : OAI22_X1 port map( A1 => n21852, A2 => n22475, B1 => n16724, B2 => 
                           n16741, ZN => n5581);
   U14246 : OAI22_X1 port map( A1 => n21852, A2 => n22481, B1 => n16724, B2 => 
                           n16740, ZN => n5582);
   U14247 : OAI22_X1 port map( A1 => n21852, A2 => n22487, B1 => n16724, B2 => 
                           n16739, ZN => n5583);
   U14248 : OAI22_X1 port map( A1 => n21852, A2 => n22493, B1 => n16724, B2 => 
                           n16738, ZN => n5584);
   U14249 : OAI22_X1 port map( A1 => n21852, A2 => n22499, B1 => n16724, B2 => 
                           n16737, ZN => n5585);
   U14250 : OAI22_X1 port map( A1 => n21853, A2 => n22505, B1 => n16724, B2 => 
                           n16736, ZN => n5586);
   U14251 : OAI22_X1 port map( A1 => n21853, A2 => n22511, B1 => n21848, B2 => 
                           n16735, ZN => n5587);
   U14252 : OAI22_X1 port map( A1 => n21853, A2 => n22517, B1 => n21848, B2 => 
                           n16734, ZN => n5588);
   U14253 : OAI22_X1 port map( A1 => n21853, A2 => n22523, B1 => n21848, B2 => 
                           n16733, ZN => n5589);
   U14254 : OAI22_X1 port map( A1 => n21939, A2 => n22382, B1 => n21938, B2 => 
                           n16553, ZN => n5886);
   U14255 : OAI22_X1 port map( A1 => n21939, A2 => n22391, B1 => n21938, B2 => 
                           n16552, ZN => n5887);
   U14256 : OAI22_X1 port map( A1 => n21939, A2 => n22397, B1 => n21938, B2 => 
                           n16551, ZN => n5888);
   U14257 : OAI22_X1 port map( A1 => n21939, A2 => n22403, B1 => n21938, B2 => 
                           n16550, ZN => n5889);
   U14258 : OAI22_X1 port map( A1 => n21939, A2 => n22409, B1 => n21938, B2 => 
                           n16549, ZN => n5890);
   U14259 : OAI22_X1 port map( A1 => n21940, A2 => n22415, B1 => n21938, B2 => 
                           n16548, ZN => n5891);
   U14260 : OAI22_X1 port map( A1 => n21940, A2 => n22421, B1 => n21938, B2 => 
                           n16547, ZN => n5892);
   U14261 : OAI22_X1 port map( A1 => n21940, A2 => n22427, B1 => n21938, B2 => 
                           n16546, ZN => n5893);
   U14262 : OAI22_X1 port map( A1 => n21940, A2 => n22433, B1 => n21938, B2 => 
                           n16545, ZN => n5894);
   U14263 : OAI22_X1 port map( A1 => n21940, A2 => n22439, B1 => n21938, B2 => 
                           n16544, ZN => n5895);
   U14264 : OAI22_X1 port map( A1 => n21941, A2 => n22445, B1 => n21938, B2 => 
                           n16543, ZN => n5896);
   U14265 : OAI22_X1 port map( A1 => n21941, A2 => n22451, B1 => n21938, B2 => 
                           n16542, ZN => n5897);
   U14266 : OAI22_X1 port map( A1 => n21941, A2 => n22457, B1 => n21938, B2 => 
                           n16541, ZN => n5898);
   U14267 : OAI22_X1 port map( A1 => n21941, A2 => n22463, B1 => n21938, B2 => 
                           n16540, ZN => n5899);
   U14268 : OAI22_X1 port map( A1 => n21941, A2 => n22469, B1 => n16521, B2 => 
                           n16539, ZN => n5900);
   U14269 : OAI22_X1 port map( A1 => n21942, A2 => n22475, B1 => n16521, B2 => 
                           n16538, ZN => n5901);
   U14270 : OAI22_X1 port map( A1 => n21942, A2 => n22481, B1 => n16521, B2 => 
                           n16537, ZN => n5902);
   U14271 : OAI22_X1 port map( A1 => n21942, A2 => n22487, B1 => n16521, B2 => 
                           n16536, ZN => n5903);
   U14272 : OAI22_X1 port map( A1 => n21942, A2 => n22493, B1 => n16521, B2 => 
                           n16535, ZN => n5904);
   U14273 : OAI22_X1 port map( A1 => n21942, A2 => n22499, B1 => n16521, B2 => 
                           n16534, ZN => n5905);
   U14274 : OAI22_X1 port map( A1 => n21943, A2 => n22505, B1 => n16521, B2 => 
                           n16533, ZN => n5906);
   U14275 : OAI22_X1 port map( A1 => n21943, A2 => n22511, B1 => n21938, B2 => 
                           n16532, ZN => n5907);
   U14276 : OAI22_X1 port map( A1 => n21943, A2 => n22517, B1 => n21938, B2 => 
                           n16531, ZN => n5908);
   U14277 : OAI22_X1 port map( A1 => n21943, A2 => n22523, B1 => n21938, B2 => 
                           n16530, ZN => n5909);
   U14278 : OAI22_X1 port map( A1 => n21948, A2 => n22382, B1 => n21947, B2 => 
                           n16519, ZN => n5918);
   U14279 : OAI22_X1 port map( A1 => n21948, A2 => n22390, B1 => n21947, B2 => 
                           n16518, ZN => n5919);
   U14280 : OAI22_X1 port map( A1 => n21948, A2 => n22396, B1 => n21947, B2 => 
                           n16517, ZN => n5920);
   U14281 : OAI22_X1 port map( A1 => n21948, A2 => n22402, B1 => n21947, B2 => 
                           n16516, ZN => n5921);
   U14282 : OAI22_X1 port map( A1 => n21948, A2 => n22408, B1 => n21947, B2 => 
                           n16515, ZN => n5922);
   U14283 : OAI22_X1 port map( A1 => n21949, A2 => n22414, B1 => n21947, B2 => 
                           n16514, ZN => n5923);
   U14284 : OAI22_X1 port map( A1 => n21949, A2 => n22420, B1 => n21947, B2 => 
                           n16513, ZN => n5924);
   U14285 : OAI22_X1 port map( A1 => n21949, A2 => n22426, B1 => n21947, B2 => 
                           n16512, ZN => n5925);
   U14286 : OAI22_X1 port map( A1 => n21949, A2 => n22432, B1 => n21947, B2 => 
                           n16511, ZN => n5926);
   U14287 : OAI22_X1 port map( A1 => n21949, A2 => n22438, B1 => n21947, B2 => 
                           n16510, ZN => n5927);
   U14288 : OAI22_X1 port map( A1 => n21950, A2 => n22444, B1 => n21947, B2 => 
                           n16509, ZN => n5928);
   U14289 : OAI22_X1 port map( A1 => n21950, A2 => n22450, B1 => n21947, B2 => 
                           n16508, ZN => n5929);
   U14290 : OAI22_X1 port map( A1 => n21950, A2 => n22456, B1 => n21947, B2 => 
                           n16507, ZN => n5930);
   U14291 : OAI22_X1 port map( A1 => n21950, A2 => n22462, B1 => n21947, B2 => 
                           n16506, ZN => n5931);
   U14292 : OAI22_X1 port map( A1 => n21950, A2 => n22468, B1 => n16487, B2 => 
                           n16505, ZN => n5932);
   U14293 : OAI22_X1 port map( A1 => n21951, A2 => n22474, B1 => n16487, B2 => 
                           n16504, ZN => n5933);
   U14294 : OAI22_X1 port map( A1 => n21951, A2 => n22480, B1 => n16487, B2 => 
                           n16503, ZN => n5934);
   U14295 : OAI22_X1 port map( A1 => n21951, A2 => n22486, B1 => n16487, B2 => 
                           n16502, ZN => n5935);
   U14296 : OAI22_X1 port map( A1 => n21951, A2 => n22492, B1 => n16487, B2 => 
                           n16501, ZN => n5936);
   U14297 : OAI22_X1 port map( A1 => n21951, A2 => n22498, B1 => n16487, B2 => 
                           n16500, ZN => n5937);
   U14298 : OAI22_X1 port map( A1 => n21952, A2 => n22504, B1 => n16487, B2 => 
                           n16499, ZN => n5938);
   U14299 : OAI22_X1 port map( A1 => n21952, A2 => n22510, B1 => n21947, B2 => 
                           n16498, ZN => n5939);
   U14300 : OAI22_X1 port map( A1 => n21952, A2 => n22516, B1 => n21947, B2 => 
                           n16497, ZN => n5940);
   U14301 : OAI22_X1 port map( A1 => n21952, A2 => n22522, B1 => n21947, B2 => 
                           n16496, ZN => n5941);
   U14302 : OAI22_X1 port map( A1 => n21984, A2 => n22382, B1 => n21983, B2 => 
                           n16382, ZN => n6046);
   U14303 : OAI22_X1 port map( A1 => n21984, A2 => n22390, B1 => n21983, B2 => 
                           n16381, ZN => n6047);
   U14304 : OAI22_X1 port map( A1 => n21984, A2 => n22396, B1 => n21983, B2 => 
                           n16380, ZN => n6048);
   U14305 : OAI22_X1 port map( A1 => n21984, A2 => n22402, B1 => n21983, B2 => 
                           n16379, ZN => n6049);
   U14306 : OAI22_X1 port map( A1 => n21984, A2 => n22408, B1 => n21983, B2 => 
                           n16378, ZN => n6050);
   U14307 : OAI22_X1 port map( A1 => n21985, A2 => n22414, B1 => n21983, B2 => 
                           n16377, ZN => n6051);
   U14308 : OAI22_X1 port map( A1 => n21985, A2 => n22420, B1 => n21983, B2 => 
                           n16376, ZN => n6052);
   U14309 : OAI22_X1 port map( A1 => n21985, A2 => n22426, B1 => n21983, B2 => 
                           n16375, ZN => n6053);
   U14310 : OAI22_X1 port map( A1 => n21985, A2 => n22432, B1 => n21983, B2 => 
                           n16374, ZN => n6054);
   U14311 : OAI22_X1 port map( A1 => n21985, A2 => n22438, B1 => n21983, B2 => 
                           n16373, ZN => n6055);
   U14312 : OAI22_X1 port map( A1 => n21986, A2 => n22444, B1 => n21983, B2 => 
                           n16372, ZN => n6056);
   U14313 : OAI22_X1 port map( A1 => n21986, A2 => n22450, B1 => n21983, B2 => 
                           n16371, ZN => n6057);
   U14314 : OAI22_X1 port map( A1 => n21986, A2 => n22456, B1 => n21983, B2 => 
                           n16370, ZN => n6058);
   U14315 : OAI22_X1 port map( A1 => n21986, A2 => n22462, B1 => n21983, B2 => 
                           n16369, ZN => n6059);
   U14316 : OAI22_X1 port map( A1 => n21986, A2 => n22468, B1 => n16350, B2 => 
                           n16368, ZN => n6060);
   U14317 : OAI22_X1 port map( A1 => n21987, A2 => n22474, B1 => n16350, B2 => 
                           n16367, ZN => n6061);
   U14318 : OAI22_X1 port map( A1 => n21987, A2 => n22480, B1 => n16350, B2 => 
                           n16366, ZN => n6062);
   U14319 : OAI22_X1 port map( A1 => n21987, A2 => n22486, B1 => n16350, B2 => 
                           n16365, ZN => n6063);
   U14320 : OAI22_X1 port map( A1 => n21987, A2 => n22492, B1 => n16350, B2 => 
                           n16364, ZN => n6064);
   U14321 : OAI22_X1 port map( A1 => n21987, A2 => n22498, B1 => n16350, B2 => 
                           n16363, ZN => n6065);
   U14322 : OAI22_X1 port map( A1 => n21988, A2 => n22504, B1 => n16350, B2 => 
                           n16362, ZN => n6066);
   U14323 : OAI22_X1 port map( A1 => n21988, A2 => n22510, B1 => n21983, B2 => 
                           n16361, ZN => n6067);
   U14324 : OAI22_X1 port map( A1 => n21988, A2 => n22516, B1 => n21983, B2 => 
                           n16360, ZN => n6068);
   U14325 : OAI22_X1 port map( A1 => n21988, A2 => n22522, B1 => n21983, B2 => 
                           n16359, ZN => n6069);
   U14326 : OAI22_X1 port map( A1 => n22020, A2 => n22383, B1 => n22019, B2 => 
                           n16341, ZN => n6174);
   U14327 : OAI22_X1 port map( A1 => n22020, A2 => n22390, B1 => n22019, B2 => 
                           n16340, ZN => n6175);
   U14328 : OAI22_X1 port map( A1 => n22020, A2 => n22396, B1 => n22019, B2 => 
                           n16339, ZN => n6176);
   U14329 : OAI22_X1 port map( A1 => n22020, A2 => n22402, B1 => n22019, B2 => 
                           n16338, ZN => n6177);
   U14330 : OAI22_X1 port map( A1 => n22020, A2 => n22408, B1 => n22019, B2 => 
                           n16337, ZN => n6178);
   U14331 : OAI22_X1 port map( A1 => n22021, A2 => n22414, B1 => n22019, B2 => 
                           n16336, ZN => n6179);
   U14332 : OAI22_X1 port map( A1 => n22021, A2 => n22420, B1 => n22019, B2 => 
                           n16335, ZN => n6180);
   U14333 : OAI22_X1 port map( A1 => n22021, A2 => n22426, B1 => n22019, B2 => 
                           n16334, ZN => n6181);
   U14334 : OAI22_X1 port map( A1 => n22021, A2 => n22432, B1 => n22019, B2 => 
                           n16333, ZN => n6182);
   U14335 : OAI22_X1 port map( A1 => n22021, A2 => n22438, B1 => n22019, B2 => 
                           n16332, ZN => n6183);
   U14336 : OAI22_X1 port map( A1 => n22022, A2 => n22444, B1 => n22019, B2 => 
                           n16331, ZN => n6184);
   U14337 : OAI22_X1 port map( A1 => n22022, A2 => n22450, B1 => n22019, B2 => 
                           n16330, ZN => n6185);
   U14338 : OAI22_X1 port map( A1 => n22022, A2 => n22456, B1 => n22019, B2 => 
                           n16329, ZN => n6186);
   U14339 : OAI22_X1 port map( A1 => n22022, A2 => n22462, B1 => n22019, B2 => 
                           n16328, ZN => n6187);
   U14340 : OAI22_X1 port map( A1 => n22022, A2 => n22468, B1 => n16309, B2 => 
                           n16327, ZN => n6188);
   U14341 : OAI22_X1 port map( A1 => n22023, A2 => n22474, B1 => n16309, B2 => 
                           n16326, ZN => n6189);
   U14342 : OAI22_X1 port map( A1 => n22023, A2 => n22480, B1 => n16309, B2 => 
                           n16325, ZN => n6190);
   U14343 : OAI22_X1 port map( A1 => n22023, A2 => n22486, B1 => n16309, B2 => 
                           n16324, ZN => n6191);
   U14344 : OAI22_X1 port map( A1 => n22023, A2 => n22492, B1 => n16309, B2 => 
                           n16323, ZN => n6192);
   U14345 : OAI22_X1 port map( A1 => n22023, A2 => n22498, B1 => n16309, B2 => 
                           n16322, ZN => n6193);
   U14346 : OAI22_X1 port map( A1 => n22024, A2 => n22504, B1 => n16309, B2 => 
                           n16321, ZN => n6194);
   U14347 : OAI22_X1 port map( A1 => n22024, A2 => n22510, B1 => n22019, B2 => 
                           n16320, ZN => n6195);
   U14348 : OAI22_X1 port map( A1 => n22024, A2 => n22516, B1 => n22019, B2 => 
                           n16319, ZN => n6196);
   U14349 : OAI22_X1 port map( A1 => n22024, A2 => n22522, B1 => n22019, B2 => 
                           n16318, ZN => n6197);
   U14350 : OAI22_X1 port map( A1 => n22038, A2 => n22383, B1 => n22037, B2 => 
                           n16273, ZN => n6238);
   U14351 : OAI22_X1 port map( A1 => n22038, A2 => n22390, B1 => n22037, B2 => 
                           n16272, ZN => n6239);
   U14352 : OAI22_X1 port map( A1 => n22038, A2 => n22396, B1 => n22037, B2 => 
                           n16271, ZN => n6240);
   U14353 : OAI22_X1 port map( A1 => n22038, A2 => n22402, B1 => n22037, B2 => 
                           n16270, ZN => n6241);
   U14354 : OAI22_X1 port map( A1 => n22038, A2 => n22408, B1 => n22037, B2 => 
                           n16269, ZN => n6242);
   U14355 : OAI22_X1 port map( A1 => n22039, A2 => n22414, B1 => n22037, B2 => 
                           n16268, ZN => n6243);
   U14356 : OAI22_X1 port map( A1 => n22039, A2 => n22420, B1 => n22037, B2 => 
                           n16267, ZN => n6244);
   U14357 : OAI22_X1 port map( A1 => n22039, A2 => n22426, B1 => n22037, B2 => 
                           n16266, ZN => n6245);
   U14358 : OAI22_X1 port map( A1 => n22039, A2 => n22432, B1 => n22037, B2 => 
                           n16265, ZN => n6246);
   U14359 : OAI22_X1 port map( A1 => n22039, A2 => n22438, B1 => n22037, B2 => 
                           n16264, ZN => n6247);
   U14360 : OAI22_X1 port map( A1 => n22040, A2 => n22444, B1 => n22037, B2 => 
                           n16263, ZN => n6248);
   U14361 : OAI22_X1 port map( A1 => n22040, A2 => n22450, B1 => n22037, B2 => 
                           n16262, ZN => n6249);
   U14362 : OAI22_X1 port map( A1 => n22040, A2 => n22456, B1 => n22037, B2 => 
                           n16261, ZN => n6250);
   U14363 : OAI22_X1 port map( A1 => n22040, A2 => n22462, B1 => n22037, B2 => 
                           n16260, ZN => n6251);
   U14364 : OAI22_X1 port map( A1 => n22040, A2 => n22468, B1 => n16241, B2 => 
                           n16259, ZN => n6252);
   U14365 : OAI22_X1 port map( A1 => n22041, A2 => n22474, B1 => n16241, B2 => 
                           n16258, ZN => n6253);
   U14366 : OAI22_X1 port map( A1 => n22041, A2 => n22480, B1 => n16241, B2 => 
                           n16257, ZN => n6254);
   U14367 : OAI22_X1 port map( A1 => n22041, A2 => n22486, B1 => n16241, B2 => 
                           n16256, ZN => n6255);
   U14368 : OAI22_X1 port map( A1 => n22041, A2 => n22492, B1 => n16241, B2 => 
                           n16255, ZN => n6256);
   U14369 : OAI22_X1 port map( A1 => n22041, A2 => n22498, B1 => n16241, B2 => 
                           n16254, ZN => n6257);
   U14370 : OAI22_X1 port map( A1 => n22042, A2 => n22504, B1 => n16241, B2 => 
                           n16253, ZN => n6258);
   U14371 : OAI22_X1 port map( A1 => n22042, A2 => n22510, B1 => n22037, B2 => 
                           n16252, ZN => n6259);
   U14372 : OAI22_X1 port map( A1 => n22042, A2 => n22516, B1 => n22037, B2 => 
                           n16251, ZN => n6260);
   U14373 : OAI22_X1 port map( A1 => n22042, A2 => n22522, B1 => n22037, B2 => 
                           n16250, ZN => n6261);
   U14374 : OAI22_X1 port map( A1 => n22047, A2 => n22383, B1 => n22046, B2 => 
                           n16238, ZN => n6270);
   U14375 : OAI22_X1 port map( A1 => n22047, A2 => n22390, B1 => n22046, B2 => 
                           n16237, ZN => n6271);
   U14376 : OAI22_X1 port map( A1 => n22047, A2 => n22396, B1 => n22046, B2 => 
                           n16236, ZN => n6272);
   U14377 : OAI22_X1 port map( A1 => n22047, A2 => n22402, B1 => n22046, B2 => 
                           n16235, ZN => n6273);
   U14378 : OAI22_X1 port map( A1 => n22047, A2 => n22408, B1 => n22046, B2 => 
                           n16234, ZN => n6274);
   U14379 : OAI22_X1 port map( A1 => n22048, A2 => n22414, B1 => n22046, B2 => 
                           n16233, ZN => n6275);
   U14380 : OAI22_X1 port map( A1 => n22048, A2 => n22420, B1 => n22046, B2 => 
                           n16232, ZN => n6276);
   U14381 : OAI22_X1 port map( A1 => n22048, A2 => n22426, B1 => n22046, B2 => 
                           n16231, ZN => n6277);
   U14382 : OAI22_X1 port map( A1 => n22048, A2 => n22432, B1 => n22046, B2 => 
                           n16230, ZN => n6278);
   U14383 : OAI22_X1 port map( A1 => n22048, A2 => n22438, B1 => n22046, B2 => 
                           n16229, ZN => n6279);
   U14384 : OAI22_X1 port map( A1 => n22049, A2 => n22444, B1 => n22046, B2 => 
                           n16228, ZN => n6280);
   U14385 : OAI22_X1 port map( A1 => n22049, A2 => n22450, B1 => n22046, B2 => 
                           n16227, ZN => n6281);
   U14386 : OAI22_X1 port map( A1 => n22049, A2 => n22456, B1 => n22046, B2 => 
                           n16226, ZN => n6282);
   U14387 : OAI22_X1 port map( A1 => n22049, A2 => n22462, B1 => n22046, B2 => 
                           n16225, ZN => n6283);
   U14388 : OAI22_X1 port map( A1 => n22049, A2 => n22468, B1 => n16206, B2 => 
                           n16224, ZN => n6284);
   U14389 : OAI22_X1 port map( A1 => n22050, A2 => n22474, B1 => n16206, B2 => 
                           n16223, ZN => n6285);
   U14390 : OAI22_X1 port map( A1 => n22050, A2 => n22480, B1 => n16206, B2 => 
                           n16222, ZN => n6286);
   U14391 : OAI22_X1 port map( A1 => n22050, A2 => n22486, B1 => n16206, B2 => 
                           n16221, ZN => n6287);
   U14392 : OAI22_X1 port map( A1 => n22050, A2 => n22492, B1 => n16206, B2 => 
                           n16220, ZN => n6288);
   U14393 : OAI22_X1 port map( A1 => n22050, A2 => n22498, B1 => n16206, B2 => 
                           n16219, ZN => n6289);
   U14394 : OAI22_X1 port map( A1 => n22051, A2 => n22504, B1 => n16206, B2 => 
                           n16218, ZN => n6290);
   U14395 : OAI22_X1 port map( A1 => n22051, A2 => n22510, B1 => n22046, B2 => 
                           n16217, ZN => n6291);
   U14396 : OAI22_X1 port map( A1 => n22051, A2 => n22516, B1 => n22046, B2 => 
                           n16216, ZN => n6292);
   U14397 : OAI22_X1 port map( A1 => n22051, A2 => n22522, B1 => n22046, B2 => 
                           n16215, ZN => n6293);
   U14398 : OAI22_X1 port map( A1 => n22056, A2 => n22383, B1 => n22055, B2 => 
                           n16203, ZN => n6302);
   U14399 : OAI22_X1 port map( A1 => n22056, A2 => n22389, B1 => n22055, B2 => 
                           n16202, ZN => n6303);
   U14400 : OAI22_X1 port map( A1 => n22056, A2 => n22395, B1 => n22055, B2 => 
                           n16201, ZN => n6304);
   U14401 : OAI22_X1 port map( A1 => n22056, A2 => n22401, B1 => n22055, B2 => 
                           n16200, ZN => n6305);
   U14402 : OAI22_X1 port map( A1 => n22056, A2 => n22407, B1 => n22055, B2 => 
                           n16199, ZN => n6306);
   U14403 : OAI22_X1 port map( A1 => n22057, A2 => n22413, B1 => n22055, B2 => 
                           n16198, ZN => n6307);
   U14404 : OAI22_X1 port map( A1 => n22057, A2 => n22419, B1 => n22055, B2 => 
                           n16197, ZN => n6308);
   U14405 : OAI22_X1 port map( A1 => n22057, A2 => n22425, B1 => n22055, B2 => 
                           n16196, ZN => n6309);
   U14406 : OAI22_X1 port map( A1 => n22057, A2 => n22431, B1 => n22055, B2 => 
                           n16195, ZN => n6310);
   U14407 : OAI22_X1 port map( A1 => n22057, A2 => n22437, B1 => n22055, B2 => 
                           n16194, ZN => n6311);
   U14408 : OAI22_X1 port map( A1 => n22058, A2 => n22443, B1 => n22055, B2 => 
                           n16193, ZN => n6312);
   U14409 : OAI22_X1 port map( A1 => n22058, A2 => n22449, B1 => n22055, B2 => 
                           n16192, ZN => n6313);
   U14410 : OAI22_X1 port map( A1 => n22058, A2 => n22455, B1 => n22055, B2 => 
                           n16191, ZN => n6314);
   U14411 : OAI22_X1 port map( A1 => n22058, A2 => n22461, B1 => n22055, B2 => 
                           n16190, ZN => n6315);
   U14412 : OAI22_X1 port map( A1 => n22058, A2 => n22467, B1 => n16171, B2 => 
                           n16189, ZN => n6316);
   U14413 : OAI22_X1 port map( A1 => n22059, A2 => n22473, B1 => n16171, B2 => 
                           n16188, ZN => n6317);
   U14414 : OAI22_X1 port map( A1 => n22059, A2 => n22479, B1 => n16171, B2 => 
                           n16187, ZN => n6318);
   U14415 : OAI22_X1 port map( A1 => n22059, A2 => n22485, B1 => n16171, B2 => 
                           n16186, ZN => n6319);
   U14416 : OAI22_X1 port map( A1 => n22059, A2 => n22491, B1 => n16171, B2 => 
                           n16185, ZN => n6320);
   U14417 : OAI22_X1 port map( A1 => n22059, A2 => n22497, B1 => n16171, B2 => 
                           n16184, ZN => n6321);
   U14418 : OAI22_X1 port map( A1 => n22060, A2 => n22503, B1 => n16171, B2 => 
                           n16183, ZN => n6322);
   U14419 : OAI22_X1 port map( A1 => n22060, A2 => n22509, B1 => n22055, B2 => 
                           n16182, ZN => n6323);
   U14420 : OAI22_X1 port map( A1 => n22060, A2 => n22515, B1 => n22055, B2 => 
                           n16181, ZN => n6324);
   U14421 : OAI22_X1 port map( A1 => n22060, A2 => n22521, B1 => n22055, B2 => 
                           n16180, ZN => n6325);
   U14422 : OAI22_X1 port map( A1 => n22074, A2 => n22383, B1 => n22073, B2 => 
                           n16167, ZN => n6366);
   U14423 : OAI22_X1 port map( A1 => n22074, A2 => n22389, B1 => n22073, B2 => 
                           n16166, ZN => n6367);
   U14424 : OAI22_X1 port map( A1 => n22074, A2 => n22395, B1 => n22073, B2 => 
                           n16165, ZN => n6368);
   U14425 : OAI22_X1 port map( A1 => n22074, A2 => n22401, B1 => n22073, B2 => 
                           n16164, ZN => n6369);
   U14426 : OAI22_X1 port map( A1 => n22074, A2 => n22407, B1 => n22073, B2 => 
                           n16163, ZN => n6370);
   U14427 : OAI22_X1 port map( A1 => n22075, A2 => n22413, B1 => n22073, B2 => 
                           n16162, ZN => n6371);
   U14428 : OAI22_X1 port map( A1 => n22075, A2 => n22419, B1 => n22073, B2 => 
                           n16161, ZN => n6372);
   U14429 : OAI22_X1 port map( A1 => n22075, A2 => n22425, B1 => n22073, B2 => 
                           n16160, ZN => n6373);
   U14430 : OAI22_X1 port map( A1 => n22075, A2 => n22431, B1 => n22073, B2 => 
                           n16159, ZN => n6374);
   U14431 : OAI22_X1 port map( A1 => n22075, A2 => n22437, B1 => n22073, B2 => 
                           n16158, ZN => n6375);
   U14432 : OAI22_X1 port map( A1 => n22076, A2 => n22443, B1 => n22073, B2 => 
                           n16157, ZN => n6376);
   U14433 : OAI22_X1 port map( A1 => n22076, A2 => n22449, B1 => n22073, B2 => 
                           n16156, ZN => n6377);
   U14434 : OAI22_X1 port map( A1 => n22076, A2 => n22455, B1 => n22073, B2 => 
                           n16155, ZN => n6378);
   U14435 : OAI22_X1 port map( A1 => n22076, A2 => n22461, B1 => n22073, B2 => 
                           n16154, ZN => n6379);
   U14436 : OAI22_X1 port map( A1 => n22076, A2 => n22467, B1 => n16135, B2 => 
                           n16153, ZN => n6380);
   U14437 : OAI22_X1 port map( A1 => n22077, A2 => n22473, B1 => n16135, B2 => 
                           n16152, ZN => n6381);
   U14438 : OAI22_X1 port map( A1 => n22077, A2 => n22479, B1 => n16135, B2 => 
                           n16151, ZN => n6382);
   U14439 : OAI22_X1 port map( A1 => n22077, A2 => n22485, B1 => n16135, B2 => 
                           n16150, ZN => n6383);
   U14440 : OAI22_X1 port map( A1 => n22077, A2 => n22491, B1 => n16135, B2 => 
                           n16149, ZN => n6384);
   U14441 : OAI22_X1 port map( A1 => n22077, A2 => n22497, B1 => n16135, B2 => 
                           n16148, ZN => n6385);
   U14442 : OAI22_X1 port map( A1 => n22078, A2 => n22503, B1 => n16135, B2 => 
                           n16147, ZN => n6386);
   U14443 : OAI22_X1 port map( A1 => n22078, A2 => n22509, B1 => n22073, B2 => 
                           n16146, ZN => n6387);
   U14444 : OAI22_X1 port map( A1 => n22078, A2 => n22515, B1 => n22073, B2 => 
                           n16145, ZN => n6388);
   U14445 : OAI22_X1 port map( A1 => n22078, A2 => n22521, B1 => n22073, B2 => 
                           n16144, ZN => n6389);
   U14446 : OAI22_X1 port map( A1 => n22083, A2 => n22383, B1 => n22082, B2 => 
                           n16132, ZN => n6398);
   U14447 : OAI22_X1 port map( A1 => n22083, A2 => n22389, B1 => n22082, B2 => 
                           n16131, ZN => n6399);
   U14448 : OAI22_X1 port map( A1 => n22083, A2 => n22395, B1 => n22082, B2 => 
                           n16130, ZN => n6400);
   U14449 : OAI22_X1 port map( A1 => n22083, A2 => n22401, B1 => n22082, B2 => 
                           n16129, ZN => n6401);
   U14450 : OAI22_X1 port map( A1 => n22083, A2 => n22407, B1 => n22082, B2 => 
                           n16128, ZN => n6402);
   U14451 : OAI22_X1 port map( A1 => n22084, A2 => n22413, B1 => n22082, B2 => 
                           n16127, ZN => n6403);
   U14452 : OAI22_X1 port map( A1 => n22084, A2 => n22419, B1 => n22082, B2 => 
                           n16126, ZN => n6404);
   U14453 : OAI22_X1 port map( A1 => n22084, A2 => n22425, B1 => n22082, B2 => 
                           n16125, ZN => n6405);
   U14454 : OAI22_X1 port map( A1 => n22084, A2 => n22431, B1 => n22082, B2 => 
                           n16124, ZN => n6406);
   U14455 : OAI22_X1 port map( A1 => n22084, A2 => n22437, B1 => n22082, B2 => 
                           n16123, ZN => n6407);
   U14456 : OAI22_X1 port map( A1 => n22085, A2 => n22443, B1 => n22082, B2 => 
                           n16122, ZN => n6408);
   U14457 : OAI22_X1 port map( A1 => n22085, A2 => n22449, B1 => n22082, B2 => 
                           n16121, ZN => n6409);
   U14458 : OAI22_X1 port map( A1 => n22085, A2 => n22455, B1 => n22082, B2 => 
                           n16120, ZN => n6410);
   U14459 : OAI22_X1 port map( A1 => n22085, A2 => n22461, B1 => n22082, B2 => 
                           n16119, ZN => n6411);
   U14460 : OAI22_X1 port map( A1 => n22085, A2 => n22467, B1 => n16100, B2 => 
                           n16118, ZN => n6412);
   U14461 : OAI22_X1 port map( A1 => n22086, A2 => n22473, B1 => n16100, B2 => 
                           n16117, ZN => n6413);
   U14462 : OAI22_X1 port map( A1 => n22086, A2 => n22479, B1 => n16100, B2 => 
                           n16116, ZN => n6414);
   U14463 : OAI22_X1 port map( A1 => n22086, A2 => n22485, B1 => n16100, B2 => 
                           n16115, ZN => n6415);
   U14464 : OAI22_X1 port map( A1 => n22086, A2 => n22491, B1 => n16100, B2 => 
                           n16114, ZN => n6416);
   U14465 : OAI22_X1 port map( A1 => n22086, A2 => n22497, B1 => n16100, B2 => 
                           n16113, ZN => n6417);
   U14466 : OAI22_X1 port map( A1 => n22087, A2 => n22503, B1 => n16100, B2 => 
                           n16112, ZN => n6418);
   U14467 : OAI22_X1 port map( A1 => n22087, A2 => n22509, B1 => n22082, B2 => 
                           n16111, ZN => n6419);
   U14468 : OAI22_X1 port map( A1 => n22087, A2 => n22515, B1 => n22082, B2 => 
                           n16110, ZN => n6420);
   U14469 : OAI22_X1 port map( A1 => n22087, A2 => n22521, B1 => n22082, B2 => 
                           n16109, ZN => n6421);
   U14470 : OAI22_X1 port map( A1 => n22092, A2 => n22383, B1 => n22091, B2 => 
                           n16098, ZN => n6430);
   U14471 : OAI22_X1 port map( A1 => n22092, A2 => n22389, B1 => n22091, B2 => 
                           n16097, ZN => n6431);
   U14472 : OAI22_X1 port map( A1 => n22092, A2 => n22395, B1 => n22091, B2 => 
                           n16096, ZN => n6432);
   U14473 : OAI22_X1 port map( A1 => n22092, A2 => n22401, B1 => n22091, B2 => 
                           n16095, ZN => n6433);
   U14474 : OAI22_X1 port map( A1 => n22092, A2 => n22407, B1 => n22091, B2 => 
                           n16094, ZN => n6434);
   U14475 : OAI22_X1 port map( A1 => n22093, A2 => n22413, B1 => n22091, B2 => 
                           n16093, ZN => n6435);
   U14476 : OAI22_X1 port map( A1 => n22093, A2 => n22419, B1 => n22091, B2 => 
                           n16092, ZN => n6436);
   U14477 : OAI22_X1 port map( A1 => n22093, A2 => n22425, B1 => n22091, B2 => 
                           n16091, ZN => n6437);
   U14478 : OAI22_X1 port map( A1 => n22093, A2 => n22431, B1 => n22091, B2 => 
                           n16090, ZN => n6438);
   U14479 : OAI22_X1 port map( A1 => n22093, A2 => n22437, B1 => n22091, B2 => 
                           n16089, ZN => n6439);
   U14480 : OAI22_X1 port map( A1 => n22094, A2 => n22443, B1 => n22091, B2 => 
                           n16088, ZN => n6440);
   U14481 : OAI22_X1 port map( A1 => n22094, A2 => n22449, B1 => n22091, B2 => 
                           n16087, ZN => n6441);
   U14482 : OAI22_X1 port map( A1 => n22094, A2 => n22455, B1 => n22091, B2 => 
                           n16086, ZN => n6442);
   U14483 : OAI22_X1 port map( A1 => n22094, A2 => n22461, B1 => n22091, B2 => 
                           n16085, ZN => n6443);
   U14484 : OAI22_X1 port map( A1 => n22094, A2 => n22467, B1 => n16066, B2 => 
                           n16084, ZN => n6444);
   U14485 : OAI22_X1 port map( A1 => n22095, A2 => n22473, B1 => n16066, B2 => 
                           n16083, ZN => n6445);
   U14486 : OAI22_X1 port map( A1 => n22095, A2 => n22479, B1 => n16066, B2 => 
                           n16082, ZN => n6446);
   U14487 : OAI22_X1 port map( A1 => n22095, A2 => n22485, B1 => n16066, B2 => 
                           n16081, ZN => n6447);
   U14488 : OAI22_X1 port map( A1 => n22095, A2 => n22491, B1 => n16066, B2 => 
                           n16080, ZN => n6448);
   U14489 : OAI22_X1 port map( A1 => n22095, A2 => n22497, B1 => n16066, B2 => 
                           n16079, ZN => n6449);
   U14490 : OAI22_X1 port map( A1 => n22096, A2 => n22503, B1 => n16066, B2 => 
                           n16078, ZN => n6450);
   U14491 : OAI22_X1 port map( A1 => n22096, A2 => n22509, B1 => n22091, B2 => 
                           n16077, ZN => n6451);
   U14492 : OAI22_X1 port map( A1 => n22096, A2 => n22515, B1 => n22091, B2 => 
                           n16076, ZN => n6452);
   U14493 : OAI22_X1 port map( A1 => n22096, A2 => n22521, B1 => n22091, B2 => 
                           n16075, ZN => n6453);
   U14494 : OAI22_X1 port map( A1 => n22101, A2 => n22383, B1 => n22100, B2 => 
                           n16064, ZN => n6462);
   U14495 : OAI22_X1 port map( A1 => n22101, A2 => n22389, B1 => n22100, B2 => 
                           n16063, ZN => n6463);
   U14496 : OAI22_X1 port map( A1 => n22101, A2 => n22395, B1 => n22100, B2 => 
                           n16062, ZN => n6464);
   U14497 : OAI22_X1 port map( A1 => n22101, A2 => n22401, B1 => n22100, B2 => 
                           n16061, ZN => n6465);
   U14498 : OAI22_X1 port map( A1 => n22101, A2 => n22407, B1 => n22100, B2 => 
                           n16060, ZN => n6466);
   U14499 : OAI22_X1 port map( A1 => n22102, A2 => n22413, B1 => n22100, B2 => 
                           n16059, ZN => n6467);
   U14500 : OAI22_X1 port map( A1 => n22102, A2 => n22419, B1 => n22100, B2 => 
                           n16058, ZN => n6468);
   U14501 : OAI22_X1 port map( A1 => n22102, A2 => n22425, B1 => n22100, B2 => 
                           n16057, ZN => n6469);
   U14502 : OAI22_X1 port map( A1 => n22102, A2 => n22431, B1 => n22100, B2 => 
                           n16056, ZN => n6470);
   U14503 : OAI22_X1 port map( A1 => n22102, A2 => n22437, B1 => n22100, B2 => 
                           n16055, ZN => n6471);
   U14504 : OAI22_X1 port map( A1 => n22103, A2 => n22443, B1 => n22100, B2 => 
                           n16054, ZN => n6472);
   U14505 : OAI22_X1 port map( A1 => n22103, A2 => n22449, B1 => n22100, B2 => 
                           n16053, ZN => n6473);
   U14506 : OAI22_X1 port map( A1 => n22103, A2 => n22455, B1 => n22100, B2 => 
                           n16052, ZN => n6474);
   U14507 : OAI22_X1 port map( A1 => n22103, A2 => n22461, B1 => n22100, B2 => 
                           n16051, ZN => n6475);
   U14508 : OAI22_X1 port map( A1 => n22103, A2 => n22467, B1 => n16032, B2 => 
                           n16050, ZN => n6476);
   U14509 : OAI22_X1 port map( A1 => n22104, A2 => n22473, B1 => n16032, B2 => 
                           n16049, ZN => n6477);
   U14510 : OAI22_X1 port map( A1 => n22104, A2 => n22479, B1 => n16032, B2 => 
                           n16048, ZN => n6478);
   U14511 : OAI22_X1 port map( A1 => n22104, A2 => n22485, B1 => n16032, B2 => 
                           n16047, ZN => n6479);
   U14512 : OAI22_X1 port map( A1 => n22104, A2 => n22491, B1 => n16032, B2 => 
                           n16046, ZN => n6480);
   U14513 : OAI22_X1 port map( A1 => n22104, A2 => n22497, B1 => n16032, B2 => 
                           n16045, ZN => n6481);
   U14514 : OAI22_X1 port map( A1 => n22105, A2 => n22503, B1 => n16032, B2 => 
                           n16044, ZN => n6482);
   U14515 : OAI22_X1 port map( A1 => n22105, A2 => n22509, B1 => n22100, B2 => 
                           n16043, ZN => n6483);
   U14516 : OAI22_X1 port map( A1 => n22105, A2 => n22515, B1 => n22100, B2 => 
                           n16042, ZN => n6484);
   U14517 : OAI22_X1 port map( A1 => n22105, A2 => n22521, B1 => n22100, B2 => 
                           n16041, ZN => n6485);
   U14518 : OAI22_X1 port map( A1 => n22137, A2 => n22384, B1 => n22136, B2 => 
                           n15927, ZN => n6590);
   U14519 : OAI22_X1 port map( A1 => n22137, A2 => n22389, B1 => n22136, B2 => 
                           n15926, ZN => n6591);
   U14520 : OAI22_X1 port map( A1 => n22137, A2 => n22395, B1 => n22136, B2 => 
                           n15925, ZN => n6592);
   U14521 : OAI22_X1 port map( A1 => n22137, A2 => n22401, B1 => n22136, B2 => 
                           n15924, ZN => n6593);
   U14522 : OAI22_X1 port map( A1 => n22137, A2 => n22407, B1 => n22136, B2 => 
                           n15923, ZN => n6594);
   U14523 : OAI22_X1 port map( A1 => n22138, A2 => n22413, B1 => n22136, B2 => 
                           n15922, ZN => n6595);
   U14524 : OAI22_X1 port map( A1 => n22138, A2 => n22419, B1 => n22136, B2 => 
                           n15921, ZN => n6596);
   U14525 : OAI22_X1 port map( A1 => n22138, A2 => n22425, B1 => n22136, B2 => 
                           n15920, ZN => n6597);
   U14526 : OAI22_X1 port map( A1 => n22138, A2 => n22431, B1 => n22136, B2 => 
                           n15919, ZN => n6598);
   U14527 : OAI22_X1 port map( A1 => n22138, A2 => n22437, B1 => n22136, B2 => 
                           n15918, ZN => n6599);
   U14528 : OAI22_X1 port map( A1 => n22139, A2 => n22443, B1 => n22136, B2 => 
                           n15917, ZN => n6600);
   U14529 : OAI22_X1 port map( A1 => n22139, A2 => n22449, B1 => n22136, B2 => 
                           n15916, ZN => n6601);
   U14530 : OAI22_X1 port map( A1 => n22139, A2 => n22455, B1 => n22136, B2 => 
                           n15915, ZN => n6602);
   U14531 : OAI22_X1 port map( A1 => n22139, A2 => n22461, B1 => n22136, B2 => 
                           n15914, ZN => n6603);
   U14532 : OAI22_X1 port map( A1 => n22139, A2 => n22467, B1 => n15895, B2 => 
                           n15913, ZN => n6604);
   U14533 : OAI22_X1 port map( A1 => n22140, A2 => n22473, B1 => n15895, B2 => 
                           n15912, ZN => n6605);
   U14534 : OAI22_X1 port map( A1 => n22140, A2 => n22479, B1 => n15895, B2 => 
                           n15911, ZN => n6606);
   U14535 : OAI22_X1 port map( A1 => n22140, A2 => n22485, B1 => n15895, B2 => 
                           n15910, ZN => n6607);
   U14536 : OAI22_X1 port map( A1 => n22140, A2 => n22491, B1 => n15895, B2 => 
                           n15909, ZN => n6608);
   U14537 : OAI22_X1 port map( A1 => n22140, A2 => n22497, B1 => n15895, B2 => 
                           n15908, ZN => n6609);
   U14538 : OAI22_X1 port map( A1 => n22141, A2 => n22503, B1 => n15895, B2 => 
                           n15907, ZN => n6610);
   U14539 : OAI22_X1 port map( A1 => n22141, A2 => n22509, B1 => n22136, B2 => 
                           n15906, ZN => n6611);
   U14540 : OAI22_X1 port map( A1 => n22141, A2 => n22515, B1 => n22136, B2 => 
                           n15905, ZN => n6612);
   U14541 : OAI22_X1 port map( A1 => n22141, A2 => n22521, B1 => n22136, B2 => 
                           n15904, ZN => n6613);
   U14542 : OAI22_X1 port map( A1 => n22173, A2 => n22384, B1 => n22172, B2 => 
                           n15854, ZN => n6718);
   U14543 : OAI22_X1 port map( A1 => n22173, A2 => n22388, B1 => n22172, B2 => 
                           n15853, ZN => n6719);
   U14544 : OAI22_X1 port map( A1 => n22173, A2 => n22394, B1 => n22172, B2 => 
                           n15852, ZN => n6720);
   U14545 : OAI22_X1 port map( A1 => n22173, A2 => n22400, B1 => n22172, B2 => 
                           n15851, ZN => n6721);
   U14546 : OAI22_X1 port map( A1 => n22173, A2 => n22406, B1 => n22172, B2 => 
                           n15850, ZN => n6722);
   U14547 : OAI22_X1 port map( A1 => n22174, A2 => n22412, B1 => n22172, B2 => 
                           n15849, ZN => n6723);
   U14548 : OAI22_X1 port map( A1 => n22174, A2 => n22418, B1 => n22172, B2 => 
                           n15848, ZN => n6724);
   U14549 : OAI22_X1 port map( A1 => n22174, A2 => n22424, B1 => n22172, B2 => 
                           n15847, ZN => n6725);
   U14550 : OAI22_X1 port map( A1 => n22174, A2 => n22430, B1 => n22172, B2 => 
                           n15846, ZN => n6726);
   U14551 : OAI22_X1 port map( A1 => n22174, A2 => n22436, B1 => n22172, B2 => 
                           n15845, ZN => n6727);
   U14552 : OAI22_X1 port map( A1 => n22175, A2 => n22442, B1 => n22172, B2 => 
                           n15844, ZN => n6728);
   U14553 : OAI22_X1 port map( A1 => n22175, A2 => n22448, B1 => n22172, B2 => 
                           n15843, ZN => n6729);
   U14554 : OAI22_X1 port map( A1 => n22175, A2 => n22454, B1 => n22172, B2 => 
                           n15842, ZN => n6730);
   U14555 : OAI22_X1 port map( A1 => n22175, A2 => n22460, B1 => n22172, B2 => 
                           n15841, ZN => n6731);
   U14556 : OAI22_X1 port map( A1 => n22175, A2 => n22466, B1 => n15822, B2 => 
                           n15840, ZN => n6732);
   U14557 : OAI22_X1 port map( A1 => n22176, A2 => n22472, B1 => n15822, B2 => 
                           n15839, ZN => n6733);
   U14558 : OAI22_X1 port map( A1 => n22176, A2 => n22478, B1 => n15822, B2 => 
                           n15838, ZN => n6734);
   U14559 : OAI22_X1 port map( A1 => n22176, A2 => n22484, B1 => n15822, B2 => 
                           n15837, ZN => n6735);
   U14560 : OAI22_X1 port map( A1 => n22176, A2 => n22490, B1 => n15822, B2 => 
                           n15836, ZN => n6736);
   U14561 : OAI22_X1 port map( A1 => n22176, A2 => n22496, B1 => n15822, B2 => 
                           n15835, ZN => n6737);
   U14562 : OAI22_X1 port map( A1 => n22177, A2 => n22502, B1 => n15822, B2 => 
                           n15834, ZN => n6738);
   U14563 : OAI22_X1 port map( A1 => n22177, A2 => n22508, B1 => n22172, B2 => 
                           n15833, ZN => n6739);
   U14564 : OAI22_X1 port map( A1 => n22177, A2 => n22514, B1 => n22172, B2 => 
                           n15832, ZN => n6740);
   U14565 : OAI22_X1 port map( A1 => n22177, A2 => n22520, B1 => n22172, B2 => 
                           n15831, ZN => n6741);
   U14566 : OAI22_X1 port map( A1 => n22182, A2 => n22384, B1 => n22181, B2 => 
                           n15820, ZN => n6750);
   U14567 : OAI22_X1 port map( A1 => n22182, A2 => n22388, B1 => n22181, B2 => 
                           n15819, ZN => n6751);
   U14568 : OAI22_X1 port map( A1 => n22182, A2 => n22394, B1 => n22181, B2 => 
                           n15818, ZN => n6752);
   U14569 : OAI22_X1 port map( A1 => n22182, A2 => n22400, B1 => n22181, B2 => 
                           n15817, ZN => n6753);
   U14570 : OAI22_X1 port map( A1 => n22182, A2 => n22406, B1 => n22181, B2 => 
                           n15816, ZN => n6754);
   U14571 : OAI22_X1 port map( A1 => n22183, A2 => n22412, B1 => n22181, B2 => 
                           n15815, ZN => n6755);
   U14572 : OAI22_X1 port map( A1 => n22183, A2 => n22418, B1 => n22181, B2 => 
                           n15814, ZN => n6756);
   U14573 : OAI22_X1 port map( A1 => n22183, A2 => n22424, B1 => n22181, B2 => 
                           n15813, ZN => n6757);
   U14574 : OAI22_X1 port map( A1 => n22183, A2 => n22430, B1 => n22181, B2 => 
                           n15812, ZN => n6758);
   U14575 : OAI22_X1 port map( A1 => n22183, A2 => n22436, B1 => n22181, B2 => 
                           n15811, ZN => n6759);
   U14576 : OAI22_X1 port map( A1 => n22184, A2 => n22442, B1 => n22181, B2 => 
                           n15810, ZN => n6760);
   U14577 : OAI22_X1 port map( A1 => n22184, A2 => n22448, B1 => n22181, B2 => 
                           n15809, ZN => n6761);
   U14578 : OAI22_X1 port map( A1 => n22184, A2 => n22454, B1 => n22181, B2 => 
                           n15808, ZN => n6762);
   U14579 : OAI22_X1 port map( A1 => n22184, A2 => n22460, B1 => n22181, B2 => 
                           n15807, ZN => n6763);
   U14580 : OAI22_X1 port map( A1 => n22184, A2 => n22466, B1 => n15788, B2 => 
                           n15806, ZN => n6764);
   U14581 : OAI22_X1 port map( A1 => n22185, A2 => n22472, B1 => n15788, B2 => 
                           n15805, ZN => n6765);
   U14582 : OAI22_X1 port map( A1 => n22185, A2 => n22478, B1 => n15788, B2 => 
                           n15804, ZN => n6766);
   U14583 : OAI22_X1 port map( A1 => n22185, A2 => n22484, B1 => n15788, B2 => 
                           n15803, ZN => n6767);
   U14584 : OAI22_X1 port map( A1 => n22185, A2 => n22490, B1 => n15788, B2 => 
                           n15802, ZN => n6768);
   U14585 : OAI22_X1 port map( A1 => n22185, A2 => n22496, B1 => n15788, B2 => 
                           n15801, ZN => n6769);
   U14586 : OAI22_X1 port map( A1 => n22186, A2 => n22502, B1 => n15788, B2 => 
                           n15800, ZN => n6770);
   U14587 : OAI22_X1 port map( A1 => n22186, A2 => n22508, B1 => n22181, B2 => 
                           n15799, ZN => n6771);
   U14588 : OAI22_X1 port map( A1 => n22186, A2 => n22514, B1 => n22181, B2 => 
                           n15798, ZN => n6772);
   U14589 : OAI22_X1 port map( A1 => n22186, A2 => n22520, B1 => n22181, B2 => 
                           n15797, ZN => n6773);
   U14590 : OAI22_X1 port map( A1 => n22191, A2 => n22384, B1 => n22190, B2 => 
                           n15785, ZN => n6782);
   U14591 : OAI22_X1 port map( A1 => n22191, A2 => n22388, B1 => n22190, B2 => 
                           n15784, ZN => n6783);
   U14592 : OAI22_X1 port map( A1 => n22191, A2 => n22394, B1 => n22190, B2 => 
                           n15783, ZN => n6784);
   U14593 : OAI22_X1 port map( A1 => n22191, A2 => n22400, B1 => n22190, B2 => 
                           n15782, ZN => n6785);
   U14594 : OAI22_X1 port map( A1 => n22191, A2 => n22406, B1 => n22190, B2 => 
                           n15781, ZN => n6786);
   U14595 : OAI22_X1 port map( A1 => n22192, A2 => n22412, B1 => n22190, B2 => 
                           n15780, ZN => n6787);
   U14596 : OAI22_X1 port map( A1 => n22192, A2 => n22418, B1 => n22190, B2 => 
                           n15779, ZN => n6788);
   U14597 : OAI22_X1 port map( A1 => n22192, A2 => n22424, B1 => n22190, B2 => 
                           n15778, ZN => n6789);
   U14598 : OAI22_X1 port map( A1 => n22192, A2 => n22430, B1 => n22190, B2 => 
                           n15777, ZN => n6790);
   U14599 : OAI22_X1 port map( A1 => n22192, A2 => n22436, B1 => n22190, B2 => 
                           n15776, ZN => n6791);
   U14600 : OAI22_X1 port map( A1 => n22193, A2 => n22442, B1 => n22190, B2 => 
                           n15775, ZN => n6792);
   U14601 : OAI22_X1 port map( A1 => n22193, A2 => n22448, B1 => n22190, B2 => 
                           n15774, ZN => n6793);
   U14602 : OAI22_X1 port map( A1 => n22193, A2 => n22454, B1 => n22190, B2 => 
                           n15773, ZN => n6794);
   U14603 : OAI22_X1 port map( A1 => n22193, A2 => n22460, B1 => n22190, B2 => 
                           n15772, ZN => n6795);
   U14604 : OAI22_X1 port map( A1 => n22193, A2 => n22466, B1 => n15753, B2 => 
                           n15771, ZN => n6796);
   U14605 : OAI22_X1 port map( A1 => n22194, A2 => n22472, B1 => n15753, B2 => 
                           n15770, ZN => n6797);
   U14606 : OAI22_X1 port map( A1 => n22194, A2 => n22478, B1 => n15753, B2 => 
                           n15769, ZN => n6798);
   U14607 : OAI22_X1 port map( A1 => n22194, A2 => n22484, B1 => n15753, B2 => 
                           n15768, ZN => n6799);
   U14608 : OAI22_X1 port map( A1 => n22194, A2 => n22490, B1 => n15753, B2 => 
                           n15767, ZN => n6800);
   U14609 : OAI22_X1 port map( A1 => n22194, A2 => n22496, B1 => n15753, B2 => 
                           n15766, ZN => n6801);
   U14610 : OAI22_X1 port map( A1 => n22195, A2 => n22502, B1 => n15753, B2 => 
                           n15765, ZN => n6802);
   U14611 : OAI22_X1 port map( A1 => n22195, A2 => n22508, B1 => n22190, B2 => 
                           n15764, ZN => n6803);
   U14612 : OAI22_X1 port map( A1 => n22195, A2 => n22514, B1 => n22190, B2 => 
                           n15763, ZN => n6804);
   U14613 : OAI22_X1 port map( A1 => n22195, A2 => n22520, B1 => n22190, B2 => 
                           n15762, ZN => n6805);
   U14614 : OAI22_X1 port map( A1 => n22218, A2 => n22384, B1 => n22217, B2 => 
                           n15714, ZN => n6878);
   U14615 : OAI22_X1 port map( A1 => n22218, A2 => n22388, B1 => n22217, B2 => 
                           n15713, ZN => n6879);
   U14616 : OAI22_X1 port map( A1 => n22218, A2 => n22394, B1 => n22217, B2 => 
                           n15712, ZN => n6880);
   U14617 : OAI22_X1 port map( A1 => n22218, A2 => n22400, B1 => n22217, B2 => 
                           n15711, ZN => n6881);
   U14618 : OAI22_X1 port map( A1 => n22218, A2 => n22406, B1 => n22217, B2 => 
                           n15710, ZN => n6882);
   U14619 : OAI22_X1 port map( A1 => n22219, A2 => n22412, B1 => n22217, B2 => 
                           n15709, ZN => n6883);
   U14620 : OAI22_X1 port map( A1 => n22219, A2 => n22418, B1 => n22217, B2 => 
                           n15708, ZN => n6884);
   U14621 : OAI22_X1 port map( A1 => n22219, A2 => n22424, B1 => n22217, B2 => 
                           n15707, ZN => n6885);
   U14622 : OAI22_X1 port map( A1 => n22219, A2 => n22430, B1 => n22217, B2 => 
                           n15706, ZN => n6886);
   U14623 : OAI22_X1 port map( A1 => n22219, A2 => n22436, B1 => n22217, B2 => 
                           n15705, ZN => n6887);
   U14624 : OAI22_X1 port map( A1 => n22220, A2 => n22442, B1 => n22217, B2 => 
                           n15704, ZN => n6888);
   U14625 : OAI22_X1 port map( A1 => n22220, A2 => n22448, B1 => n22217, B2 => 
                           n15703, ZN => n6889);
   U14626 : OAI22_X1 port map( A1 => n22220, A2 => n22454, B1 => n22217, B2 => 
                           n15702, ZN => n6890);
   U14627 : OAI22_X1 port map( A1 => n22220, A2 => n22460, B1 => n22217, B2 => 
                           n15701, ZN => n6891);
   U14628 : OAI22_X1 port map( A1 => n22220, A2 => n22466, B1 => n15682, B2 => 
                           n15700, ZN => n6892);
   U14629 : OAI22_X1 port map( A1 => n22221, A2 => n22472, B1 => n15682, B2 => 
                           n15699, ZN => n6893);
   U14630 : OAI22_X1 port map( A1 => n22221, A2 => n22478, B1 => n15682, B2 => 
                           n15698, ZN => n6894);
   U14631 : OAI22_X1 port map( A1 => n22221, A2 => n22484, B1 => n15682, B2 => 
                           n15697, ZN => n6895);
   U14632 : OAI22_X1 port map( A1 => n22221, A2 => n22490, B1 => n15682, B2 => 
                           n15696, ZN => n6896);
   U14633 : OAI22_X1 port map( A1 => n22221, A2 => n22496, B1 => n15682, B2 => 
                           n15695, ZN => n6897);
   U14634 : OAI22_X1 port map( A1 => n22222, A2 => n22502, B1 => n15682, B2 => 
                           n15694, ZN => n6898);
   U14635 : OAI22_X1 port map( A1 => n22222, A2 => n22508, B1 => n22217, B2 => 
                           n15693, ZN => n6899);
   U14636 : OAI22_X1 port map( A1 => n22222, A2 => n22514, B1 => n22217, B2 => 
                           n15692, ZN => n6900);
   U14637 : OAI22_X1 port map( A1 => n22222, A2 => n22520, B1 => n22217, B2 => 
                           n15691, ZN => n6901);
   U14638 : OAI22_X1 port map( A1 => n22227, A2 => n22384, B1 => n22226, B2 => 
                           n15679, ZN => n6910);
   U14639 : OAI22_X1 port map( A1 => n22227, A2 => n22388, B1 => n22226, B2 => 
                           n15678, ZN => n6911);
   U14640 : OAI22_X1 port map( A1 => n22227, A2 => n22394, B1 => n22226, B2 => 
                           n15677, ZN => n6912);
   U14641 : OAI22_X1 port map( A1 => n22227, A2 => n22400, B1 => n22226, B2 => 
                           n15676, ZN => n6913);
   U14642 : OAI22_X1 port map( A1 => n22227, A2 => n22406, B1 => n22226, B2 => 
                           n15675, ZN => n6914);
   U14643 : OAI22_X1 port map( A1 => n22228, A2 => n22412, B1 => n22226, B2 => 
                           n15674, ZN => n6915);
   U14644 : OAI22_X1 port map( A1 => n22228, A2 => n22418, B1 => n22226, B2 => 
                           n15673, ZN => n6916);
   U14645 : OAI22_X1 port map( A1 => n22228, A2 => n22424, B1 => n22226, B2 => 
                           n15672, ZN => n6917);
   U14646 : OAI22_X1 port map( A1 => n22228, A2 => n22430, B1 => n22226, B2 => 
                           n15671, ZN => n6918);
   U14647 : OAI22_X1 port map( A1 => n22228, A2 => n22436, B1 => n22226, B2 => 
                           n15670, ZN => n6919);
   U14648 : OAI22_X1 port map( A1 => n22229, A2 => n22442, B1 => n22226, B2 => 
                           n15669, ZN => n6920);
   U14649 : OAI22_X1 port map( A1 => n22229, A2 => n22448, B1 => n22226, B2 => 
                           n15668, ZN => n6921);
   U14650 : OAI22_X1 port map( A1 => n22229, A2 => n22454, B1 => n22226, B2 => 
                           n15667, ZN => n6922);
   U14651 : OAI22_X1 port map( A1 => n22229, A2 => n22460, B1 => n22226, B2 => 
                           n15666, ZN => n6923);
   U14652 : OAI22_X1 port map( A1 => n22229, A2 => n22466, B1 => n15647, B2 => 
                           n15665, ZN => n6924);
   U14653 : OAI22_X1 port map( A1 => n22230, A2 => n22472, B1 => n15647, B2 => 
                           n15664, ZN => n6925);
   U14654 : OAI22_X1 port map( A1 => n22230, A2 => n22478, B1 => n15647, B2 => 
                           n15663, ZN => n6926);
   U14655 : OAI22_X1 port map( A1 => n22230, A2 => n22484, B1 => n15647, B2 => 
                           n15662, ZN => n6927);
   U14656 : OAI22_X1 port map( A1 => n22230, A2 => n22490, B1 => n15647, B2 => 
                           n15661, ZN => n6928);
   U14657 : OAI22_X1 port map( A1 => n22230, A2 => n22496, B1 => n15647, B2 => 
                           n15660, ZN => n6929);
   U14658 : OAI22_X1 port map( A1 => n22231, A2 => n22502, B1 => n15647, B2 => 
                           n15659, ZN => n6930);
   U14659 : OAI22_X1 port map( A1 => n22231, A2 => n22508, B1 => n22226, B2 => 
                           n15658, ZN => n6931);
   U14660 : OAI22_X1 port map( A1 => n22231, A2 => n22514, B1 => n22226, B2 => 
                           n15657, ZN => n6932);
   U14661 : OAI22_X1 port map( A1 => n22231, A2 => n22520, B1 => n22226, B2 => 
                           n15656, ZN => n6933);
   U14662 : OAI22_X1 port map( A1 => n22245, A2 => n22385, B1 => n22244, B2 => 
                           n15607, ZN => n6974);
   U14663 : OAI22_X1 port map( A1 => n22245, A2 => n22388, B1 => n22244, B2 => 
                           n15606, ZN => n6975);
   U14664 : OAI22_X1 port map( A1 => n22245, A2 => n22394, B1 => n22244, B2 => 
                           n15605, ZN => n6976);
   U14665 : OAI22_X1 port map( A1 => n22245, A2 => n22400, B1 => n22244, B2 => 
                           n15604, ZN => n6977);
   U14666 : OAI22_X1 port map( A1 => n22245, A2 => n22406, B1 => n22244, B2 => 
                           n15603, ZN => n6978);
   U14667 : OAI22_X1 port map( A1 => n22246, A2 => n22412, B1 => n22244, B2 => 
                           n15602, ZN => n6979);
   U14668 : OAI22_X1 port map( A1 => n22246, A2 => n22418, B1 => n22244, B2 => 
                           n15601, ZN => n6980);
   U14669 : OAI22_X1 port map( A1 => n22246, A2 => n22424, B1 => n22244, B2 => 
                           n15600, ZN => n6981);
   U14670 : OAI22_X1 port map( A1 => n22246, A2 => n22430, B1 => n22244, B2 => 
                           n15599, ZN => n6982);
   U14671 : OAI22_X1 port map( A1 => n22246, A2 => n22436, B1 => n22244, B2 => 
                           n15598, ZN => n6983);
   U14672 : OAI22_X1 port map( A1 => n22247, A2 => n22442, B1 => n22244, B2 => 
                           n15597, ZN => n6984);
   U14673 : OAI22_X1 port map( A1 => n22247, A2 => n22448, B1 => n22244, B2 => 
                           n15596, ZN => n6985);
   U14674 : OAI22_X1 port map( A1 => n22247, A2 => n22454, B1 => n22244, B2 => 
                           n15595, ZN => n6986);
   U14675 : OAI22_X1 port map( A1 => n22247, A2 => n22460, B1 => n22244, B2 => 
                           n15594, ZN => n6987);
   U14676 : OAI22_X1 port map( A1 => n22247, A2 => n22466, B1 => n15575, B2 => 
                           n15593, ZN => n6988);
   U14677 : OAI22_X1 port map( A1 => n22248, A2 => n22472, B1 => n15575, B2 => 
                           n15592, ZN => n6989);
   U14678 : OAI22_X1 port map( A1 => n22248, A2 => n22478, B1 => n15575, B2 => 
                           n15591, ZN => n6990);
   U14679 : OAI22_X1 port map( A1 => n22248, A2 => n22484, B1 => n15575, B2 => 
                           n15590, ZN => n6991);
   U14680 : OAI22_X1 port map( A1 => n22248, A2 => n22490, B1 => n15575, B2 => 
                           n15589, ZN => n6992);
   U14681 : OAI22_X1 port map( A1 => n22248, A2 => n22496, B1 => n15575, B2 => 
                           n15588, ZN => n6993);
   U14682 : OAI22_X1 port map( A1 => n22249, A2 => n22502, B1 => n15575, B2 => 
                           n15587, ZN => n6994);
   U14683 : OAI22_X1 port map( A1 => n22249, A2 => n22508, B1 => n22244, B2 => 
                           n15586, ZN => n6995);
   U14684 : OAI22_X1 port map( A1 => n22249, A2 => n22514, B1 => n22244, B2 => 
                           n15585, ZN => n6996);
   U14685 : OAI22_X1 port map( A1 => n22249, A2 => n22520, B1 => n22244, B2 => 
                           n15584, ZN => n6997);
   U14686 : OAI22_X1 port map( A1 => n22272, A2 => n22385, B1 => n22271, B2 => 
                           n15503, ZN => n7070);
   U14687 : OAI22_X1 port map( A1 => n22272, A2 => n22387, B1 => n22271, B2 => 
                           n15502, ZN => n7071);
   U14688 : OAI22_X1 port map( A1 => n22272, A2 => n22393, B1 => n22271, B2 => 
                           n15501, ZN => n7072);
   U14689 : OAI22_X1 port map( A1 => n22272, A2 => n22399, B1 => n22271, B2 => 
                           n15500, ZN => n7073);
   U14690 : OAI22_X1 port map( A1 => n22272, A2 => n22405, B1 => n22271, B2 => 
                           n15499, ZN => n7074);
   U14691 : OAI22_X1 port map( A1 => n22273, A2 => n22411, B1 => n22271, B2 => 
                           n15498, ZN => n7075);
   U14692 : OAI22_X1 port map( A1 => n22273, A2 => n22417, B1 => n22271, B2 => 
                           n15497, ZN => n7076);
   U14693 : OAI22_X1 port map( A1 => n22273, A2 => n22423, B1 => n22271, B2 => 
                           n15496, ZN => n7077);
   U14694 : OAI22_X1 port map( A1 => n22273, A2 => n22429, B1 => n22271, B2 => 
                           n15495, ZN => n7078);
   U14695 : OAI22_X1 port map( A1 => n22273, A2 => n22435, B1 => n22271, B2 => 
                           n15494, ZN => n7079);
   U14696 : OAI22_X1 port map( A1 => n22274, A2 => n22441, B1 => n22271, B2 => 
                           n15493, ZN => n7080);
   U14697 : OAI22_X1 port map( A1 => n22274, A2 => n22447, B1 => n22271, B2 => 
                           n15492, ZN => n7081);
   U14698 : OAI22_X1 port map( A1 => n22274, A2 => n22453, B1 => n22271, B2 => 
                           n15491, ZN => n7082);
   U14699 : OAI22_X1 port map( A1 => n22274, A2 => n22459, B1 => n22271, B2 => 
                           n15490, ZN => n7083);
   U14700 : OAI22_X1 port map( A1 => n22274, A2 => n22465, B1 => n15471, B2 => 
                           n15489, ZN => n7084);
   U14701 : OAI22_X1 port map( A1 => n22275, A2 => n22471, B1 => n15471, B2 => 
                           n15488, ZN => n7085);
   U14702 : OAI22_X1 port map( A1 => n22275, A2 => n22477, B1 => n15471, B2 => 
                           n15487, ZN => n7086);
   U14703 : OAI22_X1 port map( A1 => n22275, A2 => n22483, B1 => n15471, B2 => 
                           n15486, ZN => n7087);
   U14704 : OAI22_X1 port map( A1 => n22275, A2 => n22489, B1 => n15471, B2 => 
                           n15485, ZN => n7088);
   U14705 : OAI22_X1 port map( A1 => n22275, A2 => n22495, B1 => n15471, B2 => 
                           n15484, ZN => n7089);
   U14706 : OAI22_X1 port map( A1 => n22276, A2 => n22501, B1 => n15471, B2 => 
                           n15483, ZN => n7090);
   U14707 : OAI22_X1 port map( A1 => n22276, A2 => n22507, B1 => n22271, B2 => 
                           n15482, ZN => n7091);
   U14708 : OAI22_X1 port map( A1 => n22276, A2 => n22513, B1 => n22271, B2 => 
                           n15481, ZN => n7092);
   U14709 : OAI22_X1 port map( A1 => n22276, A2 => n22519, B1 => n22271, B2 => 
                           n15480, ZN => n7093);
   U14710 : OAI22_X1 port map( A1 => n22281, A2 => n22385, B1 => n22280, B2 => 
                           n15469, ZN => n7102);
   U14711 : OAI22_X1 port map( A1 => n22281, A2 => n22387, B1 => n22280, B2 => 
                           n15468, ZN => n7103);
   U14712 : OAI22_X1 port map( A1 => n22281, A2 => n22393, B1 => n22280, B2 => 
                           n15467, ZN => n7104);
   U14713 : OAI22_X1 port map( A1 => n22281, A2 => n22399, B1 => n22280, B2 => 
                           n15466, ZN => n7105);
   U14714 : OAI22_X1 port map( A1 => n22281, A2 => n22405, B1 => n22280, B2 => 
                           n15465, ZN => n7106);
   U14715 : OAI22_X1 port map( A1 => n22282, A2 => n22411, B1 => n22280, B2 => 
                           n15464, ZN => n7107);
   U14716 : OAI22_X1 port map( A1 => n22282, A2 => n22417, B1 => n22280, B2 => 
                           n15463, ZN => n7108);
   U14717 : OAI22_X1 port map( A1 => n22282, A2 => n22423, B1 => n22280, B2 => 
                           n15462, ZN => n7109);
   U14718 : OAI22_X1 port map( A1 => n22282, A2 => n22429, B1 => n22280, B2 => 
                           n15461, ZN => n7110);
   U14719 : OAI22_X1 port map( A1 => n22282, A2 => n22435, B1 => n22280, B2 => 
                           n15460, ZN => n7111);
   U14720 : OAI22_X1 port map( A1 => n22283, A2 => n22441, B1 => n22280, B2 => 
                           n15459, ZN => n7112);
   U14721 : OAI22_X1 port map( A1 => n22283, A2 => n22447, B1 => n22280, B2 => 
                           n15458, ZN => n7113);
   U14722 : OAI22_X1 port map( A1 => n22283, A2 => n22453, B1 => n22280, B2 => 
                           n15457, ZN => n7114);
   U14723 : OAI22_X1 port map( A1 => n22283, A2 => n22459, B1 => n22280, B2 => 
                           n15456, ZN => n7115);
   U14724 : OAI22_X1 port map( A1 => n22283, A2 => n22465, B1 => n15437, B2 => 
                           n15455, ZN => n7116);
   U14725 : OAI22_X1 port map( A1 => n22284, A2 => n22471, B1 => n15437, B2 => 
                           n15454, ZN => n7117);
   U14726 : OAI22_X1 port map( A1 => n22284, A2 => n22477, B1 => n15437, B2 => 
                           n15453, ZN => n7118);
   U14727 : OAI22_X1 port map( A1 => n22284, A2 => n22483, B1 => n15437, B2 => 
                           n15452, ZN => n7119);
   U14728 : OAI22_X1 port map( A1 => n22284, A2 => n22489, B1 => n15437, B2 => 
                           n15451, ZN => n7120);
   U14729 : OAI22_X1 port map( A1 => n22284, A2 => n22495, B1 => n15437, B2 => 
                           n15450, ZN => n7121);
   U14730 : OAI22_X1 port map( A1 => n22285, A2 => n22501, B1 => n15437, B2 => 
                           n15449, ZN => n7122);
   U14731 : OAI22_X1 port map( A1 => n22285, A2 => n22507, B1 => n22280, B2 => 
                           n15448, ZN => n7123);
   U14732 : OAI22_X1 port map( A1 => n22285, A2 => n22513, B1 => n22280, B2 => 
                           n15447, ZN => n7124);
   U14733 : OAI22_X1 port map( A1 => n22285, A2 => n22519, B1 => n22280, B2 => 
                           n15446, ZN => n7125);
   U14734 : OAI22_X1 port map( A1 => n22290, A2 => n22385, B1 => n22289, B2 => 
                           n15435, ZN => n7134);
   U14735 : OAI22_X1 port map( A1 => n22290, A2 => n22387, B1 => n22289, B2 => 
                           n15434, ZN => n7135);
   U14736 : OAI22_X1 port map( A1 => n22290, A2 => n22393, B1 => n22289, B2 => 
                           n15433, ZN => n7136);
   U14737 : OAI22_X1 port map( A1 => n22290, A2 => n22399, B1 => n22289, B2 => 
                           n15432, ZN => n7137);
   U14738 : OAI22_X1 port map( A1 => n22290, A2 => n22405, B1 => n22289, B2 => 
                           n15431, ZN => n7138);
   U14739 : OAI22_X1 port map( A1 => n22291, A2 => n22411, B1 => n22289, B2 => 
                           n15430, ZN => n7139);
   U14740 : OAI22_X1 port map( A1 => n22291, A2 => n22417, B1 => n22289, B2 => 
                           n15429, ZN => n7140);
   U14741 : OAI22_X1 port map( A1 => n22291, A2 => n22423, B1 => n22289, B2 => 
                           n15428, ZN => n7141);
   U14742 : OAI22_X1 port map( A1 => n22291, A2 => n22429, B1 => n22289, B2 => 
                           n15427, ZN => n7142);
   U14743 : OAI22_X1 port map( A1 => n22291, A2 => n22435, B1 => n22289, B2 => 
                           n15426, ZN => n7143);
   U14744 : OAI22_X1 port map( A1 => n22292, A2 => n22441, B1 => n22289, B2 => 
                           n15425, ZN => n7144);
   U14745 : OAI22_X1 port map( A1 => n22292, A2 => n22447, B1 => n22289, B2 => 
                           n15424, ZN => n7145);
   U14746 : OAI22_X1 port map( A1 => n22292, A2 => n22453, B1 => n22289, B2 => 
                           n15423, ZN => n7146);
   U14747 : OAI22_X1 port map( A1 => n22292, A2 => n22459, B1 => n22289, B2 => 
                           n15422, ZN => n7147);
   U14748 : OAI22_X1 port map( A1 => n22292, A2 => n22465, B1 => n15403, B2 => 
                           n15421, ZN => n7148);
   U14749 : OAI22_X1 port map( A1 => n22293, A2 => n22471, B1 => n15403, B2 => 
                           n15420, ZN => n7149);
   U14750 : OAI22_X1 port map( A1 => n22293, A2 => n22477, B1 => n15403, B2 => 
                           n15419, ZN => n7150);
   U14751 : OAI22_X1 port map( A1 => n22293, A2 => n22483, B1 => n15403, B2 => 
                           n15418, ZN => n7151);
   U14752 : OAI22_X1 port map( A1 => n22293, A2 => n22489, B1 => n15403, B2 => 
                           n15417, ZN => n7152);
   U14753 : OAI22_X1 port map( A1 => n22293, A2 => n22495, B1 => n15403, B2 => 
                           n15416, ZN => n7153);
   U14754 : OAI22_X1 port map( A1 => n22294, A2 => n22501, B1 => n15403, B2 => 
                           n15415, ZN => n7154);
   U14755 : OAI22_X1 port map( A1 => n22294, A2 => n22507, B1 => n22289, B2 => 
                           n15414, ZN => n7155);
   U14756 : OAI22_X1 port map( A1 => n22294, A2 => n22513, B1 => n22289, B2 => 
                           n15413, ZN => n7156);
   U14757 : OAI22_X1 port map( A1 => n22294, A2 => n22519, B1 => n22289, B2 => 
                           n15412, ZN => n7157);
   U14758 : OAI22_X1 port map( A1 => n22299, A2 => n22385, B1 => n22298, B2 => 
                           n15400, ZN => n7166);
   U14759 : OAI22_X1 port map( A1 => n22299, A2 => n22387, B1 => n22298, B2 => 
                           n15399, ZN => n7167);
   U14760 : OAI22_X1 port map( A1 => n22299, A2 => n22393, B1 => n22298, B2 => 
                           n15398, ZN => n7168);
   U14761 : OAI22_X1 port map( A1 => n22299, A2 => n22399, B1 => n22298, B2 => 
                           n15397, ZN => n7169);
   U14762 : OAI22_X1 port map( A1 => n22299, A2 => n22405, B1 => n22298, B2 => 
                           n15396, ZN => n7170);
   U14763 : OAI22_X1 port map( A1 => n22300, A2 => n22411, B1 => n22298, B2 => 
                           n15395, ZN => n7171);
   U14764 : OAI22_X1 port map( A1 => n22300, A2 => n22417, B1 => n22298, B2 => 
                           n15394, ZN => n7172);
   U14765 : OAI22_X1 port map( A1 => n22300, A2 => n22423, B1 => n22298, B2 => 
                           n15393, ZN => n7173);
   U14766 : OAI22_X1 port map( A1 => n22300, A2 => n22429, B1 => n22298, B2 => 
                           n15392, ZN => n7174);
   U14767 : OAI22_X1 port map( A1 => n22300, A2 => n22435, B1 => n22298, B2 => 
                           n15391, ZN => n7175);
   U14768 : OAI22_X1 port map( A1 => n22301, A2 => n22441, B1 => n22298, B2 => 
                           n15390, ZN => n7176);
   U14769 : OAI22_X1 port map( A1 => n22301, A2 => n22447, B1 => n22298, B2 => 
                           n15389, ZN => n7177);
   U14770 : OAI22_X1 port map( A1 => n22301, A2 => n22453, B1 => n22298, B2 => 
                           n15388, ZN => n7178);
   U14771 : OAI22_X1 port map( A1 => n22301, A2 => n22459, B1 => n22298, B2 => 
                           n15387, ZN => n7179);
   U14772 : OAI22_X1 port map( A1 => n22301, A2 => n22465, B1 => n15368, B2 => 
                           n15386, ZN => n7180);
   U14773 : OAI22_X1 port map( A1 => n22302, A2 => n22471, B1 => n15368, B2 => 
                           n15385, ZN => n7181);
   U14774 : OAI22_X1 port map( A1 => n22302, A2 => n22477, B1 => n15368, B2 => 
                           n15384, ZN => n7182);
   U14775 : OAI22_X1 port map( A1 => n22302, A2 => n22483, B1 => n15368, B2 => 
                           n15383, ZN => n7183);
   U14776 : OAI22_X1 port map( A1 => n22302, A2 => n22489, B1 => n15368, B2 => 
                           n15382, ZN => n7184);
   U14777 : OAI22_X1 port map( A1 => n22302, A2 => n22495, B1 => n15368, B2 => 
                           n15381, ZN => n7185);
   U14778 : OAI22_X1 port map( A1 => n22303, A2 => n22501, B1 => n15368, B2 => 
                           n15380, ZN => n7186);
   U14779 : OAI22_X1 port map( A1 => n22303, A2 => n22507, B1 => n22298, B2 => 
                           n15379, ZN => n7187);
   U14780 : OAI22_X1 port map( A1 => n22303, A2 => n22513, B1 => n22298, B2 => 
                           n15378, ZN => n7188);
   U14781 : OAI22_X1 port map( A1 => n22303, A2 => n22519, B1 => n22298, B2 => 
                           n15377, ZN => n7189);
   U14782 : OAI22_X1 port map( A1 => n22326, A2 => n22385, B1 => n22325, B2 => 
                           n15297, ZN => n7262);
   U14783 : OAI22_X1 port map( A1 => n22326, A2 => n22387, B1 => n22325, B2 => 
                           n15296, ZN => n7263);
   U14784 : OAI22_X1 port map( A1 => n22326, A2 => n22393, B1 => n22325, B2 => 
                           n15295, ZN => n7264);
   U14785 : OAI22_X1 port map( A1 => n22326, A2 => n22399, B1 => n22325, B2 => 
                           n15294, ZN => n7265);
   U14786 : OAI22_X1 port map( A1 => n22326, A2 => n22405, B1 => n22325, B2 => 
                           n15293, ZN => n7266);
   U14787 : OAI22_X1 port map( A1 => n22327, A2 => n22411, B1 => n22325, B2 => 
                           n15292, ZN => n7267);
   U14788 : OAI22_X1 port map( A1 => n22327, A2 => n22417, B1 => n22325, B2 => 
                           n15291, ZN => n7268);
   U14789 : OAI22_X1 port map( A1 => n22327, A2 => n22423, B1 => n22325, B2 => 
                           n15290, ZN => n7269);
   U14790 : OAI22_X1 port map( A1 => n22327, A2 => n22429, B1 => n22325, B2 => 
                           n15289, ZN => n7270);
   U14791 : OAI22_X1 port map( A1 => n22327, A2 => n22435, B1 => n22325, B2 => 
                           n15288, ZN => n7271);
   U14792 : OAI22_X1 port map( A1 => n22328, A2 => n22441, B1 => n22325, B2 => 
                           n15287, ZN => n7272);
   U14793 : OAI22_X1 port map( A1 => n22328, A2 => n22447, B1 => n22325, B2 => 
                           n15286, ZN => n7273);
   U14794 : OAI22_X1 port map( A1 => n22328, A2 => n22453, B1 => n22325, B2 => 
                           n15285, ZN => n7274);
   U14795 : OAI22_X1 port map( A1 => n22328, A2 => n22459, B1 => n22325, B2 => 
                           n15284, ZN => n7275);
   U14796 : OAI22_X1 port map( A1 => n22328, A2 => n22465, B1 => n15265, B2 => 
                           n15283, ZN => n7276);
   U14797 : OAI22_X1 port map( A1 => n22329, A2 => n22471, B1 => n15265, B2 => 
                           n15282, ZN => n7277);
   U14798 : OAI22_X1 port map( A1 => n22329, A2 => n22477, B1 => n15265, B2 => 
                           n15281, ZN => n7278);
   U14799 : OAI22_X1 port map( A1 => n22329, A2 => n22483, B1 => n15265, B2 => 
                           n15280, ZN => n7279);
   U14800 : OAI22_X1 port map( A1 => n22329, A2 => n22489, B1 => n15265, B2 => 
                           n15279, ZN => n7280);
   U14801 : OAI22_X1 port map( A1 => n22329, A2 => n22495, B1 => n15265, B2 => 
                           n15278, ZN => n7281);
   U14802 : OAI22_X1 port map( A1 => n22330, A2 => n22501, B1 => n15265, B2 => 
                           n15277, ZN => n7282);
   U14803 : OAI22_X1 port map( A1 => n22330, A2 => n22507, B1 => n22325, B2 => 
                           n15276, ZN => n7283);
   U14804 : OAI22_X1 port map( A1 => n22330, A2 => n22513, B1 => n22325, B2 => 
                           n15275, ZN => n7284);
   U14805 : OAI22_X1 port map( A1 => n22330, A2 => n22519, B1 => n22325, B2 => 
                           n15274, ZN => n7285);
   U14806 : OAI22_X1 port map( A1 => n22335, A2 => n22385, B1 => n22334, B2 => 
                           n15262, ZN => n7294);
   U14807 : OAI22_X1 port map( A1 => n22335, A2 => n22387, B1 => n22334, B2 => 
                           n15261, ZN => n7295);
   U14808 : OAI22_X1 port map( A1 => n22335, A2 => n22393, B1 => n22334, B2 => 
                           n15260, ZN => n7296);
   U14809 : OAI22_X1 port map( A1 => n22335, A2 => n22399, B1 => n22334, B2 => 
                           n15259, ZN => n7297);
   U14810 : OAI22_X1 port map( A1 => n22335, A2 => n22405, B1 => n22334, B2 => 
                           n15258, ZN => n7298);
   U14811 : OAI22_X1 port map( A1 => n22336, A2 => n22411, B1 => n22334, B2 => 
                           n15257, ZN => n7299);
   U14812 : OAI22_X1 port map( A1 => n22336, A2 => n22417, B1 => n22334, B2 => 
                           n15256, ZN => n7300);
   U14813 : OAI22_X1 port map( A1 => n22336, A2 => n22423, B1 => n22334, B2 => 
                           n15255, ZN => n7301);
   U14814 : OAI22_X1 port map( A1 => n22336, A2 => n22429, B1 => n22334, B2 => 
                           n15254, ZN => n7302);
   U14815 : OAI22_X1 port map( A1 => n22336, A2 => n22435, B1 => n22334, B2 => 
                           n15253, ZN => n7303);
   U14816 : OAI22_X1 port map( A1 => n22337, A2 => n22441, B1 => n22334, B2 => 
                           n15252, ZN => n7304);
   U14817 : OAI22_X1 port map( A1 => n22337, A2 => n22447, B1 => n22334, B2 => 
                           n15251, ZN => n7305);
   U14818 : OAI22_X1 port map( A1 => n22337, A2 => n22453, B1 => n22334, B2 => 
                           n15250, ZN => n7306);
   U14819 : OAI22_X1 port map( A1 => n22337, A2 => n22459, B1 => n22334, B2 => 
                           n15249, ZN => n7307);
   U14820 : OAI22_X1 port map( A1 => n22337, A2 => n22465, B1 => n15230, B2 => 
                           n15248, ZN => n7308);
   U14821 : OAI22_X1 port map( A1 => n22338, A2 => n22471, B1 => n15230, B2 => 
                           n15247, ZN => n7309);
   U14822 : OAI22_X1 port map( A1 => n22338, A2 => n22477, B1 => n15230, B2 => 
                           n15246, ZN => n7310);
   U14823 : OAI22_X1 port map( A1 => n22338, A2 => n22483, B1 => n15230, B2 => 
                           n15245, ZN => n7311);
   U14824 : OAI22_X1 port map( A1 => n22338, A2 => n22489, B1 => n15230, B2 => 
                           n15244, ZN => n7312);
   U14825 : OAI22_X1 port map( A1 => n22338, A2 => n22495, B1 => n15230, B2 => 
                           n15243, ZN => n7313);
   U14826 : OAI22_X1 port map( A1 => n22339, A2 => n22501, B1 => n15230, B2 => 
                           n15242, ZN => n7314);
   U14827 : OAI22_X1 port map( A1 => n22339, A2 => n22507, B1 => n22334, B2 => 
                           n15241, ZN => n7315);
   U14828 : OAI22_X1 port map( A1 => n22339, A2 => n22513, B1 => n22334, B2 => 
                           n15240, ZN => n7316);
   U14829 : OAI22_X1 port map( A1 => n22339, A2 => n22519, B1 => n22334, B2 => 
                           n15239, ZN => n7317);
   U14830 : BUF_X1 port map( A => n18472, Z => n20796);
   U14831 : BUF_X1 port map( A => n16893, Z => n21353);
   U14832 : BUF_X1 port map( A => n18477, Z => n20863);
   U14833 : BUF_X1 port map( A => n16898, Z => n21420);
   U14834 : BUF_X1 port map( A => n18472, Z => n20795);
   U14835 : BUF_X1 port map( A => n16893, Z => n21352);
   U14836 : BUF_X1 port map( A => n18472, Z => n20792);
   U14837 : BUF_X1 port map( A => n18477, Z => n20859);
   U14838 : BUF_X1 port map( A => n18472, Z => n20794);
   U14839 : BUF_X1 port map( A => n18477, Z => n20861);
   U14840 : BUF_X1 port map( A => n18472, Z => n20793);
   U14841 : BUF_X1 port map( A => n18477, Z => n20860);
   U14842 : BUF_X1 port map( A => n18477, Z => n20862);
   U14843 : BUF_X1 port map( A => n16893, Z => n21349);
   U14844 : BUF_X1 port map( A => n16898, Z => n21416);
   U14845 : BUF_X1 port map( A => n16893, Z => n21351);
   U14846 : BUF_X1 port map( A => n16898, Z => n21418);
   U14847 : BUF_X1 port map( A => n16893, Z => n21350);
   U14848 : BUF_X1 port map( A => n16898, Z => n21417);
   U14849 : BUF_X1 port map( A => n16898, Z => n21419);
   U14850 : BUF_X1 port map( A => n18468, Z => n20992);
   U14851 : BUF_X1 port map( A => n16888, Z => n21549);
   U14852 : BUF_X1 port map( A => n18463, Z => n21037);
   U14853 : BUF_X1 port map( A => n16882, Z => n21594);
   U14854 : BUF_X1 port map( A => n18472, Z => n20797);
   U14855 : BUF_X1 port map( A => n18477, Z => n20864);
   U14856 : BUF_X1 port map( A => n16893, Z => n21354);
   U14857 : BUF_X1 port map( A => n16898, Z => n21421);
   U14858 : NAND2_X1 port map( A1 => n16611, A2 => n15642, ZN => n16793);
   U14859 : NAND2_X1 port map( A1 => n16611, A2 => n15504, ZN => n16688);
   U14860 : NAND2_X1 port map( A1 => n16611, A2 => n15366, ZN => n16614);
   U14861 : NAND2_X1 port map( A1 => n16611, A2 => n15228, ZN => n16554);
   U14862 : NAND2_X1 port map( A1 => n16204, A2 => n15642, ZN => n16417);
   U14863 : NAND2_X1 port map( A1 => n16204, A2 => n15504, ZN => n16344);
   U14864 : NAND2_X1 port map( A1 => n16204, A2 => n15366, ZN => n16239);
   U14865 : NAND2_X1 port map( A1 => n16204, A2 => n15228, ZN => n16133);
   U14866 : NAND2_X1 port map( A1 => n15751, A2 => n15642, ZN => n15996);
   U14867 : NAND2_X1 port map( A1 => n15751, A2 => n15504, ZN => n15891);
   U14868 : NAND2_X1 port map( A1 => n15751, A2 => n15366, ZN => n15786);
   U14869 : NAND2_X1 port map( A1 => n15751, A2 => n15228, ZN => n15680);
   U14870 : NAND2_X1 port map( A1 => n15642, A2 => n15227, ZN => n15539);
   U14871 : NAND2_X1 port map( A1 => n15504, A2 => n15227, ZN => n15401);
   U14872 : NAND2_X1 port map( A1 => n15366, A2 => n15227, ZN => n15263);
   U14873 : AND3_X1 port map( A1 => n15643, A2 => n15644, A3 => n15645, ZN => 
                           n15227);
   U14874 : NAND2_X1 port map( A1 => n15227, A2 => n15228, ZN => n15151);
   U14875 : AND2_X1 port map( A1 => n19625, A2 => n20932, ZN => n18450);
   U14876 : AND2_X1 port map( A1 => n19625, A2 => n19673, ZN => n18490);
   U14877 : AND2_X1 port map( A1 => n19625, A2 => n19674, ZN => n18491);
   U14878 : AND2_X1 port map( A1 => n19625, A2 => n19634, ZN => n18501);
   U14879 : AND2_X1 port map( A1 => n19625, A2 => n19637, ZN => n18431);
   U14880 : AND2_X1 port map( A1 => n19625, A2 => n19626, ZN => n18441);
   U14881 : AND2_X1 port map( A1 => n18352, A2 => n21489, ZN => n16868);
   U14882 : AND2_X1 port map( A1 => n18352, A2 => n18409, ZN => n16915);
   U14883 : AND2_X1 port map( A1 => n18352, A2 => n18410, ZN => n16916);
   U14884 : AND2_X1 port map( A1 => n18352, A2 => n18361, ZN => n16928);
   U14885 : AND2_X1 port map( A1 => n18352, A2 => n18365, ZN => n16848);
   U14886 : AND2_X1 port map( A1 => n18352, A2 => n18353, ZN => n16859);
   U14887 : AND2_X1 port map( A1 => n19670, A2 => n19661, ZN => n20945);
   U14888 : AND2_X1 port map( A1 => n19677, A2 => n19661, ZN => n20806);
   U14889 : AND2_X1 port map( A1 => n19662, A2 => n19661, ZN => n20993);
   U14890 : AND2_X1 port map( A1 => n18405, A2 => n18394, ZN => n21502);
   U14891 : AND2_X1 port map( A1 => n18414, A2 => n18394, ZN => n21363);
   U14892 : AND2_X1 port map( A1 => n18395, A2 => n18394, ZN => n21550);
   U14893 : AND2_X1 port map( A1 => n19662, A2 => n19661, ZN => n18470);
   U14894 : AND2_X1 port map( A1 => n19677, A2 => n19661, ZN => n18476);
   U14895 : AND2_X1 port map( A1 => n18395, A2 => n18394, ZN => n16890);
   U14896 : AND2_X1 port map( A1 => n18414, A2 => n18394, ZN => n16897);
   U14897 : AND2_X1 port map( A1 => n19670, A2 => n19661, ZN => n18480);
   U14898 : AND2_X1 port map( A1 => n18405, A2 => n18394, ZN => n16901);
   U14899 : AND2_X1 port map( A1 => n19660, A2 => n19661, ZN => n21071);
   U14900 : AND2_X1 port map( A1 => n18393, A2 => n18394, ZN => n21628);
   U14901 : AND2_X1 port map( A1 => n19660, A2 => n19661, ZN => n18466);
   U14902 : AND2_X1 port map( A1 => n18393, A2 => n18394, ZN => n16885);
   U14903 : AND2_X1 port map( A1 => n19625, A2 => n20974, ZN => n18451);
   U14904 : AND2_X1 port map( A1 => n19625, A2 => n21100, ZN => n18437);
   U14905 : AND2_X1 port map( A1 => n18352, A2 => n21531, ZN => n16869);
   U14906 : AND2_X1 port map( A1 => n18352, A2 => n21657, ZN => n16855);
   U14907 : OAI21_X1 port map( B1 => n15226, B2 => n16793, A => n22375, ZN => 
                           n16832);
   U14908 : INV_X1 port map( A => n16797, ZN => n21829);
   U14909 : OAI21_X1 port map( B1 => n15156, B2 => n16793, A => n22380, ZN => 
                           n16797);
   U14910 : INV_X1 port map( A => n16758, ZN => n21847);
   U14911 : OAI21_X1 port map( B1 => n15226, B2 => n16688, A => n22380, ZN => 
                           n16758);
   U14912 : INV_X1 port map( A => n16690, ZN => n21865);
   U14913 : OAI21_X1 port map( B1 => n15156, B2 => n16688, A => n22379, ZN => 
                           n16690);
   U14914 : INV_X1 port map( A => n16620, ZN => n21883);
   U14915 : OAI21_X1 port map( B1 => n15226, B2 => n16614, A => n22380, ZN => 
                           n16620);
   U14916 : INV_X1 port map( A => n16616, ZN => n21901);
   U14917 : OAI21_X1 port map( B1 => n15156, B2 => n16614, A => n22379, ZN => 
                           n16616);
   U14918 : INV_X1 port map( A => n16610, ZN => n21919);
   U14919 : OAI21_X1 port map( B1 => n15226, B2 => n16554, A => n22379, ZN => 
                           n16610);
   U14920 : INV_X1 port map( A => n16556, ZN => n21937);
   U14921 : OAI21_X1 port map( B1 => n15156, B2 => n16554, A => n22379, ZN => 
                           n16556);
   U14922 : INV_X1 port map( A => n16487, ZN => n21955);
   U14923 : OAI21_X1 port map( B1 => n15226, B2 => n16417, A => n22379, ZN => 
                           n16487);
   U14924 : INV_X1 port map( A => n16419, ZN => n21973);
   U14925 : OAI21_X1 port map( B1 => n15156, B2 => n16417, A => n22378, ZN => 
                           n16419);
   U14926 : INV_X1 port map( A => n16350, ZN => n21991);
   U14927 : OAI21_X1 port map( B1 => n15226, B2 => n16344, A => n22379, ZN => 
                           n16350);
   U14928 : INV_X1 port map( A => n16346, ZN => n22009);
   U14929 : OAI21_X1 port map( B1 => n15156, B2 => n16344, A => n22379, ZN => 
                           n16346);
   U14930 : INV_X1 port map( A => n16309, ZN => n22027);
   U14931 : OAI21_X1 port map( B1 => n15226, B2 => n16239, A => n22378, ZN => 
                           n16309);
   U14932 : INV_X1 port map( A => n16241, ZN => n22045);
   U14933 : OAI21_X1 port map( B1 => n15156, B2 => n16239, A => n22378, ZN => 
                           n16241);
   U14934 : INV_X1 port map( A => n16171, ZN => n22063);
   U14935 : OAI21_X1 port map( B1 => n15226, B2 => n16133, A => n22378, ZN => 
                           n16171);
   U14936 : INV_X1 port map( A => n16135, ZN => n22081);
   U14937 : OAI21_X1 port map( B1 => n15156, B2 => n16133, A => n22378, ZN => 
                           n16135);
   U14938 : INV_X1 port map( A => n16066, ZN => n22099);
   U14939 : OAI21_X1 port map( B1 => n15226, B2 => n15996, A => n22378, ZN => 
                           n16066);
   U14940 : INV_X1 port map( A => n15998, ZN => n22117);
   U14941 : OAI21_X1 port map( B1 => n15156, B2 => n15996, A => n22377, ZN => 
                           n15998);
   U14942 : INV_X1 port map( A => n15929, ZN => n22135);
   U14943 : OAI21_X1 port map( B1 => n15226, B2 => n15891, A => n22377, ZN => 
                           n15929);
   U14944 : INV_X1 port map( A => n15893, ZN => n22153);
   U14945 : OAI21_X1 port map( B1 => n15156, B2 => n15891, A => n22377, ZN => 
                           n15893);
   U14946 : INV_X1 port map( A => n15856, ZN => n22171);
   U14947 : OAI21_X1 port map( B1 => n15226, B2 => n15786, A => n22377, ZN => 
                           n15856);
   U14948 : INV_X1 port map( A => n15788, ZN => n22189);
   U14949 : OAI21_X1 port map( B1 => n15156, B2 => n15786, A => n22377, ZN => 
                           n15788);
   U14950 : INV_X1 port map( A => n15750, ZN => n22207);
   U14951 : OAI21_X1 port map( B1 => n15226, B2 => n15680, A => n22377, ZN => 
                           n15750);
   U14952 : INV_X1 port map( A => n15682, ZN => n22225);
   U14953 : OAI21_X1 port map( B1 => n15156, B2 => n15680, A => n22377, ZN => 
                           n15682);
   U14954 : INV_X1 port map( A => n15609, ZN => n22243);
   U14955 : OAI21_X1 port map( B1 => n15226, B2 => n15539, A => n22376, ZN => 
                           n15609);
   U14956 : INV_X1 port map( A => n15541, ZN => n22261);
   U14957 : OAI21_X1 port map( B1 => n15156, B2 => n15539, A => n22376, ZN => 
                           n15541);
   U14958 : INV_X1 port map( A => n15471, ZN => n22279);
   U14959 : OAI21_X1 port map( B1 => n15226, B2 => n15401, A => n22376, ZN => 
                           n15471);
   U14960 : INV_X1 port map( A => n15403, ZN => n22297);
   U14961 : OAI21_X1 port map( B1 => n15156, B2 => n15401, A => n22376, ZN => 
                           n15403);
   U14962 : INV_X1 port map( A => n15333, ZN => n22315);
   U14963 : OAI21_X1 port map( B1 => n15226, B2 => n15263, A => n22376, ZN => 
                           n15333);
   U14964 : INV_X1 port map( A => n15265, ZN => n22333);
   U14965 : OAI21_X1 port map( B1 => n15156, B2 => n15263, A => n22376, ZN => 
                           n15265);
   U14966 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => n19645, ZN => n21104);
   U14967 : NAND2_X1 port map( A1 => ADD_RD1(0), A2 => n19645, ZN => n18454);
   U14968 : NAND2_X1 port map( A1 => ADD_RD2(0), A2 => n18374, ZN => n21661);
   U14969 : NAND2_X1 port map( A1 => ADD_RD2(0), A2 => n18374, ZN => n16873);
   U14970 : NOR2_X2 port map( A1 => n19645, A2 => ADD_RD1(0), ZN => n19625);
   U14971 : NOR2_X2 port map( A1 => n18374, A2 => ADD_RD2(0), ZN => n18352);
   U14972 : NOR3_X1 port map( A1 => n19665, A2 => ADD_RD1(5), A3 => n19666, ZN 
                           => n19662);
   U14973 : NOR3_X1 port map( A1 => n18399, A2 => ADD_RD2(5), A3 => n18400, ZN 
                           => n18395);
   U14974 : NOR3_X1 port map( A1 => n19671, A2 => ADD_RD1(4), A3 => n19665, ZN 
                           => n19670);
   U14975 : NOR3_X1 port map( A1 => n18406, A2 => ADD_RD2(4), A3 => n18399, ZN 
                           => n18405);
   U14976 : AOI221_X1 port map( B1 => n18450, B2 => n8915, C1 => n20979, C2 => 
                           n19692, A => n19642, ZN => n19641);
   U14977 : OAI222_X1 port map( A1 => n19643, A2 => n21104, B1 => n19644, B2 =>
                           n21105, C1 => n16382, C2 => n21108, ZN => n19642);
   U14978 : NOR4_X1 port map( A1 => n19655, A2 => n19656, A3 => n19657, A4 => 
                           n19658, ZN => n19643);
   U14979 : NOR4_X1 port map( A1 => n19647, A2 => n19648, A3 => n19649, A4 => 
                           n19650, ZN => n19644);
   U14980 : AOI221_X1 port map( B1 => n20938, B2 => n8904, C1 => n20980, C2 => 
                           n19693, A => n19593, ZN => n19592);
   U14981 : OAI222_X1 port map( A1 => n19594, A2 => n18454, B1 => n19595, B2 =>
                           n21106, C1 => n16381, C2 => n21109, ZN => n19593);
   U14982 : NOR4_X1 port map( A1 => n19604, A2 => n19605, A3 => n19606, A4 => 
                           n19607, ZN => n19594);
   U14983 : NOR4_X1 port map( A1 => n19596, A2 => n19597, A3 => n19598, A4 => 
                           n19599, ZN => n19595);
   U14984 : AOI221_X1 port map( B1 => n20938, B2 => n8893, C1 => n20978, C2 => 
                           n19694, A => n19556, ZN => n19555);
   U14985 : OAI222_X1 port map( A1 => n19557, A2 => n21104, B1 => n19558, B2 =>
                           n18456, C1 => n16380, C2 => n21107, ZN => n19556);
   U14986 : NOR4_X1 port map( A1 => n19567, A2 => n19568, A3 => n19569, A4 => 
                           n19570, ZN => n19557);
   U14987 : NOR4_X1 port map( A1 => n19559, A2 => n19560, A3 => n19561, A4 => 
                           n19562, ZN => n19558);
   U14988 : AOI221_X1 port map( B1 => n20939, B2 => n8882, C1 => n20978, C2 => 
                           n19695, A => n19519, ZN => n19518);
   U14989 : OAI222_X1 port map( A1 => n19520, A2 => n18454, B1 => n19521, B2 =>
                           n21105, C1 => n16379, C2 => n21107, ZN => n19519);
   U14990 : NOR4_X1 port map( A1 => n19530, A2 => n19531, A3 => n19532, A4 => 
                           n19533, ZN => n19520);
   U14991 : NOR4_X1 port map( A1 => n19522, A2 => n19523, A3 => n19524, A4 => 
                           n19525, ZN => n19521);
   U14992 : AOI221_X1 port map( B1 => n20940, B2 => n8871, C1 => n20979, C2 => 
                           n19696, A => n19482, ZN => n19481);
   U14993 : OAI222_X1 port map( A1 => n19483, A2 => n21104, B1 => n19484, B2 =>
                           n21106, C1 => n16378, C2 => n21108, ZN => n19482);
   U14994 : NOR4_X1 port map( A1 => n19493, A2 => n19494, A3 => n19495, A4 => 
                           n19496, ZN => n19483);
   U14995 : NOR4_X1 port map( A1 => n19485, A2 => n19486, A3 => n19487, A4 => 
                           n19488, ZN => n19484);
   U14996 : AOI221_X1 port map( B1 => n20940, B2 => n8860, C1 => n20979, C2 => 
                           n19697, A => n19445, ZN => n19444);
   U14997 : OAI222_X1 port map( A1 => n19446, A2 => n18454, B1 => n19447, B2 =>
                           n18456, C1 => n16377, C2 => n21108, ZN => n19445);
   U14998 : NOR4_X1 port map( A1 => n19456, A2 => n19457, A3 => n19458, A4 => 
                           n19459, ZN => n19446);
   U14999 : NOR4_X1 port map( A1 => n19448, A2 => n19449, A3 => n19450, A4 => 
                           n19451, ZN => n19447);
   U15000 : AOI221_X1 port map( B1 => n20943, B2 => n8849, C1 => n20980, C2 => 
                           n19698, A => n19408, ZN => n19407);
   U15001 : OAI222_X1 port map( A1 => n19409, A2 => n21104, B1 => n19410, B2 =>
                           n21105, C1 => n16376, C2 => n21109, ZN => n19408);
   U15002 : NOR4_X1 port map( A1 => n19419, A2 => n19420, A3 => n19421, A4 => 
                           n19422, ZN => n19409);
   U15003 : NOR4_X1 port map( A1 => n19411, A2 => n19412, A3 => n19413, A4 => 
                           n19414, ZN => n19410);
   U15004 : AOI221_X1 port map( B1 => n20940, B2 => n8838, C1 => n20978, C2 => 
                           n19699, A => n19371, ZN => n19370);
   U15005 : OAI222_X1 port map( A1 => n19372, A2 => n18454, B1 => n19373, B2 =>
                           n21106, C1 => n16375, C2 => n21107, ZN => n19371);
   U15006 : NOR4_X1 port map( A1 => n19382, A2 => n19383, A3 => n19384, A4 => 
                           n19385, ZN => n19372);
   U15007 : NOR4_X1 port map( A1 => n19374, A2 => n19375, A3 => n19376, A4 => 
                           n19377, ZN => n19373);
   U15008 : AOI221_X1 port map( B1 => n20944, B2 => n8827, C1 => n20980, C2 => 
                           n19700, A => n19334, ZN => n19333);
   U15009 : OAI222_X1 port map( A1 => n19335, A2 => n21104, B1 => n19336, B2 =>
                           n18456, C1 => n16374, C2 => n21109, ZN => n19334);
   U15010 : NOR4_X1 port map( A1 => n19345, A2 => n19346, A3 => n19347, A4 => 
                           n19348, ZN => n19335);
   U15011 : NOR4_X1 port map( A1 => n19337, A2 => n19338, A3 => n19339, A4 => 
                           n19340, ZN => n19336);
   U15012 : AOI221_X1 port map( B1 => n20941, B2 => n8816, C1 => n20979, C2 => 
                           n19701, A => n19297, ZN => n19296);
   U15013 : OAI222_X1 port map( A1 => n19298, A2 => n18454, B1 => n19299, B2 =>
                           n21105, C1 => n16373, C2 => n21108, ZN => n19297);
   U15014 : NOR4_X1 port map( A1 => n19308, A2 => n19309, A3 => n19310, A4 => 
                           n19311, ZN => n19298);
   U15015 : NOR4_X1 port map( A1 => n19300, A2 => n19301, A3 => n19302, A4 => 
                           n19303, ZN => n19299);
   U15016 : AOI221_X1 port map( B1 => n20941, B2 => n8805, C1 => n20980, C2 => 
                           n19702, A => n19260, ZN => n19259);
   U15017 : OAI222_X1 port map( A1 => n19261, A2 => n21104, B1 => n19262, B2 =>
                           n21106, C1 => n16372, C2 => n21109, ZN => n19260);
   U15018 : NOR4_X1 port map( A1 => n19271, A2 => n19272, A3 => n19273, A4 => 
                           n19274, ZN => n19261);
   U15019 : NOR4_X1 port map( A1 => n19263, A2 => n19264, A3 => n19265, A4 => 
                           n19266, ZN => n19262);
   U15020 : AOI221_X1 port map( B1 => n20942, B2 => n8794, C1 => n20978, C2 => 
                           n19703, A => n19223, ZN => n19222);
   U15021 : OAI222_X1 port map( A1 => n19224, A2 => n18454, B1 => n19225, B2 =>
                           n18456, C1 => n16371, C2 => n21107, ZN => n19223);
   U15022 : NOR4_X1 port map( A1 => n19234, A2 => n19235, A3 => n19236, A4 => 
                           n19237, ZN => n19224);
   U15023 : NOR4_X1 port map( A1 => n19226, A2 => n19227, A3 => n19228, A4 => 
                           n19229, ZN => n19225);
   U15024 : AOI221_X1 port map( B1 => n20943, B2 => n8783, C1 => n20978, C2 => 
                           n19704, A => n19186, ZN => n19185);
   U15025 : OAI222_X1 port map( A1 => n19187, A2 => n21104, B1 => n19188, B2 =>
                           n21105, C1 => n16370, C2 => n21107, ZN => n19186);
   U15026 : NOR4_X1 port map( A1 => n19197, A2 => n19198, A3 => n19199, A4 => 
                           n19200, ZN => n19187);
   U15027 : NOR4_X1 port map( A1 => n19189, A2 => n19190, A3 => n19191, A4 => 
                           n19192, ZN => n19188);
   U15028 : AOI221_X1 port map( B1 => n20943, B2 => n8772, C1 => n20979, C2 => 
                           n19705, A => n19149, ZN => n19148);
   U15029 : OAI222_X1 port map( A1 => n19150, A2 => n18454, B1 => n19151, B2 =>
                           n21106, C1 => n16369, C2 => n21108, ZN => n19149);
   U15030 : NOR4_X1 port map( A1 => n19160, A2 => n19161, A3 => n19162, A4 => 
                           n19163, ZN => n19150);
   U15031 : NOR4_X1 port map( A1 => n19152, A2 => n19153, A3 => n19154, A4 => 
                           n19155, ZN => n19151);
   U15032 : AOI221_X1 port map( B1 => n20941, B2 => n8761, C1 => n20979, C2 => 
                           n19706, A => n19112, ZN => n19111);
   U15033 : OAI222_X1 port map( A1 => n19113, A2 => n21104, B1 => n19114, B2 =>
                           n18456, C1 => n16368, C2 => n21108, ZN => n19112);
   U15034 : NOR4_X1 port map( A1 => n19123, A2 => n19124, A3 => n19125, A4 => 
                           n19126, ZN => n19113);
   U15035 : NOR4_X1 port map( A1 => n19115, A2 => n19116, A3 => n19117, A4 => 
                           n19118, ZN => n19114);
   U15036 : AOI221_X1 port map( B1 => n20942, B2 => n8750, C1 => n20980, C2 => 
                           n19707, A => n19075, ZN => n19074);
   U15037 : OAI222_X1 port map( A1 => n19076, A2 => n18454, B1 => n19077, B2 =>
                           n21105, C1 => n16367, C2 => n21109, ZN => n19075);
   U15038 : NOR4_X1 port map( A1 => n19086, A2 => n19087, A3 => n19088, A4 => 
                           n19089, ZN => n19076);
   U15039 : NOR4_X1 port map( A1 => n19078, A2 => n19079, A3 => n19080, A4 => 
                           n19081, ZN => n19077);
   U15040 : AOI221_X1 port map( B1 => n20943, B2 => n8739, C1 => n20978, C2 => 
                           n19708, A => n19038, ZN => n19037);
   U15041 : OAI222_X1 port map( A1 => n19039, A2 => n21104, B1 => n19040, B2 =>
                           n21106, C1 => n16366, C2 => n21107, ZN => n19038);
   U15042 : NOR4_X1 port map( A1 => n19049, A2 => n19050, A3 => n19051, A4 => 
                           n19052, ZN => n19039);
   U15043 : NOR4_X1 port map( A1 => n19041, A2 => n19042, A3 => n19043, A4 => 
                           n19044, ZN => n19040);
   U15044 : AOI221_X1 port map( B1 => n20943, B2 => n8728, C1 => n20980, C2 => 
                           n19709, A => n19001, ZN => n19000);
   U15045 : OAI222_X1 port map( A1 => n19002, A2 => n18454, B1 => n19003, B2 =>
                           n18456, C1 => n16365, C2 => n21109, ZN => n19001);
   U15046 : NOR4_X1 port map( A1 => n19012, A2 => n19013, A3 => n19014, A4 => 
                           n19015, ZN => n19002);
   U15047 : NOR4_X1 port map( A1 => n19004, A2 => n19005, A3 => n19006, A4 => 
                           n19007, ZN => n19003);
   U15048 : AOI221_X1 port map( B1 => n20944, B2 => n8717, C1 => n20979, C2 => 
                           n19710, A => n18964, ZN => n18963);
   U15049 : OAI222_X1 port map( A1 => n18965, A2 => n21104, B1 => n18966, B2 =>
                           n21105, C1 => n16364, C2 => n21108, ZN => n18964);
   U15050 : NOR4_X1 port map( A1 => n18975, A2 => n18976, A3 => n18977, A4 => 
                           n18978, ZN => n18965);
   U15051 : AOI221_X1 port map( B1 => n20944, B2 => n8706, C1 => n20980, C2 => 
                           n19711, A => n18927, ZN => n18926);
   U15052 : OAI222_X1 port map( A1 => n18928, A2 => n18454, B1 => n18929, B2 =>
                           n21106, C1 => n16363, C2 => n21109, ZN => n18927);
   U15053 : NOR4_X1 port map( A1 => n18938, A2 => n18939, A3 => n18940, A4 => 
                           n18941, ZN => n18928);
   U15054 : AOI221_X1 port map( B1 => n20944, B2 => n8695, C1 => n20978, C2 => 
                           n19712, A => n18890, ZN => n18889);
   U15055 : OAI222_X1 port map( A1 => n18891, A2 => n21104, B1 => n18892, B2 =>
                           n18456, C1 => n16362, C2 => n21107, ZN => n18890);
   U15056 : NOR4_X1 port map( A1 => n18901, A2 => n18902, A3 => n18903, A4 => 
                           n18904, ZN => n18891);
   U15057 : AOI221_X1 port map( B1 => n20944, B2 => n8684, C1 => n20978, C2 => 
                           n19681, A => n18853, ZN => n18852);
   U15058 : OAI222_X1 port map( A1 => n18854, A2 => n18454, B1 => n18855, B2 =>
                           n21105, C1 => n16361, C2 => n21107, ZN => n18853);
   U15059 : NOR4_X1 port map( A1 => n18864, A2 => n18865, A3 => n18866, A4 => 
                           n18867, ZN => n18854);
   U15060 : AOI221_X1 port map( B1 => n20938, B2 => n8673, C1 => n20979, C2 => 
                           n19713, A => n18816, ZN => n18815);
   U15061 : OAI222_X1 port map( A1 => n18817, A2 => n21104, B1 => n18818, B2 =>
                           n21106, C1 => n16360, C2 => n21108, ZN => n18816);
   U15062 : NOR4_X1 port map( A1 => n18827, A2 => n18828, A3 => n18829, A4 => 
                           n18830, ZN => n18817);
   U15063 : NOR4_X1 port map( A1 => n18819, A2 => n18820, A3 => n18821, A4 => 
                           n18822, ZN => n18818);
   U15064 : AOI221_X1 port map( B1 => n20938, B2 => n8662, C1 => n20979, C2 => 
                           n19714, A => n18779, ZN => n18778);
   U15065 : OAI222_X1 port map( A1 => n18780, A2 => n18454, B1 => n18781, B2 =>
                           n18456, C1 => n16359, C2 => n21108, ZN => n18779);
   U15066 : NOR4_X1 port map( A1 => n18790, A2 => n18791, A3 => n18792, A4 => 
                           n18793, ZN => n18780);
   U15067 : NOR4_X1 port map( A1 => n18782, A2 => n18783, A3 => n18784, A4 => 
                           n18785, ZN => n18781);
   U15068 : AOI221_X1 port map( B1 => n20938, B2 => n8651, C1 => n20980, C2 => 
                           n19715, A => n18742, ZN => n18741);
   U15069 : OAI222_X1 port map( A1 => n18743, A2 => n21104, B1 => n18744, B2 =>
                           n21105, C1 => n16358, C2 => n21109, ZN => n18742);
   U15070 : NOR4_X1 port map( A1 => n18753, A2 => n18754, A3 => n18755, A4 => 
                           n18756, ZN => n18743);
   U15071 : NOR4_X1 port map( A1 => n18745, A2 => n18746, A3 => n18747, A4 => 
                           n18748, ZN => n18744);
   U15072 : AOI221_X1 port map( B1 => n20939, B2 => n8640, C1 => n20978, C2 => 
                           n19716, A => n18705, ZN => n18704);
   U15073 : OAI222_X1 port map( A1 => n18706, A2 => n18454, B1 => n18707, B2 =>
                           n21106, C1 => n16357, C2 => n21107, ZN => n18705);
   U15074 : NOR4_X1 port map( A1 => n18716, A2 => n18717, A3 => n18718, A4 => 
                           n18719, ZN => n18706);
   U15075 : NOR4_X1 port map( A1 => n18708, A2 => n18709, A3 => n18710, A4 => 
                           n18711, ZN => n18707);
   U15076 : AOI221_X1 port map( B1 => n20940, B2 => n8629, C1 => n20980, C2 => 
                           n19717, A => n18668, ZN => n18667);
   U15077 : OAI222_X1 port map( A1 => n18669, A2 => n21104, B1 => n18670, B2 =>
                           n18456, C1 => n16356, C2 => n21109, ZN => n18668);
   U15078 : NOR4_X1 port map( A1 => n18679, A2 => n18680, A3 => n18681, A4 => 
                           n18682, ZN => n18669);
   U15079 : NOR4_X1 port map( A1 => n18671, A2 => n18672, A3 => n18673, A4 => 
                           n18674, ZN => n18670);
   U15080 : AOI221_X1 port map( B1 => n20939, B2 => n8618, C1 => n20979, C2 => 
                           n19718, A => n18631, ZN => n18630);
   U15081 : OAI222_X1 port map( A1 => n18632, A2 => n18454, B1 => n18633, B2 =>
                           n21105, C1 => n16355, C2 => n21108, ZN => n18631);
   U15082 : NOR4_X1 port map( A1 => n18642, A2 => n18643, A3 => n18644, A4 => 
                           n18645, ZN => n18632);
   U15083 : NOR4_X1 port map( A1 => n18634, A2 => n18635, A3 => n18636, A4 => 
                           n18637, ZN => n18633);
   U15084 : AOI221_X1 port map( B1 => n20943, B2 => n8607, C1 => n20980, C2 => 
                           n19719, A => n18594, ZN => n18593);
   U15085 : OAI222_X1 port map( A1 => n18595, A2 => n21104, B1 => n18596, B2 =>
                           n21106, C1 => n16354, C2 => n21109, ZN => n18594);
   U15086 : NOR4_X1 port map( A1 => n18605, A2 => n18606, A3 => n18607, A4 => 
                           n18608, ZN => n18595);
   U15087 : NOR4_X1 port map( A1 => n18597, A2 => n18598, A3 => n18599, A4 => 
                           n18600, ZN => n18596);
   U15088 : AOI221_X1 port map( B1 => n20940, B2 => n8596, C1 => n20978, C2 => 
                           n19720, A => n18557, ZN => n18556);
   U15089 : OAI222_X1 port map( A1 => n18558, A2 => n18454, B1 => n18559, B2 =>
                           n18456, C1 => n16353, C2 => n21107, ZN => n18557);
   U15090 : NOR4_X1 port map( A1 => n18568, A2 => n18569, A3 => n18570, A4 => 
                           n18571, ZN => n18558);
   U15091 : NOR4_X1 port map( A1 => n18560, A2 => n18561, A3 => n18562, A4 => 
                           n18563, ZN => n18559);
   U15092 : AOI221_X1 port map( B1 => n20939, B2 => n8585, C1 => n20978, C2 => 
                           n19721, A => n18520, ZN => n18519);
   U15093 : OAI222_X1 port map( A1 => n18521, A2 => n21104, B1 => n18522, B2 =>
                           n21105, C1 => n16352, C2 => n21107, ZN => n18520);
   U15094 : NOR4_X1 port map( A1 => n18531, A2 => n18532, A3 => n18533, A4 => 
                           n18534, ZN => n18521);
   U15095 : NOR4_X1 port map( A1 => n18523, A2 => n18524, A3 => n18525, A4 => 
                           n18526, ZN => n18522);
   U15096 : AOI221_X1 port map( B1 => n20942, B2 => n8574, C1 => n20979, C2 => 
                           n19722, A => n18452, ZN => n18449);
   U15097 : OAI222_X1 port map( A1 => n18453, A2 => n18454, B1 => n18455, B2 =>
                           n21106, C1 => n16351, C2 => n21108, ZN => n18452);
   U15098 : NOR4_X1 port map( A1 => n18482, A2 => n18483, A3 => n18484, A4 => 
                           n18485, ZN => n18453);
   U15099 : NOR4_X1 port map( A1 => n18458, A2 => n18459, A3 => n18460, A4 => 
                           n18461, ZN => n18455);
   U15100 : AOI221_X1 port map( B1 => n16868, B2 => n8915, C1 => n21536, C2 => 
                           n19692, A => n18371, ZN => n18369);
   U15101 : OAI222_X1 port map( A1 => n18372, A2 => n21661, B1 => n18373, B2 =>
                           n21662, C1 => n16382, C2 => n21665, ZN => n18371);
   U15102 : NOR4_X1 port map( A1 => n18387, A2 => n18388, A3 => n18389, A4 => 
                           n18390, ZN => n18372);
   U15103 : NOR4_X1 port map( A1 => n18376, A2 => n18377, A3 => n18378, A4 => 
                           n18379, ZN => n18373);
   U15104 : AOI221_X1 port map( B1 => n21495, B2 => n8904, C1 => n21537, C2 => 
                           n19693, A => n18312, ZN => n18310);
   U15105 : OAI222_X1 port map( A1 => n18313, A2 => n16873, B1 => n18314, B2 =>
                           n21663, C1 => n16381, C2 => n21666, ZN => n18312);
   U15106 : NOR4_X1 port map( A1 => n18326, A2 => n18327, A3 => n18328, A4 => 
                           n18329, ZN => n18313);
   U15107 : NOR4_X1 port map( A1 => n18315, A2 => n18316, A3 => n18317, A4 => 
                           n18318, ZN => n18314);
   U15108 : AOI221_X1 port map( B1 => n21495, B2 => n8893, C1 => n21535, C2 => 
                           n19694, A => n18265, ZN => n18263);
   U15109 : OAI222_X1 port map( A1 => n18266, A2 => n21661, B1 => n18267, B2 =>
                           n16875, C1 => n16380, C2 => n21664, ZN => n18265);
   U15110 : NOR4_X1 port map( A1 => n18279, A2 => n18280, A3 => n18281, A4 => 
                           n18282, ZN => n18266);
   U15111 : NOR4_X1 port map( A1 => n18268, A2 => n18269, A3 => n18270, A4 => 
                           n18271, ZN => n18267);
   U15112 : AOI221_X1 port map( B1 => n21496, B2 => n8882, C1 => n21535, C2 => 
                           n19695, A => n18218, ZN => n18216);
   U15113 : OAI222_X1 port map( A1 => n18219, A2 => n16873, B1 => n18220, B2 =>
                           n21662, C1 => n16379, C2 => n21664, ZN => n18218);
   U15114 : NOR4_X1 port map( A1 => n18232, A2 => n18233, A3 => n18234, A4 => 
                           n18235, ZN => n18219);
   U15115 : NOR4_X1 port map( A1 => n18221, A2 => n18222, A3 => n18223, A4 => 
                           n18224, ZN => n18220);
   U15116 : AOI221_X1 port map( B1 => n21497, B2 => n8871, C1 => n21536, C2 => 
                           n19696, A => n18171, ZN => n18169);
   U15117 : OAI222_X1 port map( A1 => n18172, A2 => n21661, B1 => n18173, B2 =>
                           n21663, C1 => n16378, C2 => n21665, ZN => n18171);
   U15118 : NOR4_X1 port map( A1 => n18185, A2 => n18186, A3 => n18187, A4 => 
                           n18188, ZN => n18172);
   U15119 : NOR4_X1 port map( A1 => n18174, A2 => n18175, A3 => n18176, A4 => 
                           n18177, ZN => n18173);
   U15120 : AOI221_X1 port map( B1 => n21497, B2 => n8860, C1 => n21536, C2 => 
                           n19697, A => n18124, ZN => n18122);
   U15121 : OAI222_X1 port map( A1 => n18125, A2 => n16873, B1 => n18126, B2 =>
                           n16875, C1 => n16377, C2 => n21665, ZN => n18124);
   U15122 : NOR4_X1 port map( A1 => n18138, A2 => n18139, A3 => n18140, A4 => 
                           n18141, ZN => n18125);
   U15123 : NOR4_X1 port map( A1 => n18127, A2 => n18128, A3 => n18129, A4 => 
                           n18130, ZN => n18126);
   U15124 : AOI221_X1 port map( B1 => n21500, B2 => n8849, C1 => n21537, C2 => 
                           n19698, A => n18077, ZN => n18075);
   U15125 : OAI222_X1 port map( A1 => n18078, A2 => n21661, B1 => n18079, B2 =>
                           n21662, C1 => n16376, C2 => n21666, ZN => n18077);
   U15126 : NOR4_X1 port map( A1 => n18091, A2 => n18092, A3 => n18093, A4 => 
                           n18094, ZN => n18078);
   U15127 : NOR4_X1 port map( A1 => n18080, A2 => n18081, A3 => n18082, A4 => 
                           n18083, ZN => n18079);
   U15128 : AOI221_X1 port map( B1 => n21497, B2 => n8838, C1 => n21535, C2 => 
                           n19699, A => n18030, ZN => n18028);
   U15129 : OAI222_X1 port map( A1 => n18031, A2 => n16873, B1 => n18032, B2 =>
                           n21663, C1 => n16375, C2 => n21664, ZN => n18030);
   U15130 : NOR4_X1 port map( A1 => n18044, A2 => n18045, A3 => n18046, A4 => 
                           n18047, ZN => n18031);
   U15131 : NOR4_X1 port map( A1 => n18033, A2 => n18034, A3 => n18035, A4 => 
                           n18036, ZN => n18032);
   U15132 : AOI221_X1 port map( B1 => n21501, B2 => n8827, C1 => n21537, C2 => 
                           n19700, A => n17983, ZN => n17981);
   U15133 : OAI222_X1 port map( A1 => n17984, A2 => n21661, B1 => n17985, B2 =>
                           n16875, C1 => n16374, C2 => n21666, ZN => n17983);
   U15134 : NOR4_X1 port map( A1 => n17997, A2 => n17998, A3 => n17999, A4 => 
                           n18000, ZN => n17984);
   U15135 : NOR4_X1 port map( A1 => n17986, A2 => n17987, A3 => n17988, A4 => 
                           n17989, ZN => n17985);
   U15136 : AOI221_X1 port map( B1 => n21498, B2 => n8816, C1 => n21536, C2 => 
                           n19701, A => n17936, ZN => n17934);
   U15137 : OAI222_X1 port map( A1 => n17937, A2 => n16873, B1 => n17938, B2 =>
                           n21662, C1 => n16373, C2 => n21665, ZN => n17936);
   U15138 : NOR4_X1 port map( A1 => n17950, A2 => n17951, A3 => n17952, A4 => 
                           n17953, ZN => n17937);
   U15139 : NOR4_X1 port map( A1 => n17939, A2 => n17940, A3 => n17941, A4 => 
                           n17942, ZN => n17938);
   U15140 : AOI221_X1 port map( B1 => n21498, B2 => n8805, C1 => n21537, C2 => 
                           n19702, A => n17889, ZN => n17887);
   U15141 : OAI222_X1 port map( A1 => n17890, A2 => n21661, B1 => n17891, B2 =>
                           n21663, C1 => n16372, C2 => n21666, ZN => n17889);
   U15142 : NOR4_X1 port map( A1 => n17903, A2 => n17904, A3 => n17905, A4 => 
                           n17906, ZN => n17890);
   U15143 : NOR4_X1 port map( A1 => n17892, A2 => n17893, A3 => n17894, A4 => 
                           n17895, ZN => n17891);
   U15144 : AOI221_X1 port map( B1 => n21499, B2 => n8794, C1 => n21535, C2 => 
                           n19703, A => n17842, ZN => n17840);
   U15145 : OAI222_X1 port map( A1 => n17843, A2 => n16873, B1 => n17844, B2 =>
                           n16875, C1 => n16371, C2 => n21664, ZN => n17842);
   U15146 : NOR4_X1 port map( A1 => n17856, A2 => n17857, A3 => n17858, A4 => 
                           n17859, ZN => n17843);
   U15147 : NOR4_X1 port map( A1 => n17845, A2 => n17846, A3 => n17847, A4 => 
                           n17848, ZN => n17844);
   U15148 : AOI221_X1 port map( B1 => n21500, B2 => n8783, C1 => n21535, C2 => 
                           n19704, A => n17795, ZN => n17793);
   U15149 : OAI222_X1 port map( A1 => n17796, A2 => n21661, B1 => n17797, B2 =>
                           n21662, C1 => n16370, C2 => n21664, ZN => n17795);
   U15150 : NOR4_X1 port map( A1 => n17809, A2 => n17810, A3 => n17811, A4 => 
                           n17812, ZN => n17796);
   U15151 : NOR4_X1 port map( A1 => n17798, A2 => n17799, A3 => n17800, A4 => 
                           n17801, ZN => n17797);
   U15152 : AOI221_X1 port map( B1 => n21500, B2 => n8772, C1 => n21536, C2 => 
                           n19705, A => n17748, ZN => n17746);
   U15153 : OAI222_X1 port map( A1 => n17749, A2 => n16873, B1 => n17750, B2 =>
                           n21663, C1 => n16369, C2 => n21665, ZN => n17748);
   U15154 : NOR4_X1 port map( A1 => n17762, A2 => n17763, A3 => n17764, A4 => 
                           n17765, ZN => n17749);
   U15155 : NOR4_X1 port map( A1 => n17751, A2 => n17752, A3 => n17753, A4 => 
                           n17754, ZN => n17750);
   U15156 : AOI221_X1 port map( B1 => n21498, B2 => n8761, C1 => n21536, C2 => 
                           n19706, A => n17701, ZN => n17699);
   U15157 : OAI222_X1 port map( A1 => n17702, A2 => n21661, B1 => n17703, B2 =>
                           n16875, C1 => n16368, C2 => n21665, ZN => n17701);
   U15158 : NOR4_X1 port map( A1 => n17715, A2 => n17716, A3 => n17717, A4 => 
                           n17718, ZN => n17702);
   U15159 : NOR4_X1 port map( A1 => n17704, A2 => n17705, A3 => n17706, A4 => 
                           n17707, ZN => n17703);
   U15160 : AOI221_X1 port map( B1 => n21499, B2 => n8750, C1 => n21537, C2 => 
                           n19707, A => n17654, ZN => n17652);
   U15161 : OAI222_X1 port map( A1 => n17655, A2 => n16873, B1 => n17656, B2 =>
                           n21662, C1 => n16367, C2 => n21666, ZN => n17654);
   U15162 : NOR4_X1 port map( A1 => n17668, A2 => n17669, A3 => n17670, A4 => 
                           n17671, ZN => n17655);
   U15163 : NOR4_X1 port map( A1 => n17657, A2 => n17658, A3 => n17659, A4 => 
                           n17660, ZN => n17656);
   U15164 : AOI221_X1 port map( B1 => n21500, B2 => n8739, C1 => n21535, C2 => 
                           n19708, A => n17607, ZN => n17605);
   U15165 : OAI222_X1 port map( A1 => n17608, A2 => n21661, B1 => n17609, B2 =>
                           n21663, C1 => n16366, C2 => n21664, ZN => n17607);
   U15166 : NOR4_X1 port map( A1 => n17621, A2 => n17622, A3 => n17623, A4 => 
                           n17624, ZN => n17608);
   U15167 : NOR4_X1 port map( A1 => n17610, A2 => n17611, A3 => n17612, A4 => 
                           n17613, ZN => n17609);
   U15168 : AOI221_X1 port map( B1 => n21500, B2 => n8728, C1 => n21537, C2 => 
                           n19709, A => n17560, ZN => n17558);
   U15169 : OAI222_X1 port map( A1 => n17561, A2 => n16873, B1 => n17562, B2 =>
                           n16875, C1 => n16365, C2 => n21666, ZN => n17560);
   U15170 : NOR4_X1 port map( A1 => n17574, A2 => n17575, A3 => n17576, A4 => 
                           n17577, ZN => n17561);
   U15171 : NOR4_X1 port map( A1 => n17563, A2 => n17564, A3 => n17565, A4 => 
                           n17566, ZN => n17562);
   U15172 : AOI221_X1 port map( B1 => n21501, B2 => n8717, C1 => n21536, C2 => 
                           n19710, A => n17513, ZN => n17511);
   U15173 : OAI222_X1 port map( A1 => n17514, A2 => n21661, B1 => n17515, B2 =>
                           n21662, C1 => n16364, C2 => n21665, ZN => n17513);
   U15174 : NOR4_X1 port map( A1 => n17527, A2 => n17528, A3 => n17529, A4 => 
                           n17530, ZN => n17514);
   U15175 : AOI221_X1 port map( B1 => n21501, B2 => n8706, C1 => n21537, C2 => 
                           n19711, A => n17466, ZN => n17464);
   U15176 : OAI222_X1 port map( A1 => n17467, A2 => n16873, B1 => n17468, B2 =>
                           n21663, C1 => n16363, C2 => n21666, ZN => n17466);
   U15177 : NOR4_X1 port map( A1 => n17480, A2 => n17481, A3 => n17482, A4 => 
                           n17483, ZN => n17467);
   U15178 : AOI221_X1 port map( B1 => n21501, B2 => n8695, C1 => n21535, C2 => 
                           n19712, A => n17419, ZN => n17417);
   U15179 : OAI222_X1 port map( A1 => n17420, A2 => n21661, B1 => n17421, B2 =>
                           n16875, C1 => n16362, C2 => n21664, ZN => n17419);
   U15180 : NOR4_X1 port map( A1 => n17433, A2 => n17434, A3 => n17435, A4 => 
                           n17436, ZN => n17420);
   U15181 : AOI221_X1 port map( B1 => n21501, B2 => n8684, C1 => n21535, C2 => 
                           n19681, A => n17372, ZN => n17370);
   U15182 : OAI222_X1 port map( A1 => n17373, A2 => n16873, B1 => n17374, B2 =>
                           n21662, C1 => n16361, C2 => n21664, ZN => n17372);
   U15183 : NOR4_X1 port map( A1 => n17386, A2 => n17387, A3 => n17388, A4 => 
                           n17389, ZN => n17373);
   U15184 : AOI221_X1 port map( B1 => n21495, B2 => n8673, C1 => n21536, C2 => 
                           n19713, A => n17325, ZN => n17323);
   U15185 : OAI222_X1 port map( A1 => n17326, A2 => n21661, B1 => n17327, B2 =>
                           n21663, C1 => n16360, C2 => n21665, ZN => n17325);
   U15186 : NOR4_X1 port map( A1 => n17339, A2 => n17340, A3 => n17341, A4 => 
                           n17342, ZN => n17326);
   U15187 : NOR4_X1 port map( A1 => n17328, A2 => n17329, A3 => n17330, A4 => 
                           n17331, ZN => n17327);
   U15188 : AOI221_X1 port map( B1 => n21495, B2 => n8662, C1 => n21536, C2 => 
                           n19714, A => n17278, ZN => n17276);
   U15189 : OAI222_X1 port map( A1 => n17279, A2 => n16873, B1 => n17280, B2 =>
                           n16875, C1 => n16359, C2 => n21665, ZN => n17278);
   U15190 : NOR4_X1 port map( A1 => n17292, A2 => n17293, A3 => n17294, A4 => 
                           n17295, ZN => n17279);
   U15191 : NOR4_X1 port map( A1 => n17281, A2 => n17282, A3 => n17283, A4 => 
                           n17284, ZN => n17280);
   U15192 : AOI221_X1 port map( B1 => n21495, B2 => n8651, C1 => n21537, C2 => 
                           n19715, A => n17231, ZN => n17229);
   U15193 : OAI222_X1 port map( A1 => n17232, A2 => n21661, B1 => n17233, B2 =>
                           n21662, C1 => n16358, C2 => n21666, ZN => n17231);
   U15194 : NOR4_X1 port map( A1 => n17245, A2 => n17246, A3 => n17247, A4 => 
                           n17248, ZN => n17232);
   U15195 : NOR4_X1 port map( A1 => n17234, A2 => n17235, A3 => n17236, A4 => 
                           n17237, ZN => n17233);
   U15196 : AOI221_X1 port map( B1 => n21496, B2 => n8640, C1 => n21535, C2 => 
                           n19716, A => n17184, ZN => n17182);
   U15197 : OAI222_X1 port map( A1 => n17185, A2 => n16873, B1 => n17186, B2 =>
                           n21663, C1 => n16357, C2 => n21664, ZN => n17184);
   U15198 : NOR4_X1 port map( A1 => n17198, A2 => n17199, A3 => n17200, A4 => 
                           n17201, ZN => n17185);
   U15199 : NOR4_X1 port map( A1 => n17187, A2 => n17188, A3 => n17189, A4 => 
                           n17190, ZN => n17186);
   U15200 : AOI221_X1 port map( B1 => n21497, B2 => n8629, C1 => n21537, C2 => 
                           n19717, A => n17137, ZN => n17135);
   U15201 : OAI222_X1 port map( A1 => n17138, A2 => n21661, B1 => n17139, B2 =>
                           n16875, C1 => n16356, C2 => n21666, ZN => n17137);
   U15202 : NOR4_X1 port map( A1 => n17151, A2 => n17152, A3 => n17153, A4 => 
                           n17154, ZN => n17138);
   U15203 : NOR4_X1 port map( A1 => n17140, A2 => n17141, A3 => n17142, A4 => 
                           n17143, ZN => n17139);
   U15204 : AOI221_X1 port map( B1 => n21496, B2 => n8618, C1 => n21536, C2 => 
                           n19718, A => n17090, ZN => n17088);
   U15205 : OAI222_X1 port map( A1 => n17091, A2 => n16873, B1 => n17092, B2 =>
                           n21662, C1 => n16355, C2 => n21665, ZN => n17090);
   U15206 : NOR4_X1 port map( A1 => n17104, A2 => n17105, A3 => n17106, A4 => 
                           n17107, ZN => n17091);
   U15207 : NOR4_X1 port map( A1 => n17093, A2 => n17094, A3 => n17095, A4 => 
                           n17096, ZN => n17092);
   U15208 : AOI221_X1 port map( B1 => n21500, B2 => n8607, C1 => n21537, C2 => 
                           n19719, A => n17043, ZN => n17041);
   U15209 : OAI222_X1 port map( A1 => n17044, A2 => n21661, B1 => n17045, B2 =>
                           n21663, C1 => n16354, C2 => n21666, ZN => n17043);
   U15210 : NOR4_X1 port map( A1 => n17057, A2 => n17058, A3 => n17059, A4 => 
                           n17060, ZN => n17044);
   U15211 : NOR4_X1 port map( A1 => n17046, A2 => n17047, A3 => n17048, A4 => 
                           n17049, ZN => n17045);
   U15212 : AOI221_X1 port map( B1 => n21497, B2 => n8596, C1 => n21535, C2 => 
                           n19720, A => n16996, ZN => n16994);
   U15213 : OAI222_X1 port map( A1 => n16997, A2 => n16873, B1 => n16998, B2 =>
                           n16875, C1 => n16353, C2 => n21664, ZN => n16996);
   U15214 : NOR4_X1 port map( A1 => n17010, A2 => n17011, A3 => n17012, A4 => 
                           n17013, ZN => n16997);
   U15215 : NOR4_X1 port map( A1 => n16999, A2 => n17000, A3 => n17001, A4 => 
                           n17002, ZN => n16998);
   U15216 : AOI221_X1 port map( B1 => n21496, B2 => n8585, C1 => n21535, C2 => 
                           n19721, A => n16949, ZN => n16947);
   U15217 : OAI222_X1 port map( A1 => n16950, A2 => n21661, B1 => n16951, B2 =>
                           n21662, C1 => n16352, C2 => n21664, ZN => n16949);
   U15218 : NOR4_X1 port map( A1 => n16963, A2 => n16964, A3 => n16965, A4 => 
                           n16966, ZN => n16950);
   U15219 : NOR4_X1 port map( A1 => n16952, A2 => n16953, A3 => n16954, A4 => 
                           n16955, ZN => n16951);
   U15220 : AOI221_X1 port map( B1 => n21499, B2 => n8574, C1 => n21536, C2 => 
                           n19722, A => n16871, ZN => n16867);
   U15221 : OAI222_X1 port map( A1 => n16872, A2 => n16873, B1 => n16874, B2 =>
                           n21663, C1 => n16351, C2 => n21665, ZN => n16871);
   U15222 : NOR4_X1 port map( A1 => n16904, A2 => n16905, A3 => n16906, A4 => 
                           n16907, ZN => n16872);
   U15223 : NOR4_X1 port map( A1 => n16877, A2 => n16878, A3 => n16879, A4 => 
                           n16880, ZN => n16874);
   U15224 : AOI221_X1 port map( B1 => n21144, B2 => n9532, C1 => n21155, C2 => 
                           n9628, A => n19585, ZN => n19584);
   U15225 : OAI222_X1 port map( A1 => n4479, A2 => n21182, B1 => n4511, B2 => 
                           n21170, C1 => n15926, C2 => n21161, ZN => n19585);
   U15226 : AOI221_X1 port map( B1 => n21149, B2 => n9531, C1 => n21153, C2 => 
                           n9627, A => n19548, ZN => n19547);
   U15227 : OAI222_X1 port map( A1 => n4480, A2 => n21178, B1 => n4512, B2 => 
                           n21169, C1 => n15925, C2 => n21166, ZN => n19548);
   U15228 : AOI221_X1 port map( B1 => n21150, B2 => n9530, C1 => n21153, C2 => 
                           n9626, A => n19511, ZN => n19510);
   U15229 : OAI222_X1 port map( A1 => n4481, A2 => n21178, B1 => n4513, B2 => 
                           n21170, C1 => n15924, C2 => n21162, ZN => n19511);
   U15230 : AOI221_X1 port map( B1 => n21145, B2 => n9529, C1 => n21154, C2 => 
                           n9625, A => n19474, ZN => n19473);
   U15231 : OAI222_X1 port map( A1 => n4482, A2 => n21179, B1 => n4514, B2 => 
                           n21171, C1 => n15923, C2 => n21164, ZN => n19474);
   U15232 : AOI221_X1 port map( B1 => n21144, B2 => n9528, C1 => n21154, C2 => 
                           n9624, A => n19437, ZN => n19436);
   U15233 : OAI222_X1 port map( A1 => n4483, A2 => n21180, B1 => n4515, B2 => 
                           n21171, C1 => n15922, C2 => n21163, ZN => n19437);
   U15234 : AOI221_X1 port map( B1 => n21148, B2 => n9527, C1 => n21154, C2 => 
                           n9623, A => n19400, ZN => n19399);
   U15235 : OAI222_X1 port map( A1 => n4484, A2 => n21180, B1 => n4516, B2 => 
                           n21175, C1 => n15921, C2 => n21164, ZN => n19400);
   U15236 : AOI221_X1 port map( B1 => n21146, B2 => n9526, C1 => n21155, C2 => 
                           n9622, A => n19363, ZN => n19362);
   U15237 : OAI222_X1 port map( A1 => n4485, A2 => n21183, B1 => n4517, B2 => 
                           n21171, C1 => n15920, C2 => n21164, ZN => n19363);
   U15238 : AOI221_X1 port map( B1 => n21147, B2 => n9525, C1 => n21155, C2 => 
                           n9621, A => n19326, ZN => n19325);
   U15239 : OAI222_X1 port map( A1 => n4486, A2 => n21179, B1 => n4518, B2 => 
                           n21172, C1 => n15919, C2 => n21162, ZN => n19326);
   U15240 : AOI221_X1 port map( B1 => n21146, B2 => n9524, C1 => n21156, C2 => 
                           n9620, A => n19289, ZN => n19288);
   U15241 : OAI222_X1 port map( A1 => n4487, A2 => n21181, B1 => n4519, B2 => 
                           n21173, C1 => n15918, C2 => n21165, ZN => n19289);
   U15242 : AOI221_X1 port map( B1 => n21147, B2 => n9523, C1 => n21157, C2 => 
                           n9619, A => n19252, ZN => n19251);
   U15243 : OAI222_X1 port map( A1 => n4488, A2 => n21182, B1 => n4520, B2 => 
                           n21174, C1 => n15917, C2 => n21166, ZN => n19252);
   U15244 : AOI221_X1 port map( B1 => n21148, B2 => n9522, C1 => n21157, C2 => 
                           n9618, A => n19215, ZN => n19214);
   U15245 : OAI222_X1 port map( A1 => n4489, A2 => n21182, B1 => n4521, B2 => 
                           n21173, C1 => n15916, C2 => n21167, ZN => n19215);
   U15246 : AOI221_X1 port map( B1 => n21148, B2 => n9521, C1 => n21157, C2 => 
                           n9617, A => n19178, ZN => n19177);
   U15247 : OAI222_X1 port map( A1 => n4490, A2 => n21177, B1 => n4522, B2 => 
                           n21170, C1 => n15915, C2 => n21162, ZN => n19178);
   U15248 : AOI221_X1 port map( B1 => n21149, B2 => n9520, C1 => n21156, C2 => 
                           n9616, A => n19141, ZN => n19140);
   U15249 : OAI222_X1 port map( A1 => n4491, A2 => n21178, B1 => n4523, B2 => 
                           n21170, C1 => n15914, C2 => n21162, ZN => n19141);
   U15250 : AOI221_X1 port map( B1 => n21148, B2 => n9519, C1 => n21157, C2 => 
                           n9615, A => n19104, ZN => n19103);
   U15251 : OAI222_X1 port map( A1 => n4492, A2 => n21179, B1 => n4524, B2 => 
                           n21171, C1 => n15913, C2 => n21163, ZN => n19104);
   U15252 : AOI221_X1 port map( B1 => n21147, B2 => n9518, C1 => n21157, C2 => 
                           n9614, A => n19067, ZN => n19066);
   U15253 : OAI222_X1 port map( A1 => n4493, A2 => n21180, B1 => n4525, B2 => 
                           n21172, C1 => n15912, C2 => n21163, ZN => n19067);
   U15254 : AOI221_X1 port map( B1 => n21149, B2 => n9517, C1 => n21154, C2 => 
                           n9613, A => n19030, ZN => n19029);
   U15255 : OAI222_X1 port map( A1 => n4494, A2 => n21179, B1 => n4526, B2 => 
                           n21173, C1 => n15911, C2 => n21164, ZN => n19030);
   U15256 : AOI221_X1 port map( B1 => n21149, B2 => n9516, C1 => n21153, C2 => 
                           n9612, A => n18993, ZN => n18992);
   U15257 : OAI222_X1 port map( A1 => n4495, A2 => n21181, B1 => n4527, B2 => 
                           n21172, C1 => n15910, C2 => n21163, ZN => n18993);
   U15258 : AOI221_X1 port map( B1 => n21146, B2 => n9515, C1 => n21156, C2 => 
                           n9611, A => n18956, ZN => n18955);
   U15259 : OAI222_X1 port map( A1 => n4496, A2 => n21180, B1 => n4528, B2 => 
                           n21172, C1 => n15909, C2 => n21161, ZN => n18956);
   U15260 : AOI221_X1 port map( B1 => n21149, B2 => n9514, C1 => n21155, C2 => 
                           n9610, A => n18919, ZN => n18918);
   U15261 : OAI222_X1 port map( A1 => n4497, A2 => n21181, B1 => n4529, B2 => 
                           n21170, C1 => n15908, C2 => n21165, ZN => n18919);
   U15262 : AOI221_X1 port map( B1 => n21150, B2 => n9513, C1 => n21158, C2 => 
                           n9609, A => n18882, ZN => n18881);
   U15263 : OAI222_X1 port map( A1 => n4498, A2 => n21181, B1 => n4530, B2 => 
                           n21171, C1 => n15907, C2 => n21166, ZN => n18882);
   U15264 : AOI221_X1 port map( B1 => n21150, B2 => n9512, C1 => n21158, C2 => 
                           n9608, A => n18845, ZN => n18844);
   U15265 : OAI222_X1 port map( A1 => n4499, A2 => n21182, B1 => n4531, B2 => 
                           n21174, C1 => n15906, C2 => n21165, ZN => n18845);
   U15266 : AOI221_X1 port map( B1 => n21150, B2 => n9511, C1 => n21158, C2 => 
                           n9607, A => n18808, ZN => n18807);
   U15267 : OAI222_X1 port map( A1 => n4500, A2 => n21183, B1 => n4532, B2 => 
                           n21173, C1 => n15905, C2 => n21166, ZN => n18808);
   U15268 : AOI221_X1 port map( B1 => n21150, B2 => n9510, C1 => n21158, C2 => 
                           n9606, A => n18771, ZN => n18770);
   U15269 : OAI222_X1 port map( A1 => n4501, A2 => n21183, B1 => n4533, B2 => 
                           n21175, C1 => n15904, C2 => n21166, ZN => n18771);
   U15270 : AOI221_X1 port map( B1 => n21144, B2 => n9509, C1 => n21153, C2 => 
                           n9605, A => n18734, ZN => n18733);
   U15271 : OAI222_X1 port map( A1 => n4502, A2 => n21183, B1 => n4534, B2 => 
                           n21174, C1 => n15903, C2 => n21167, ZN => n18734);
   U15272 : AOI221_X1 port map( B1 => n21149, B2 => n9508, C1 => n21153, C2 => 
                           n9604, A => n18697, ZN => n18696);
   U15273 : OAI222_X1 port map( A1 => n4503, A2 => n21182, B1 => n4535, B2 => 
                           n21175, C1 => n15902, C2 => n21167, ZN => n18697);
   U15274 : AOI221_X1 port map( B1 => n21144, B2 => n9507, C1 => n21158, C2 => 
                           n9603, A => n18660, ZN => n18659);
   U15275 : OAI222_X1 port map( A1 => n4504, A2 => n21183, B1 => n4536, B2 => 
                           n21174, C1 => n15901, C2 => n21165, ZN => n18660);
   U15276 : AOI221_X1 port map( B1 => n21145, B2 => n9506, C1 => n21154, C2 => 
                           n9602, A => n18623, ZN => n18622);
   U15277 : OAI222_X1 port map( A1 => n4505, A2 => n21178, B1 => n4537, B2 => 
                           n21175, C1 => n15900, C2 => n21165, ZN => n18623);
   U15278 : AOI221_X1 port map( B1 => n21145, B2 => n9505, C1 => n21154, C2 => 
                           n9601, A => n18586, ZN => n18585);
   U15279 : OAI222_X1 port map( A1 => n4506, A2 => n21178, B1 => n4538, B2 => 
                           n21173, C1 => n15899, C2 => n21161, ZN => n18586);
   U15280 : AOI221_X1 port map( B1 => n21145, B2 => n9504, C1 => n21156, C2 => 
                           n9600, A => n18549, ZN => n18548);
   U15281 : OAI222_X1 port map( A1 => n4507, A2 => n21177, B1 => n4539, B2 => 
                           n21169, C1 => n15898, C2 => n21161, ZN => n18549);
   U15282 : AOI221_X1 port map( B1 => n21146, B2 => n9503, C1 => n21155, C2 => 
                           n9599, A => n18512, ZN => n18511);
   U15283 : OAI222_X1 port map( A1 => n4508, A2 => n21180, B1 => n4540, B2 => 
                           n21169, C1 => n15897, C2 => n21165, ZN => n18512);
   U15284 : AOI221_X1 port map( B1 => n21146, B2 => n9502, C1 => n21156, C2 => 
                           n9598, A => n18427, ZN => n18424);
   U15285 : OAI222_X1 port map( A1 => n4509, A2 => n21177, B1 => n4541, B2 => 
                           n21169, C1 => n15896, C2 => n21167, ZN => n18427);
   U15286 : AOI221_X1 port map( B1 => n21701, B2 => n9532, C1 => n21712, C2 => 
                           n9628, A => n18302, ZN => n18301);
   U15287 : OAI222_X1 port map( A1 => n4479, A2 => n21739, B1 => n4511, B2 => 
                           n21727, C1 => n15926, C2 => n21718, ZN => n18302);
   U15288 : AOI221_X1 port map( B1 => n21706, B2 => n9531, C1 => n21710, C2 => 
                           n9627, A => n18255, ZN => n18254);
   U15289 : OAI222_X1 port map( A1 => n4480, A2 => n21735, B1 => n4512, B2 => 
                           n21726, C1 => n15925, C2 => n21723, ZN => n18255);
   U15290 : AOI221_X1 port map( B1 => n21707, B2 => n9530, C1 => n21710, C2 => 
                           n9626, A => n18208, ZN => n18207);
   U15291 : OAI222_X1 port map( A1 => n4481, A2 => n21735, B1 => n4513, B2 => 
                           n21727, C1 => n15924, C2 => n21719, ZN => n18208);
   U15292 : AOI221_X1 port map( B1 => n21702, B2 => n9529, C1 => n21711, C2 => 
                           n9625, A => n18161, ZN => n18160);
   U15293 : OAI222_X1 port map( A1 => n4482, A2 => n21736, B1 => n4514, B2 => 
                           n21728, C1 => n15923, C2 => n21721, ZN => n18161);
   U15294 : AOI221_X1 port map( B1 => n21701, B2 => n9528, C1 => n21711, C2 => 
                           n9624, A => n18114, ZN => n18113);
   U15295 : OAI222_X1 port map( A1 => n4483, A2 => n21737, B1 => n4515, B2 => 
                           n21728, C1 => n15922, C2 => n21720, ZN => n18114);
   U15296 : AOI221_X1 port map( B1 => n21705, B2 => n9527, C1 => n21711, C2 => 
                           n9623, A => n18067, ZN => n18066);
   U15297 : OAI222_X1 port map( A1 => n4484, A2 => n21737, B1 => n4516, B2 => 
                           n21732, C1 => n15921, C2 => n21721, ZN => n18067);
   U15298 : AOI221_X1 port map( B1 => n21703, B2 => n9526, C1 => n21712, C2 => 
                           n9622, A => n18020, ZN => n18019);
   U15299 : OAI222_X1 port map( A1 => n4485, A2 => n21740, B1 => n4517, B2 => 
                           n21728, C1 => n15920, C2 => n21721, ZN => n18020);
   U15300 : AOI221_X1 port map( B1 => n21704, B2 => n9525, C1 => n21712, C2 => 
                           n9621, A => n17973, ZN => n17972);
   U15301 : OAI222_X1 port map( A1 => n4486, A2 => n21736, B1 => n4518, B2 => 
                           n21729, C1 => n15919, C2 => n21719, ZN => n17973);
   U15302 : AOI221_X1 port map( B1 => n21703, B2 => n9524, C1 => n21713, C2 => 
                           n9620, A => n17926, ZN => n17925);
   U15303 : OAI222_X1 port map( A1 => n4487, A2 => n21738, B1 => n4519, B2 => 
                           n21730, C1 => n15918, C2 => n21722, ZN => n17926);
   U15304 : AOI221_X1 port map( B1 => n21704, B2 => n9523, C1 => n21714, C2 => 
                           n9619, A => n17879, ZN => n17878);
   U15305 : OAI222_X1 port map( A1 => n4488, A2 => n21739, B1 => n4520, B2 => 
                           n21731, C1 => n15917, C2 => n21723, ZN => n17879);
   U15306 : AOI221_X1 port map( B1 => n21705, B2 => n9522, C1 => n21714, C2 => 
                           n9618, A => n17832, ZN => n17831);
   U15307 : OAI222_X1 port map( A1 => n4489, A2 => n21739, B1 => n4521, B2 => 
                           n21730, C1 => n15916, C2 => n21724, ZN => n17832);
   U15308 : AOI221_X1 port map( B1 => n21705, B2 => n9521, C1 => n21714, C2 => 
                           n9617, A => n17785, ZN => n17784);
   U15309 : OAI222_X1 port map( A1 => n4490, A2 => n21734, B1 => n4522, B2 => 
                           n21727, C1 => n15915, C2 => n21719, ZN => n17785);
   U15310 : AOI221_X1 port map( B1 => n21706, B2 => n9520, C1 => n21713, C2 => 
                           n9616, A => n17738, ZN => n17737);
   U15311 : OAI222_X1 port map( A1 => n4491, A2 => n21735, B1 => n4523, B2 => 
                           n21727, C1 => n15914, C2 => n21719, ZN => n17738);
   U15312 : AOI221_X1 port map( B1 => n21705, B2 => n9519, C1 => n21714, C2 => 
                           n9615, A => n17691, ZN => n17690);
   U15313 : OAI222_X1 port map( A1 => n4492, A2 => n21736, B1 => n4524, B2 => 
                           n21728, C1 => n15913, C2 => n21720, ZN => n17691);
   U15314 : AOI221_X1 port map( B1 => n21704, B2 => n9518, C1 => n21714, C2 => 
                           n9614, A => n17644, ZN => n17643);
   U15315 : OAI222_X1 port map( A1 => n4493, A2 => n21737, B1 => n4525, B2 => 
                           n21729, C1 => n15912, C2 => n21720, ZN => n17644);
   U15316 : AOI221_X1 port map( B1 => n21706, B2 => n9517, C1 => n21711, C2 => 
                           n9613, A => n17597, ZN => n17596);
   U15317 : OAI222_X1 port map( A1 => n4494, A2 => n21736, B1 => n4526, B2 => 
                           n21730, C1 => n15911, C2 => n21721, ZN => n17597);
   U15318 : AOI221_X1 port map( B1 => n21706, B2 => n9516, C1 => n21710, C2 => 
                           n9612, A => n17550, ZN => n17549);
   U15319 : OAI222_X1 port map( A1 => n4495, A2 => n21738, B1 => n4527, B2 => 
                           n21729, C1 => n15910, C2 => n21720, ZN => n17550);
   U15320 : AOI221_X1 port map( B1 => n21703, B2 => n9515, C1 => n21713, C2 => 
                           n9611, A => n17503, ZN => n17502);
   U15321 : OAI222_X1 port map( A1 => n4496, A2 => n21737, B1 => n4528, B2 => 
                           n21729, C1 => n15909, C2 => n21718, ZN => n17503);
   U15322 : AOI221_X1 port map( B1 => n21706, B2 => n9514, C1 => n21712, C2 => 
                           n9610, A => n17456, ZN => n17455);
   U15323 : OAI222_X1 port map( A1 => n4497, A2 => n21738, B1 => n4529, B2 => 
                           n21727, C1 => n15908, C2 => n21722, ZN => n17456);
   U15324 : AOI221_X1 port map( B1 => n21707, B2 => n9513, C1 => n21715, C2 => 
                           n9609, A => n17409, ZN => n17408);
   U15325 : OAI222_X1 port map( A1 => n4498, A2 => n21738, B1 => n4530, B2 => 
                           n21728, C1 => n15907, C2 => n21723, ZN => n17409);
   U15326 : AOI221_X1 port map( B1 => n21707, B2 => n9512, C1 => n21715, C2 => 
                           n9608, A => n17362, ZN => n17361);
   U15327 : OAI222_X1 port map( A1 => n4499, A2 => n21739, B1 => n4531, B2 => 
                           n21731, C1 => n15906, C2 => n21722, ZN => n17362);
   U15328 : AOI221_X1 port map( B1 => n21707, B2 => n9511, C1 => n21715, C2 => 
                           n9607, A => n17315, ZN => n17314);
   U15329 : OAI222_X1 port map( A1 => n4500, A2 => n21740, B1 => n4532, B2 => 
                           n21730, C1 => n15905, C2 => n21723, ZN => n17315);
   U15330 : AOI221_X1 port map( B1 => n21707, B2 => n9510, C1 => n21715, C2 => 
                           n9606, A => n17268, ZN => n17267);
   U15331 : OAI222_X1 port map( A1 => n4501, A2 => n21740, B1 => n4533, B2 => 
                           n21732, C1 => n15904, C2 => n21723, ZN => n17268);
   U15332 : AOI221_X1 port map( B1 => n21701, B2 => n9509, C1 => n21710, C2 => 
                           n9605, A => n17221, ZN => n17220);
   U15333 : OAI222_X1 port map( A1 => n4502, A2 => n21740, B1 => n4534, B2 => 
                           n21731, C1 => n15903, C2 => n21724, ZN => n17221);
   U15334 : AOI221_X1 port map( B1 => n21706, B2 => n9508, C1 => n21710, C2 => 
                           n9604, A => n17174, ZN => n17173);
   U15335 : OAI222_X1 port map( A1 => n4503, A2 => n21739, B1 => n4535, B2 => 
                           n21732, C1 => n15902, C2 => n21724, ZN => n17174);
   U15336 : AOI221_X1 port map( B1 => n21701, B2 => n9507, C1 => n21715, C2 => 
                           n9603, A => n17127, ZN => n17126);
   U15337 : OAI222_X1 port map( A1 => n4504, A2 => n21740, B1 => n4536, B2 => 
                           n21731, C1 => n15901, C2 => n21722, ZN => n17127);
   U15338 : AOI221_X1 port map( B1 => n21702, B2 => n9506, C1 => n21711, C2 => 
                           n9602, A => n17080, ZN => n17079);
   U15339 : OAI222_X1 port map( A1 => n4505, A2 => n21735, B1 => n4537, B2 => 
                           n21732, C1 => n15900, C2 => n21722, ZN => n17080);
   U15340 : AOI221_X1 port map( B1 => n21702, B2 => n9505, C1 => n21711, C2 => 
                           n9601, A => n17033, ZN => n17032);
   U15341 : OAI222_X1 port map( A1 => n4506, A2 => n21735, B1 => n4538, B2 => 
                           n21730, C1 => n15899, C2 => n21718, ZN => n17033);
   U15342 : AOI221_X1 port map( B1 => n21702, B2 => n9504, C1 => n21713, C2 => 
                           n9600, A => n16986, ZN => n16985);
   U15343 : OAI222_X1 port map( A1 => n4507, A2 => n21734, B1 => n4539, B2 => 
                           n21726, C1 => n15898, C2 => n21718, ZN => n16986);
   U15344 : AOI221_X1 port map( B1 => n21703, B2 => n9503, C1 => n21712, C2 => 
                           n9599, A => n16939, ZN => n16938);
   U15345 : OAI222_X1 port map( A1 => n4508, A2 => n21737, B1 => n4540, B2 => 
                           n21726, C1 => n15897, C2 => n21722, ZN => n16939);
   U15346 : AOI221_X1 port map( B1 => n21703, B2 => n9502, C1 => n21713, C2 => 
                           n9598, A => n16844, ZN => n16841);
   U15347 : OAI222_X1 port map( A1 => n4509, A2 => n21734, B1 => n4541, B2 => 
                           n21726, C1 => n15896, C2 => n21724, ZN => n16844);
   U15348 : NOR4_X1 port map( A1 => n18967, A2 => n18968, A3 => n18969, A4 => 
                           n18970, ZN => n18966);
   U15349 : OAI221_X1 port map( B1 => n16220, B2 => n20863, C1 => n16114, C2 =>
                           n20873, A => n18974, ZN => n18967);
   U15350 : OAI221_X1 port map( B1 => n8033, B2 => n20796, C1 => n16535, C2 => 
                           n20729, A => n18973, ZN => n18968);
   U15351 : OAI221_X1 port map( B1 => n15382, B2 => n21030, C1 => n15244, C2 =>
                           n21032, A => n18971, ZN => n18970);
   U15352 : NOR4_X1 port map( A1 => n18930, A2 => n18931, A3 => n18932, A4 => 
                           n18933, ZN => n18929);
   U15353 : OAI221_X1 port map( B1 => n16219, B2 => n20859, C1 => n16113, C2 =>
                           n20875, A => n18937, ZN => n18930);
   U15354 : OAI221_X1 port map( B1 => n8065, B2 => n20792, C1 => n16534, C2 => 
                           n20731, A => n18936, ZN => n18931);
   U15355 : OAI221_X1 port map( B1 => n15381, B2 => n21026, C1 => n15243, C2 =>
                           n21034, A => n18934, ZN => n18933);
   U15356 : NOR4_X1 port map( A1 => n18893, A2 => n18894, A3 => n18895, A4 => 
                           n18896, ZN => n18892);
   U15357 : OAI221_X1 port map( B1 => n16218, B2 => n20859, C1 => n16112, C2 =>
                           n20873, A => n18900, ZN => n18893);
   U15358 : OAI221_X1 port map( B1 => n8097, B2 => n20792, C1 => n16533, C2 => 
                           n20729, A => n18899, ZN => n18894);
   U15359 : OAI221_X1 port map( B1 => n15659, B2 => n20981, C1 => n15765, C2 =>
                           n20987, A => n18898, ZN => n18895);
   U15360 : NOR4_X1 port map( A1 => n17516, A2 => n17517, A3 => n17518, A4 => 
                           n17519, ZN => n17515);
   U15361 : OAI221_X1 port map( B1 => n16220, B2 => n21420, C1 => n16114, C2 =>
                           n21430, A => n17525, ZN => n17516);
   U15362 : OAI221_X1 port map( B1 => n8033, B2 => n21353, C1 => n16535, C2 => 
                           n21286, A => n17524, ZN => n17517);
   U15363 : OAI221_X1 port map( B1 => n15382, B2 => n21587, C1 => n15244, C2 =>
                           n21589, A => n17520, ZN => n17519);
   U15364 : NOR4_X1 port map( A1 => n17469, A2 => n17470, A3 => n17471, A4 => 
                           n17472, ZN => n17468);
   U15365 : OAI221_X1 port map( B1 => n16219, B2 => n21416, C1 => n16113, C2 =>
                           n21432, A => n17478, ZN => n17469);
   U15366 : OAI221_X1 port map( B1 => n8065, B2 => n21349, C1 => n16534, C2 => 
                           n21288, A => n17477, ZN => n17470);
   U15367 : OAI221_X1 port map( B1 => n15381, B2 => n21583, C1 => n15243, C2 =>
                           n21591, A => n17473, ZN => n17472);
   U15368 : NOR4_X1 port map( A1 => n17422, A2 => n17423, A3 => n17424, A4 => 
                           n17425, ZN => n17421);
   U15369 : OAI221_X1 port map( B1 => n16218, B2 => n21416, C1 => n16112, C2 =>
                           n21430, A => n17431, ZN => n17422);
   U15370 : OAI221_X1 port map( B1 => n8097, B2 => n21349, C1 => n16533, C2 => 
                           n21286, A => n17430, ZN => n17423);
   U15371 : OAI221_X1 port map( B1 => n15659, B2 => n21538, C1 => n15765, C2 =>
                           n21544, A => n17428, ZN => n17424);
   U15372 : NOR4_X1 port map( A1 => n18856, A2 => n18857, A3 => n18858, A4 => 
                           n18859, ZN => n18855);
   U15373 : OAI221_X1 port map( B1 => n16217, B2 => n20861, C1 => n16111, C2 =>
                           n20878, A => n18863, ZN => n18856);
   U15374 : OAI221_X1 port map( B1 => n8129, B2 => n20794, C1 => n16532, C2 => 
                           n20734, A => n18862, ZN => n18857);
   U15375 : OAI221_X1 port map( B1 => n15379, B2 => n21028, C1 => n15241, C2 =>
                           n21037, A => n18860, ZN => n18859);
   U15376 : NOR4_X1 port map( A1 => n17375, A2 => n17376, A3 => n17377, A4 => 
                           n17378, ZN => n17374);
   U15377 : OAI221_X1 port map( B1 => n16217, B2 => n21418, C1 => n16111, C2 =>
                           n21435, A => n17384, ZN => n17375);
   U15378 : OAI221_X1 port map( B1 => n8129, B2 => n21351, C1 => n16532, C2 => 
                           n21291, A => n17383, ZN => n17376);
   U15379 : OAI221_X1 port map( B1 => n15379, B2 => n21585, C1 => n15241, C2 =>
                           n21594, A => n17379, ZN => n17378);
   U15380 : NOR2_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), ZN => n15228);
   U15381 : AOI221_X1 port map( B1 => n20866, B2 => n8905, C1 => n20881, C2 => 
                           n19723, A => n19612, ZN => n19591);
   U15382 : OAI22_X1 port map( A1 => n16202, A2 => n20888, B1 => n16340, B2 => 
                           n20896, ZN => n19612);
   U15383 : AOI221_X1 port map( B1 => n21112, B2 => n9468, C1 => n21121, C2 => 
                           n19724, A => n19586, ZN => n19583);
   U15384 : OAI22_X1 port map( A1 => n16518, A2 => n21135, B1 => n15853, B2 => 
                           n21132, ZN => n19586);
   U15385 : AOI221_X1 port map( B1 => n20866, B2 => n8894, C1 => n20881, C2 => 
                           n19725, A => n19575, ZN => n19554);
   U15386 : OAI22_X1 port map( A1 => n16201, A2 => n20888, B1 => n16339, B2 => 
                           n20901, ZN => n19575);
   U15387 : AOI221_X1 port map( B1 => n21117, B2 => n9467, C1 => n21120, C2 => 
                           n19726, A => n19549, ZN => n19546);
   U15388 : OAI22_X1 port map( A1 => n16517, A2 => n21139, B1 => n15852, B2 => 
                           n21127, ZN => n19549);
   U15389 : AOI221_X1 port map( B1 => n20868, B2 => n8883, C1 => n20882, C2 => 
                           n19727, A => n19538, ZN => n19517);
   U15390 : OAI22_X1 port map( A1 => n16200, A2 => n20893, B1 => n16338, B2 => 
                           n20896, ZN => n19538);
   U15391 : AOI221_X1 port map( B1 => n21116, B2 => n9466, C1 => n21120, C2 => 
                           n19728, A => n19512, ZN => n19509);
   U15392 : OAI22_X1 port map( A1 => n16516, A2 => n21135, B1 => n15851, B2 => 
                           n21127, ZN => n19512);
   U15393 : AOI221_X1 port map( B1 => n20867, B2 => n8872, C1 => n20882, C2 => 
                           n19729, A => n19501, ZN => n19480);
   U15394 : OAI22_X1 port map( A1 => n16199, A2 => n20888, B1 => n16337, B2 => 
                           n20896, ZN => n19501);
   U15395 : AOI221_X1 port map( B1 => n21112, B2 => n9465, C1 => n21125, C2 => 
                           n19730, A => n19475, ZN => n19472);
   U15396 : OAI22_X1 port map( A1 => n16515, A2 => n21136, B1 => n15850, B2 => 
                           n21128, ZN => n19475);
   U15397 : AOI221_X1 port map( B1 => n20868, B2 => n8861, C1 => n20882, C2 => 
                           n19731, A => n19464, ZN => n19443);
   U15398 : OAI22_X1 port map( A1 => n16198, A2 => n20889, B1 => n16336, B2 => 
                           n20897, ZN => n19464);
   U15399 : AOI221_X1 port map( B1 => n21114, B2 => n9464, C1 => n21121, C2 => 
                           n19732, A => n19438, ZN => n19435);
   U15400 : OAI22_X1 port map( A1 => n16514, A2 => n21136, B1 => n15849, B2 => 
                           n21129, ZN => n19438);
   U15401 : AOI221_X1 port map( B1 => n20868, B2 => n8850, C1 => n20883, C2 => 
                           n19733, A => n19427, ZN => n19406);
   U15402 : OAI22_X1 port map( A1 => n16197, A2 => n20889, B1 => n16335, B2 => 
                           n20898, ZN => n19427);
   U15403 : AOI221_X1 port map( B1 => n21115, B2 => n9463, C1 => n21122, C2 => 
                           n19734, A => n19401, ZN => n19398);
   U15404 : OAI22_X1 port map( A1 => n16513, A2 => n21137, B1 => n15848, B2 => 
                           n21130, ZN => n19401);
   U15405 : AOI221_X1 port map( B1 => n20869, B2 => n8839, C1 => n20884, C2 => 
                           n19735, A => n19390, ZN => n19369);
   U15406 : OAI22_X1 port map( A1 => n16196, A2 => n20890, B1 => n16334, B2 => 
                           n20897, ZN => n19390);
   U15407 : AOI221_X1 port map( B1 => n21113, B2 => n9462, C1 => n21122, C2 => 
                           n19736, A => n19364, ZN => n19361);
   U15408 : OAI22_X1 port map( A1 => n16512, A2 => n21138, B1 => n15847, B2 => 
                           n21131, ZN => n19364);
   U15409 : AOI221_X1 port map( B1 => n20869, B2 => n8828, C1 => n20883, C2 => 
                           n19737, A => n19353, ZN => n19332);
   U15410 : OAI22_X1 port map( A1 => n16195, A2 => n20890, B1 => n16333, B2 => 
                           n20902, ZN => n19353);
   U15411 : AOI221_X1 port map( B1 => n21113, B2 => n9461, C1 => n21123, C2 => 
                           n19738, A => n19327, ZN => n19324);
   U15412 : OAI22_X1 port map( A1 => n16511, A2 => n21138, B1 => n15846, B2 => 
                           n21131, ZN => n19327);
   U15413 : AOI221_X1 port map( B1 => n20871, B2 => n8817, C1 => n20886, C2 => 
                           n19739, A => n19316, ZN => n19295);
   U15414 : OAI22_X1 port map( A1 => n16194, A2 => n20888, B1 => n16332, B2 => 
                           n20899, ZN => n19316);
   U15415 : AOI221_X1 port map( B1 => n21113, B2 => n9460, C1 => n21123, C2 => 
                           n19740, A => n19290, ZN => n19287);
   U15416 : OAI22_X1 port map( A1 => n16510, A2 => n21137, B1 => n15845, B2 => 
                           n21130, ZN => n19290);
   U15417 : AOI221_X1 port map( B1 => n20870, B2 => n8806, C1 => n20883, C2 => 
                           n19741, A => n19279, ZN => n19258);
   U15418 : OAI22_X1 port map( A1 => n16193, A2 => n20891, B1 => n16331, B2 => 
                           n20899, ZN => n19279);
   U15419 : AOI221_X1 port map( B1 => n21114, B2 => n9459, C1 => n21124, C2 => 
                           n19742, A => n19253, ZN => n19250);
   U15420 : OAI22_X1 port map( A1 => n16509, A2 => n21136, B1 => n15844, B2 => 
                           n21128, ZN => n19253);
   U15421 : AOI221_X1 port map( B1 => n20871, B2 => n8795, C1 => n20884, C2 => 
                           n19743, A => n19242, ZN => n19221);
   U15422 : OAI22_X1 port map( A1 => n16192, A2 => n20892, B1 => n16330, B2 => 
                           n20900, ZN => n19242);
   U15423 : AOI221_X1 port map( B1 => n21115, B2 => n9458, C1 => n21124, C2 => 
                           n19744, A => n19216, ZN => n19213);
   U15424 : OAI22_X1 port map( A1 => n16508, A2 => n21139, B1 => n15843, B2 => 
                           n21132, ZN => n19216);
   U15425 : AOI221_X1 port map( B1 => n20871, B2 => n8784, C1 => n20885, C2 => 
                           n19745, A => n19205, ZN => n19184);
   U15426 : OAI22_X1 port map( A1 => n16191, A2 => n20889, B1 => n16329, B2 => 
                           n20897, ZN => n19205);
   U15427 : AOI221_X1 port map( B1 => n21115, B2 => n9457, C1 => n21124, C2 => 
                           n19746, A => n19179, ZN => n19176);
   U15428 : OAI22_X1 port map( A1 => n16507, A2 => n21136, B1 => n15842, B2 => 
                           n21129, ZN => n19179);
   U15429 : AOI221_X1 port map( B1 => n20867, B2 => n8773, C1 => n20885, C2 => 
                           n19747, A => n19168, ZN => n19147);
   U15430 : OAI22_X1 port map( A1 => n16190, A2 => n20890, B1 => n16328, B2 => 
                           n20897, ZN => n19168);
   U15431 : AOI221_X1 port map( B1 => n21116, B2 => n9456, C1 => n21123, C2 => 
                           n19748, A => n19142, ZN => n19139);
   U15432 : OAI22_X1 port map( A1 => n16506, A2 => n21137, B1 => n15841, B2 => 
                           n21130, ZN => n19142);
   U15433 : AOI221_X1 port map( B1 => n20870, B2 => n8762, C1 => n20885, C2 => 
                           n19749, A => n19131, ZN => n19110);
   U15434 : OAI22_X1 port map( A1 => n16189, A2 => n20889, B1 => n16327, B2 => 
                           n20898, ZN => n19131);
   U15435 : AOI221_X1 port map( B1 => n21115, B2 => n9455, C1 => n21124, C2 => 
                           n19750, A => n19105, ZN => n19102);
   U15436 : OAI22_X1 port map( A1 => n16505, A2 => n21137, B1 => n15840, B2 => 
                           n21130, ZN => n19105);
   U15437 : AOI221_X1 port map( B1 => n20871, B2 => n8751, C1 => n20884, C2 => 
                           n19751, A => n19094, ZN => n19073);
   U15438 : OAI22_X1 port map( A1 => n16188, A2 => n20890, B1 => n16326, B2 => 
                           n20898, ZN => n19094);
   U15439 : AOI221_X1 port map( B1 => n21114, B2 => n9454, C1 => n21124, C2 => 
                           n19752, A => n19068, ZN => n19065);
   U15440 : OAI22_X1 port map( A1 => n16504, A2 => n21138, B1 => n15839, B2 => 
                           n21131, ZN => n19068);
   U15441 : AOI221_X1 port map( B1 => n20869, B2 => n8740, C1 => n20885, C2 => 
                           n19753, A => n19057, ZN => n19036);
   U15442 : OAI22_X1 port map( A1 => n16187, A2 => n20889, B1 => n16325, B2 => 
                           n20898, ZN => n19057);
   U15443 : AOI221_X1 port map( B1 => n21116, B2 => n9453, C1 => n21121, C2 => 
                           n19754, A => n19031, ZN => n19028);
   U15444 : OAI22_X1 port map( A1 => n16503, A2 => n21138, B1 => n15838, B2 => 
                           n21131, ZN => n19031);
   U15445 : AOI221_X1 port map( B1 => n20870, B2 => n8729, C1 => n20885, C2 => 
                           n19755, A => n19020, ZN => n18999);
   U15446 : OAI22_X1 port map( A1 => n16186, A2 => n20892, B1 => n16324, B2 => 
                           n20900, ZN => n19020);
   U15447 : AOI221_X1 port map( B1 => n21116, B2 => n9452, C1 => n21120, C2 => 
                           n19756, A => n18994, ZN => n18991);
   U15448 : OAI22_X1 port map( A1 => n16502, A2 => n21135, B1 => n15837, B2 => 
                           n21133, ZN => n18994);
   U15449 : AOI221_X1 port map( B1 => n20872, B2 => n8718, C1 => n20886, C2 => 
                           n19757, A => n18983, ZN => n18962);
   U15450 : OAI22_X1 port map( A1 => n16185, A2 => n20891, B1 => n16323, B2 => 
                           n20899, ZN => n18983);
   U15451 : AOI221_X1 port map( B1 => n21113, B2 => n9451, C1 => n21123, C2 => 
                           n19758, A => n18957, ZN => n18954);
   U15452 : OAI22_X1 port map( A1 => n16501, A2 => n21139, B1 => n15836, B2 => 
                           n21132, ZN => n18957);
   U15453 : AOI221_X1 port map( B1 => n20872, B2 => n8707, C1 => n20886, C2 => 
                           n19759, A => n18946, ZN => n18925);
   U15454 : OAI22_X1 port map( A1 => n16184, A2 => n20892, B1 => n16322, B2 => 
                           n20899, ZN => n18946);
   U15455 : AOI221_X1 port map( B1 => n21116, B2 => n9450, C1 => n21122, C2 => 
                           n19760, A => n18920, ZN => n18917);
   U15456 : OAI22_X1 port map( A1 => n16500, A2 => n21140, B1 => n15835, B2 => 
                           n21131, ZN => n18920);
   U15457 : AOI221_X1 port map( B1 => n21117, B2 => n9449, C1 => n21125, C2 => 
                           n19761, A => n18883, ZN => n18880);
   U15458 : OAI22_X1 port map( A1 => n16499, A2 => n21135, B1 => n15834, B2 => 
                           n21127, ZN => n18883);
   U15459 : AOI221_X1 port map( B1 => n21117, B2 => n9448, C1 => n21125, C2 => 
                           n19762, A => n18846, ZN => n18843);
   U15460 : OAI22_X1 port map( A1 => n16498, A2 => n21140, B1 => n15833, B2 => 
                           n21132, ZN => n18846);
   U15461 : AOI221_X1 port map( B1 => n20868, B2 => n8608, C1 => n20883, C2 => 
                           n19763, A => n18613, ZN => n18592);
   U15462 : OAI22_X1 port map( A1 => n16175, A2 => n20891, B1 => n16313, B2 => 
                           n20896, ZN => n18613);
   U15463 : AOI221_X1 port map( B1 => n20869, B2 => n8597, C1 => n20884, C2 => 
                           n19764, A => n18576, ZN => n18555);
   U15464 : OAI22_X1 port map( A1 => n16174, A2 => n20888, B1 => n16312, B2 => 
                           n20896, ZN => n18576);
   U15465 : AOI221_X1 port map( B1 => n20868, B2 => n8586, C1 => n20883, C2 => 
                           n19765, A => n18539, ZN => n18518);
   U15466 : OAI22_X1 port map( A1 => n16173, A2 => n20888, B1 => n16311, B2 => 
                           n20902, ZN => n18539);
   U15467 : AOI221_X1 port map( B1 => n21113, B2 => n9439, C1 => n21122, C2 => 
                           n19766, A => n18513, ZN => n18510);
   U15468 : OAI22_X1 port map( A1 => n16489, A2 => n21136, B1 => n15824, B2 => 
                           n21133, ZN => n18513);
   U15469 : AOI221_X1 port map( B1 => n20870, B2 => n8575, C1 => n20884, C2 => 
                           n19767, A => n18492, ZN => n18448);
   U15470 : OAI22_X1 port map( A1 => n16172, A2 => n20894, B1 => n16310, B2 => 
                           n20896, ZN => n18492);
   U15471 : AOI221_X1 port map( B1 => n21114, B2 => n9438, C1 => n21122, C2 => 
                           n19768, A => n18433, ZN => n18423);
   U15472 : OAI22_X1 port map( A1 => n16488, A2 => n21140, B1 => n15823, B2 => 
                           n21129, ZN => n18433);
   U15473 : AOI221_X1 port map( B1 => n21423, B2 => n8905, C1 => n21438, C2 => 
                           n19723, A => n18338, ZN => n18309);
   U15474 : OAI22_X1 port map( A1 => n16202, A2 => n21445, B1 => n16340, B2 => 
                           n21453, ZN => n18338);
   U15475 : AOI221_X1 port map( B1 => n21669, B2 => n9468, C1 => n21678, C2 => 
                           n19724, A => n18304, ZN => n18300);
   U15476 : OAI22_X1 port map( A1 => n16518, A2 => n21692, B1 => n15853, B2 => 
                           n21689, ZN => n18304);
   U15477 : AOI221_X1 port map( B1 => n21423, B2 => n8894, C1 => n21438, C2 => 
                           n19725, A => n18291, ZN => n18262);
   U15478 : OAI22_X1 port map( A1 => n16201, A2 => n21445, B1 => n16339, B2 => 
                           n21458, ZN => n18291);
   U15479 : AOI221_X1 port map( B1 => n21674, B2 => n9467, C1 => n21677, C2 => 
                           n19726, A => n18257, ZN => n18253);
   U15480 : OAI22_X1 port map( A1 => n16517, A2 => n21696, B1 => n15852, B2 => 
                           n21684, ZN => n18257);
   U15481 : AOI221_X1 port map( B1 => n21425, B2 => n8883, C1 => n21439, C2 => 
                           n19727, A => n18244, ZN => n18215);
   U15482 : OAI22_X1 port map( A1 => n16200, A2 => n21450, B1 => n16338, B2 => 
                           n21453, ZN => n18244);
   U15483 : AOI221_X1 port map( B1 => n21673, B2 => n9466, C1 => n21677, C2 => 
                           n19728, A => n18210, ZN => n18206);
   U15484 : OAI22_X1 port map( A1 => n16516, A2 => n21692, B1 => n15851, B2 => 
                           n21684, ZN => n18210);
   U15485 : AOI221_X1 port map( B1 => n21424, B2 => n8872, C1 => n21439, C2 => 
                           n19729, A => n18197, ZN => n18168);
   U15486 : OAI22_X1 port map( A1 => n16199, A2 => n21445, B1 => n16337, B2 => 
                           n21453, ZN => n18197);
   U15487 : AOI221_X1 port map( B1 => n21669, B2 => n9465, C1 => n21682, C2 => 
                           n19730, A => n18163, ZN => n18159);
   U15488 : OAI22_X1 port map( A1 => n16515, A2 => n21693, B1 => n15850, B2 => 
                           n21685, ZN => n18163);
   U15489 : AOI221_X1 port map( B1 => n21425, B2 => n8861, C1 => n21439, C2 => 
                           n19731, A => n18150, ZN => n18121);
   U15490 : OAI22_X1 port map( A1 => n16198, A2 => n21446, B1 => n16336, B2 => 
                           n21454, ZN => n18150);
   U15491 : AOI221_X1 port map( B1 => n21671, B2 => n9464, C1 => n21678, C2 => 
                           n19732, A => n18116, ZN => n18112);
   U15492 : OAI22_X1 port map( A1 => n16514, A2 => n21693, B1 => n15849, B2 => 
                           n21686, ZN => n18116);
   U15493 : AOI221_X1 port map( B1 => n21425, B2 => n8850, C1 => n21440, C2 => 
                           n19733, A => n18103, ZN => n18074);
   U15494 : OAI22_X1 port map( A1 => n16197, A2 => n21446, B1 => n16335, B2 => 
                           n21455, ZN => n18103);
   U15495 : AOI221_X1 port map( B1 => n21672, B2 => n9463, C1 => n21679, C2 => 
                           n19734, A => n18069, ZN => n18065);
   U15496 : OAI22_X1 port map( A1 => n16513, A2 => n21694, B1 => n15848, B2 => 
                           n21687, ZN => n18069);
   U15497 : AOI221_X1 port map( B1 => n21426, B2 => n8839, C1 => n21441, C2 => 
                           n19735, A => n18056, ZN => n18027);
   U15498 : OAI22_X1 port map( A1 => n16196, A2 => n21447, B1 => n16334, B2 => 
                           n21454, ZN => n18056);
   U15499 : AOI221_X1 port map( B1 => n21670, B2 => n9462, C1 => n21679, C2 => 
                           n19736, A => n18022, ZN => n18018);
   U15500 : OAI22_X1 port map( A1 => n16512, A2 => n21695, B1 => n15847, B2 => 
                           n21688, ZN => n18022);
   U15501 : AOI221_X1 port map( B1 => n21426, B2 => n8828, C1 => n21440, C2 => 
                           n19737, A => n18009, ZN => n17980);
   U15502 : OAI22_X1 port map( A1 => n16195, A2 => n21447, B1 => n16333, B2 => 
                           n21459, ZN => n18009);
   U15503 : AOI221_X1 port map( B1 => n21670, B2 => n9461, C1 => n21680, C2 => 
                           n19738, A => n17975, ZN => n17971);
   U15504 : OAI22_X1 port map( A1 => n16511, A2 => n21695, B1 => n15846, B2 => 
                           n21688, ZN => n17975);
   U15505 : AOI221_X1 port map( B1 => n21428, B2 => n8817, C1 => n21443, C2 => 
                           n19739, A => n17962, ZN => n17933);
   U15506 : OAI22_X1 port map( A1 => n16194, A2 => n21445, B1 => n16332, B2 => 
                           n21456, ZN => n17962);
   U15507 : AOI221_X1 port map( B1 => n21670, B2 => n9460, C1 => n21680, C2 => 
                           n19740, A => n17928, ZN => n17924);
   U15508 : OAI22_X1 port map( A1 => n16510, A2 => n21694, B1 => n15845, B2 => 
                           n21687, ZN => n17928);
   U15509 : AOI221_X1 port map( B1 => n21427, B2 => n8806, C1 => n21440, C2 => 
                           n19741, A => n17915, ZN => n17886);
   U15510 : OAI22_X1 port map( A1 => n16193, A2 => n21448, B1 => n16331, B2 => 
                           n21456, ZN => n17915);
   U15511 : AOI221_X1 port map( B1 => n21671, B2 => n9459, C1 => n21681, C2 => 
                           n19742, A => n17881, ZN => n17877);
   U15512 : OAI22_X1 port map( A1 => n16509, A2 => n21693, B1 => n15844, B2 => 
                           n21685, ZN => n17881);
   U15513 : AOI221_X1 port map( B1 => n21428, B2 => n8795, C1 => n21441, C2 => 
                           n19743, A => n17868, ZN => n17839);
   U15514 : OAI22_X1 port map( A1 => n16192, A2 => n21449, B1 => n16330, B2 => 
                           n21457, ZN => n17868);
   U15515 : AOI221_X1 port map( B1 => n21672, B2 => n9458, C1 => n21681, C2 => 
                           n19744, A => n17834, ZN => n17830);
   U15516 : OAI22_X1 port map( A1 => n16508, A2 => n21696, B1 => n15843, B2 => 
                           n21689, ZN => n17834);
   U15517 : AOI221_X1 port map( B1 => n21428, B2 => n8784, C1 => n21442, C2 => 
                           n19745, A => n17821, ZN => n17792);
   U15518 : OAI22_X1 port map( A1 => n16191, A2 => n21446, B1 => n16329, B2 => 
                           n21454, ZN => n17821);
   U15519 : AOI221_X1 port map( B1 => n21672, B2 => n9457, C1 => n21681, C2 => 
                           n19746, A => n17787, ZN => n17783);
   U15520 : OAI22_X1 port map( A1 => n16507, A2 => n21693, B1 => n15842, B2 => 
                           n21686, ZN => n17787);
   U15521 : AOI221_X1 port map( B1 => n21424, B2 => n8773, C1 => n21442, C2 => 
                           n19747, A => n17774, ZN => n17745);
   U15522 : OAI22_X1 port map( A1 => n16190, A2 => n21447, B1 => n16328, B2 => 
                           n21454, ZN => n17774);
   U15523 : AOI221_X1 port map( B1 => n21673, B2 => n9456, C1 => n21680, C2 => 
                           n19748, A => n17740, ZN => n17736);
   U15524 : OAI22_X1 port map( A1 => n16506, A2 => n21694, B1 => n15841, B2 => 
                           n21687, ZN => n17740);
   U15525 : AOI221_X1 port map( B1 => n21427, B2 => n8762, C1 => n21442, C2 => 
                           n19749, A => n17727, ZN => n17698);
   U15526 : OAI22_X1 port map( A1 => n16189, A2 => n21446, B1 => n16327, B2 => 
                           n21455, ZN => n17727);
   U15527 : AOI221_X1 port map( B1 => n21672, B2 => n9455, C1 => n21681, C2 => 
                           n19750, A => n17693, ZN => n17689);
   U15528 : OAI22_X1 port map( A1 => n16505, A2 => n21694, B1 => n15840, B2 => 
                           n21687, ZN => n17693);
   U15529 : AOI221_X1 port map( B1 => n21428, B2 => n8751, C1 => n21441, C2 => 
                           n19751, A => n17680, ZN => n17651);
   U15530 : OAI22_X1 port map( A1 => n16188, A2 => n21447, B1 => n16326, B2 => 
                           n21455, ZN => n17680);
   U15531 : AOI221_X1 port map( B1 => n21671, B2 => n9454, C1 => n21681, C2 => 
                           n19752, A => n17646, ZN => n17642);
   U15532 : OAI22_X1 port map( A1 => n16504, A2 => n21695, B1 => n15839, B2 => 
                           n21688, ZN => n17646);
   U15533 : AOI221_X1 port map( B1 => n21426, B2 => n8740, C1 => n21442, C2 => 
                           n19753, A => n17633, ZN => n17604);
   U15534 : OAI22_X1 port map( A1 => n16187, A2 => n21446, B1 => n16325, B2 => 
                           n21455, ZN => n17633);
   U15535 : AOI221_X1 port map( B1 => n21673, B2 => n9453, C1 => n21678, C2 => 
                           n19754, A => n17599, ZN => n17595);
   U15536 : OAI22_X1 port map( A1 => n16503, A2 => n21695, B1 => n15838, B2 => 
                           n21688, ZN => n17599);
   U15537 : AOI221_X1 port map( B1 => n21427, B2 => n8729, C1 => n21442, C2 => 
                           n19755, A => n17586, ZN => n17557);
   U15538 : OAI22_X1 port map( A1 => n16186, A2 => n21449, B1 => n16324, B2 => 
                           n21457, ZN => n17586);
   U15539 : AOI221_X1 port map( B1 => n21673, B2 => n9452, C1 => n21677, C2 => 
                           n19756, A => n17552, ZN => n17548);
   U15540 : OAI22_X1 port map( A1 => n16502, A2 => n21692, B1 => n15837, B2 => 
                           n21690, ZN => n17552);
   U15541 : AOI221_X1 port map( B1 => n21429, B2 => n8718, C1 => n21443, C2 => 
                           n19757, A => n17539, ZN => n17510);
   U15542 : OAI22_X1 port map( A1 => n16185, A2 => n21448, B1 => n16323, B2 => 
                           n21456, ZN => n17539);
   U15543 : AOI221_X1 port map( B1 => n21670, B2 => n9451, C1 => n21680, C2 => 
                           n19758, A => n17505, ZN => n17501);
   U15544 : OAI22_X1 port map( A1 => n16501, A2 => n21696, B1 => n15836, B2 => 
                           n21689, ZN => n17505);
   U15545 : AOI221_X1 port map( B1 => n21429, B2 => n8707, C1 => n21443, C2 => 
                           n19759, A => n17492, ZN => n17463);
   U15546 : OAI22_X1 port map( A1 => n16184, A2 => n21449, B1 => n16322, B2 => 
                           n21456, ZN => n17492);
   U15547 : AOI221_X1 port map( B1 => n21673, B2 => n9450, C1 => n21679, C2 => 
                           n19760, A => n17458, ZN => n17454);
   U15548 : OAI22_X1 port map( A1 => n16500, A2 => n21697, B1 => n15835, B2 => 
                           n21688, ZN => n17458);
   U15549 : AOI221_X1 port map( B1 => n21674, B2 => n9449, C1 => n21682, C2 => 
                           n19761, A => n17411, ZN => n17407);
   U15550 : OAI22_X1 port map( A1 => n16499, A2 => n21692, B1 => n15834, B2 => 
                           n21684, ZN => n17411);
   U15551 : AOI221_X1 port map( B1 => n21674, B2 => n9448, C1 => n21682, C2 => 
                           n19762, A => n17364, ZN => n17360);
   U15552 : OAI22_X1 port map( A1 => n16498, A2 => n21697, B1 => n15833, B2 => 
                           n21689, ZN => n17364);
   U15553 : AOI221_X1 port map( B1 => n21425, B2 => n8608, C1 => n21440, C2 => 
                           n19763, A => n17069, ZN => n17040);
   U15554 : OAI22_X1 port map( A1 => n16175, A2 => n21448, B1 => n16313, B2 => 
                           n21453, ZN => n17069);
   U15555 : AOI221_X1 port map( B1 => n21426, B2 => n8597, C1 => n21441, C2 => 
                           n19764, A => n17022, ZN => n16993);
   U15556 : OAI22_X1 port map( A1 => n16174, A2 => n21445, B1 => n16312, B2 => 
                           n21453, ZN => n17022);
   U15557 : AOI221_X1 port map( B1 => n21425, B2 => n8586, C1 => n21440, C2 => 
                           n19765, A => n16975, ZN => n16946);
   U15558 : OAI22_X1 port map( A1 => n16173, A2 => n21445, B1 => n16311, B2 => 
                           n21459, ZN => n16975);
   U15559 : AOI221_X1 port map( B1 => n21670, B2 => n9439, C1 => n21679, C2 => 
                           n19766, A => n16941, ZN => n16937);
   U15560 : OAI22_X1 port map( A1 => n16489, A2 => n21693, B1 => n15824, B2 => 
                           n21690, ZN => n16941);
   U15561 : AOI221_X1 port map( B1 => n21427, B2 => n8575, C1 => n21441, C2 => 
                           n19767, A => n16918, ZN => n16866);
   U15562 : OAI22_X1 port map( A1 => n16172, A2 => n21451, B1 => n16310, B2 => 
                           n21453, ZN => n16918);
   U15563 : AOI221_X1 port map( B1 => n21671, B2 => n9438, C1 => n21679, C2 => 
                           n19768, A => n16851, ZN => n16840);
   U15564 : OAI22_X1 port map( A1 => n16488, A2 => n21697, B1 => n15823, B2 => 
                           n21686, ZN => n16851);
   U15565 : AOI221_X1 port map( B1 => n20872, B2 => n8696, C1 => n20886, C2 => 
                           n19682, A => n18909, ZN => n18888);
   U15566 : OAI22_X1 port map( A1 => n16183, A2 => n20892, B1 => n16321, B2 => 
                           n20900, ZN => n18909);
   U15567 : AOI221_X1 port map( B1 => n20872, B2 => n8685, C1 => n20886, C2 => 
                           n19683, A => n18872, ZN => n18851);
   U15568 : OAI22_X1 port map( A1 => n16182, A2 => n20891, B1 => n16320, B2 => 
                           n20900, ZN => n18872);
   U15569 : AOI221_X1 port map( B1 => n20866, B2 => n8674, C1 => n20881, C2 => 
                           n19769, A => n18835, ZN => n18814);
   U15570 : OAI22_X1 port map( A1 => n16181, A2 => n20893, B1 => n16319, B2 => 
                           n20902, ZN => n18835);
   U15571 : AOI221_X1 port map( B1 => n21117, B2 => n9447, C1 => n21125, C2 => 
                           n19684, A => n18809, ZN => n18806);
   U15572 : OAI22_X1 port map( A1 => n16497, A2 => n21139, B1 => n15832, B2 => 
                           n21130, ZN => n18809);
   U15573 : AOI221_X1 port map( B1 => n20866, B2 => n8663, C1 => n20881, C2 => 
                           n19770, A => n18798, ZN => n18777);
   U15574 : OAI22_X1 port map( A1 => n16180, A2 => n20893, B1 => n16318, B2 => 
                           n20901, ZN => n18798);
   U15575 : AOI221_X1 port map( B1 => n21117, B2 => n9446, C1 => n21125, C2 => 
                           n19685, A => n18772, ZN => n18769);
   U15576 : OAI22_X1 port map( A1 => n16496, A2 => n21140, B1 => n15831, B2 => 
                           n21132, ZN => n18772);
   U15577 : AOI221_X1 port map( B1 => n20866, B2 => n8652, C1 => n20881, C2 => 
                           n19771, A => n18761, ZN => n18740);
   U15578 : OAI22_X1 port map( A1 => n16179, A2 => n20894, B1 => n16317, B2 => 
                           n20902, ZN => n18761);
   U15579 : AOI221_X1 port map( B1 => n21112, B2 => n9445, C1 => n21121, C2 => 
                           n19772, A => n18735, ZN => n18732);
   U15580 : OAI22_X1 port map( A1 => n16495, A2 => n21138, B1 => n15830, B2 => 
                           n21128, ZN => n18735);
   U15581 : AOI221_X1 port map( B1 => n20872, B2 => n8641, C1 => n20882, C2 => 
                           n19773, A => n18724, ZN => n18703);
   U15582 : OAI22_X1 port map( A1 => n16178, A2 => n20894, B1 => n16316, B2 => 
                           n20901, ZN => n18724);
   U15583 : AOI221_X1 port map( B1 => n21117, B2 => n9444, C1 => n21120, C2 => 
                           n19774, A => n18698, ZN => n18695);
   U15584 : OAI22_X1 port map( A1 => n16494, A2 => n21141, B1 => n15829, B2 => 
                           n21127, ZN => n18698);
   U15585 : AOI221_X1 port map( B1 => n20867, B2 => n8630, C1 => n20882, C2 => 
                           n19775, A => n18687, ZN => n18666);
   U15586 : OAI22_X1 port map( A1 => n16177, A2 => n20893, B1 => n16315, B2 => 
                           n20902, ZN => n18687);
   U15587 : AOI221_X1 port map( B1 => n21112, B2 => n9443, C1 => n21120, C2 => 
                           n19776, A => n18661, ZN => n18658);
   U15588 : OAI22_X1 port map( A1 => n16493, A2 => n21140, B1 => n15828, B2 => 
                           n21133, ZN => n18661);
   U15589 : AOI221_X1 port map( B1 => n20867, B2 => n8619, C1 => n20882, C2 => 
                           n19777, A => n18650, ZN => n18629);
   U15590 : OAI22_X1 port map( A1 => n16176, A2 => n20894, B1 => n16314, B2 => 
                           n20901, ZN => n18650);
   U15591 : AOI221_X1 port map( B1 => n21112, B2 => n9442, C1 => n21123, C2 => 
                           n19778, A => n18624, ZN => n18621);
   U15592 : OAI22_X1 port map( A1 => n16492, A2 => n21135, B1 => n15827, B2 => 
                           n21133, ZN => n18624);
   U15593 : AOI221_X1 port map( B1 => n21113, B2 => n9441, C1 => n21121, C2 => 
                           n19779, A => n18587, ZN => n18584);
   U15594 : OAI22_X1 port map( A1 => n16491, A2 => n21141, B1 => n15826, B2 => 
                           n21133, ZN => n18587);
   U15595 : AOI221_X1 port map( B1 => n21114, B2 => n9440, C1 => n21121, C2 => 
                           n19780, A => n18550, ZN => n18547);
   U15596 : OAI22_X1 port map( A1 => n16490, A2 => n21141, B1 => n15825, B2 => 
                           n21129, ZN => n18550);
   U15597 : AOI221_X1 port map( B1 => n21429, B2 => n8696, C1 => n21443, C2 => 
                           n19682, A => n17445, ZN => n17416);
   U15598 : OAI22_X1 port map( A1 => n16183, A2 => n21449, B1 => n16321, B2 => 
                           n21457, ZN => n17445);
   U15599 : AOI221_X1 port map( B1 => n21429, B2 => n8685, C1 => n21443, C2 => 
                           n19683, A => n17398, ZN => n17369);
   U15600 : OAI22_X1 port map( A1 => n16182, A2 => n21448, B1 => n16320, B2 => 
                           n21457, ZN => n17398);
   U15601 : AOI221_X1 port map( B1 => n21423, B2 => n8674, C1 => n21438, C2 => 
                           n19769, A => n17351, ZN => n17322);
   U15602 : OAI22_X1 port map( A1 => n16181, A2 => n21450, B1 => n16319, B2 => 
                           n21459, ZN => n17351);
   U15603 : AOI221_X1 port map( B1 => n21674, B2 => n9447, C1 => n21682, C2 => 
                           n19684, A => n17317, ZN => n17313);
   U15604 : OAI22_X1 port map( A1 => n16497, A2 => n21696, B1 => n15832, B2 => 
                           n21687, ZN => n17317);
   U15605 : AOI221_X1 port map( B1 => n21423, B2 => n8663, C1 => n21438, C2 => 
                           n19770, A => n17304, ZN => n17275);
   U15606 : OAI22_X1 port map( A1 => n16180, A2 => n21450, B1 => n16318, B2 => 
                           n21458, ZN => n17304);
   U15607 : AOI221_X1 port map( B1 => n21674, B2 => n9446, C1 => n21682, C2 => 
                           n19685, A => n17270, ZN => n17266);
   U15608 : OAI22_X1 port map( A1 => n16496, A2 => n21697, B1 => n15831, B2 => 
                           n21689, ZN => n17270);
   U15609 : AOI221_X1 port map( B1 => n21423, B2 => n8652, C1 => n21438, C2 => 
                           n19771, A => n17257, ZN => n17228);
   U15610 : OAI22_X1 port map( A1 => n16179, A2 => n21451, B1 => n16317, B2 => 
                           n21459, ZN => n17257);
   U15611 : AOI221_X1 port map( B1 => n21669, B2 => n9445, C1 => n21678, C2 => 
                           n19772, A => n17223, ZN => n17219);
   U15612 : OAI22_X1 port map( A1 => n16495, A2 => n21695, B1 => n15830, B2 => 
                           n21685, ZN => n17223);
   U15613 : AOI221_X1 port map( B1 => n21429, B2 => n8641, C1 => n21439, C2 => 
                           n19773, A => n17210, ZN => n17181);
   U15614 : OAI22_X1 port map( A1 => n16178, A2 => n21451, B1 => n16316, B2 => 
                           n21458, ZN => n17210);
   U15615 : AOI221_X1 port map( B1 => n21674, B2 => n9444, C1 => n21677, C2 => 
                           n19774, A => n17176, ZN => n17172);
   U15616 : OAI22_X1 port map( A1 => n16494, A2 => n21698, B1 => n15829, B2 => 
                           n21684, ZN => n17176);
   U15617 : AOI221_X1 port map( B1 => n21424, B2 => n8630, C1 => n21439, C2 => 
                           n19775, A => n17163, ZN => n17134);
   U15618 : OAI22_X1 port map( A1 => n16177, A2 => n21450, B1 => n16315, B2 => 
                           n21459, ZN => n17163);
   U15619 : AOI221_X1 port map( B1 => n21669, B2 => n9443, C1 => n21677, C2 => 
                           n19776, A => n17129, ZN => n17125);
   U15620 : OAI22_X1 port map( A1 => n16493, A2 => n21697, B1 => n15828, B2 => 
                           n21690, ZN => n17129);
   U15621 : AOI221_X1 port map( B1 => n21424, B2 => n8619, C1 => n21439, C2 => 
                           n19777, A => n17116, ZN => n17087);
   U15622 : OAI22_X1 port map( A1 => n16176, A2 => n21451, B1 => n16314, B2 => 
                           n21458, ZN => n17116);
   U15623 : AOI221_X1 port map( B1 => n21669, B2 => n9442, C1 => n21680, C2 => 
                           n19778, A => n17082, ZN => n17078);
   U15624 : OAI22_X1 port map( A1 => n16492, A2 => n21692, B1 => n15827, B2 => 
                           n21690, ZN => n17082);
   U15625 : AOI221_X1 port map( B1 => n21670, B2 => n9441, C1 => n21678, C2 => 
                           n19779, A => n17035, ZN => n17031);
   U15626 : OAI22_X1 port map( A1 => n16491, A2 => n21698, B1 => n15826, B2 => 
                           n21690, ZN => n17035);
   U15627 : AOI221_X1 port map( B1 => n21671, B2 => n9440, C1 => n21678, C2 => 
                           n19780, A => n16988, ZN => n16984);
   U15628 : OAI22_X1 port map( A1 => n16490, A2 => n21698, B1 => n15825, B2 => 
                           n21686, ZN => n16988);
   U15629 : NOR2_X1 port map( A1 => n16653, A2 => ADD_WR(3), ZN => n15366);
   U15630 : AOI221_X1 port map( B1 => n20800, B2 => n8906, C1 => n20841, C2 => 
                           n19781, A => n19613, ZN => n19590);
   U15631 : OAI22_X1 port map( A1 => n16755, A2 => n20849, B1 => n4289, B2 => 
                           n20852, ZN => n19613);
   U15632 : AOI221_X1 port map( B1 => n21205, B2 => n8570, C1 => n21210, C2 => 
                           n9018, A => n19587, ZN => n19582);
   U15633 : OAI22_X1 port map( A1 => n16063, A2 => n21199, B1 => n16097, B2 => 
                           n21187, ZN => n19587);
   U15634 : AOI221_X1 port map( B1 => n20800, B2 => n8895, C1 => n20839, C2 => 
                           n19782, A => n19576, ZN => n19553);
   U15635 : OAI22_X1 port map( A1 => n16754, A2 => n20843, B1 => n4291, B2 => 
                           n20853, ZN => n19576);
   U15636 : AOI221_X1 port map( B1 => n21208, B2 => n8568, C1 => n21209, C2 => 
                           n9016, A => n19550, ZN => n19545);
   U15637 : OAI22_X1 port map( A1 => n16062, A2 => n21195, B1 => n16096, B2 => 
                           n21191, ZN => n19550);
   U15638 : AOI221_X1 port map( B1 => n20803, B2 => n8884, C1 => n20839, C2 => 
                           n19783, A => n19539, ZN => n19516);
   U15639 : OAI22_X1 port map( A1 => n16753, A2 => n20844, B1 => n4293, B2 => 
                           n20856, ZN => n19539);
   U15640 : AOI221_X1 port map( B1 => n21207, B2 => n8566, C1 => n21209, C2 => 
                           n9014, A => n19513, ZN => n19508);
   U15641 : OAI22_X1 port map( A1 => n16061, A2 => n21194, B1 => n16095, B2 => 
                           n21188, ZN => n19513);
   U15642 : AOI221_X1 port map( B1 => n20801, B2 => n8873, C1 => n20840, C2 => 
                           n19784, A => n19502, ZN => n19479);
   U15643 : OAI22_X1 port map( A1 => n16752, A2 => n20844, B1 => n4295, B2 => 
                           n20853, ZN => n19502);
   U15644 : AOI221_X1 port map( B1 => n21203, B2 => n8564, C1 => n21211, C2 => 
                           n9012, A => n19476, ZN => n19471);
   U15645 : OAI22_X1 port map( A1 => n16060, A2 => n21198, B1 => n16094, B2 => 
                           n21192, ZN => n19476);
   U15646 : AOI221_X1 port map( B1 => n20801, B2 => n8862, C1 => n20840, C2 => 
                           n19785, A => n19465, ZN => n19442);
   U15647 : OAI22_X1 port map( A1 => n16751, A2 => n20846, B1 => n4297, B2 => 
                           n20854, ZN => n19465);
   U15648 : AOI221_X1 port map( B1 => n21203, B2 => n8562, C1 => n21210, C2 => 
                           n9010, A => n19439, ZN => n19434);
   U15649 : OAI22_X1 port map( A1 => n16059, A2 => n21195, B1 => n16093, B2 => 
                           n21186, ZN => n19439);
   U15650 : AOI221_X1 port map( B1 => n20802, B2 => n8851, C1 => n20841, C2 => 
                           n19786, A => n19428, ZN => n19405);
   U15651 : OAI22_X1 port map( A1 => n16750, A2 => n20845, B1 => n4299, B2 => 
                           n20854, ZN => n19428);
   U15652 : AOI221_X1 port map( B1 => n21203, B2 => n8560, C1 => n21210, C2 => 
                           n9008, A => n19402, ZN => n19397);
   U15653 : OAI22_X1 port map( A1 => n16058, A2 => n21196, B1 => n16092, B2 => 
                           n21187, ZN => n19402);
   U15654 : AOI221_X1 port map( B1 => n20802, B2 => n8840, C1 => n20839, C2 => 
                           n19787, A => n19391, ZN => n19368);
   U15655 : OAI22_X1 port map( A1 => n16749, A2 => n20845, B1 => n4301, B2 => 
                           n20856, ZN => n19391);
   U15656 : AOI221_X1 port map( B1 => n21204, B2 => n8558, C1 => n21209, C2 => 
                           n9006, A => n19365, ZN => n19360);
   U15657 : OAI22_X1 port map( A1 => n16057, A2 => n21196, B1 => n16091, B2 => 
                           n21187, ZN => n19365);
   U15658 : AOI221_X1 port map( B1 => n20802, B2 => n8829, C1 => n20841, C2 => 
                           n19788, A => n19354, ZN => n19331);
   U15659 : OAI22_X1 port map( A1 => n16748, A2 => n20845, B1 => n4303, B2 => 
                           n20853, ZN => n19354);
   U15660 : AOI221_X1 port map( B1 => n21204, B2 => n8556, C1 => n21211, C2 => 
                           n9004, A => n19328, ZN => n19323);
   U15661 : OAI22_X1 port map( A1 => n16056, A2 => n21197, B1 => n16090, B2 => 
                           n21188, ZN => n19328);
   U15662 : AOI221_X1 port map( B1 => n20803, B2 => n8818, C1 => n20840, C2 => 
                           n19789, A => n19317, ZN => n19294);
   U15663 : OAI22_X1 port map( A1 => n16747, A2 => n20844, B1 => n4305, B2 => 
                           n20857, ZN => n19317);
   U15664 : AOI221_X1 port map( B1 => n21205, B2 => n8554, C1 => n21211, C2 => 
                           n9002, A => n19291, ZN => n19286);
   U15665 : OAI22_X1 port map( A1 => n16055, A2 => n21196, B1 => n16089, B2 => 
                           n21186, ZN => n19291);
   U15666 : AOI221_X1 port map( B1 => n20803, B2 => n8807, C1 => n20841, C2 => 
                           n19790, A => n19280, ZN => n19257);
   U15667 : OAI22_X1 port map( A1 => n16746, A2 => n20846, B1 => n4307, B2 => 
                           n20855, ZN => n19280);
   U15668 : AOI221_X1 port map( B1 => n21204, B2 => n8552, C1 => n21210, C2 => 
                           n9000, A => n19254, ZN => n19249);
   U15669 : OAI22_X1 port map( A1 => n16054, A2 => n21195, B1 => n16088, B2 => 
                           n21188, ZN => n19254);
   U15670 : AOI221_X1 port map( B1 => n20804, B2 => n8796, C1 => n20839, C2 => 
                           n19791, A => n19243, ZN => n19220);
   U15671 : OAI22_X1 port map( A1 => n16745, A2 => n20847, B1 => n4309, B2 => 
                           n20856, ZN => n19243);
   U15672 : AOI221_X1 port map( B1 => n21206, B2 => n8550, C1 => n21209, C2 => 
                           n8998, A => n19217, ZN => n19212);
   U15673 : OAI22_X1 port map( A1 => n16053, A2 => n21198, B1 => n16087, B2 => 
                           n21189, ZN => n19217);
   U15674 : AOI221_X1 port map( B1 => n20804, B2 => n8785, C1 => n20839, C2 => 
                           n19792, A => n19206, ZN => n19183);
   U15675 : OAI22_X1 port map( A1 => n16744, A2 => n20844, B1 => n4311, B2 => 
                           n20853, ZN => n19206);
   U15676 : AOI221_X1 port map( B1 => n21206, B2 => n8548, C1 => n21209, C2 => 
                           n8996, A => n19180, ZN => n19175);
   U15677 : OAI22_X1 port map( A1 => n16052, A2 => n21195, B1 => n16086, B2 => 
                           n21186, ZN => n19180);
   U15678 : AOI221_X1 port map( B1 => n20801, B2 => n8774, C1 => n20840, C2 => 
                           n19793, A => n19169, ZN => n19146);
   U15679 : OAI22_X1 port map( A1 => n16743, A2 => n20845, B1 => n4313, B2 => 
                           n20854, ZN => n19169);
   U15680 : AOI221_X1 port map( B1 => n21207, B2 => n8546, C1 => n21211, C2 => 
                           n8994, A => n19143, ZN => n19138);
   U15681 : OAI22_X1 port map( A1 => n16051, A2 => n21197, B1 => n16085, B2 => 
                           n21187, ZN => n19143);
   U15682 : AOI221_X1 port map( B1 => n20803, B2 => n8763, C1 => n20840, C2 => 
                           n19794, A => n19132, ZN => n19109);
   U15683 : OAI22_X1 port map( A1 => n16742, A2 => n20845, B1 => n4315, B2 => 
                           n20854, ZN => n19132);
   U15684 : AOI221_X1 port map( B1 => n21206, B2 => n8544, C1 => n21210, C2 => 
                           n8992, A => n19106, ZN => n19101);
   U15685 : OAI22_X1 port map( A1 => n16050, A2 => n21196, B1 => n16084, B2 => 
                           n21188, ZN => n19106);
   U15686 : AOI221_X1 port map( B1 => n20804, B2 => n8752, C1 => n20841, C2 => 
                           n19795, A => n19095, ZN => n19072);
   U15687 : OAI22_X1 port map( A1 => n16741, A2 => n20848, B1 => n4317, B2 => 
                           n20852, ZN => n19095);
   U15688 : AOI221_X1 port map( B1 => n21206, B2 => n8542, C1 => n21210, C2 => 
                           n8990, A => n19069, ZN => n19064);
   U15689 : OAI22_X1 port map( A1 => n16049, A2 => n21197, B1 => n16083, B2 => 
                           n21188, ZN => n19069);
   U15690 : AOI221_X1 port map( B1 => n20802, B2 => n8741, C1 => n20839, C2 => 
                           n19796, A => n19058, ZN => n19035);
   U15691 : OAI22_X1 port map( A1 => n16740, A2 => n20845, B1 => n4319, B2 => 
                           n20852, ZN => n19058);
   U15692 : AOI221_X1 port map( B1 => n21207, B2 => n8540, C1 => n21209, C2 => 
                           n8988, A => n19032, ZN => n19027);
   U15693 : OAI22_X1 port map( A1 => n16048, A2 => n21197, B1 => n16082, B2 => 
                           n21192, ZN => n19032);
   U15694 : AOI221_X1 port map( B1 => n20803, B2 => n8730, C1 => n20841, C2 => 
                           n19797, A => n19021, ZN => n18998);
   U15695 : OAI22_X1 port map( A1 => n16739, A2 => n20843, B1 => n4321, B2 => 
                           n20854, ZN => n19021);
   U15696 : AOI221_X1 port map( B1 => n21207, B2 => n8538, C1 => n21211, C2 => 
                           n8986, A => n18995, ZN => n18990);
   U15697 : OAI22_X1 port map( A1 => n16047, A2 => n21194, B1 => n16081, B2 => 
                           n21187, ZN => n18995);
   U15698 : AOI221_X1 port map( B1 => n20805, B2 => n8719, C1 => n20840, C2 => 
                           n19798, A => n18984, ZN => n18961);
   U15699 : OAI22_X1 port map( A1 => n16738, A2 => n20846, B1 => n4323, B2 => 
                           n20855, ZN => n18984);
   U15700 : AOI221_X1 port map( B1 => n21205, B2 => n8536, C1 => n21211, C2 => 
                           n8984, A => n18958, ZN => n18953);
   U15701 : OAI22_X1 port map( A1 => n16046, A2 => n21198, B1 => n16080, B2 => 
                           n21189, ZN => n18958);
   U15702 : AOI221_X1 port map( B1 => n20805, B2 => n8708, C1 => n20841, C2 => 
                           n19799, A => n18947, ZN => n18924);
   U15703 : OAI22_X1 port map( A1 => n16737, A2 => n20847, B1 => n4325, B2 => 
                           n20855, ZN => n18947);
   U15704 : AOI221_X1 port map( B1 => n21207, B2 => n8534, C1 => n21210, C2 => 
                           n8982, A => n18921, ZN => n18916);
   U15705 : OAI22_X1 port map( A1 => n16045, A2 => n21199, B1 => n16079, B2 => 
                           n21190, ZN => n18921);
   U15706 : AOI221_X1 port map( B1 => n20805, B2 => n8697, C1 => n20839, C2 => 
                           n19800, A => n18910, ZN => n18887);
   U15707 : OAI22_X1 port map( A1 => n16736, A2 => n20846, B1 => n4327, B2 => 
                           n20856, ZN => n18910);
   U15708 : AOI221_X1 port map( B1 => n21208, B2 => n8532, C1 => n21209, C2 => 
                           n8980, A => n18884, ZN => n18879);
   U15709 : OAI22_X1 port map( A1 => n16044, A2 => n21194, B1 => n16078, B2 => 
                           n21186, ZN => n18884);
   U15710 : AOI221_X1 port map( B1 => n20805, B2 => n8686, C1 => n20839, C2 => 
                           n19686, A => n18873, ZN => n18850);
   U15711 : OAI22_X1 port map( A1 => n16735, A2 => n20847, B1 => n4329, B2 => 
                           n20858, ZN => n18873);
   U15712 : AOI221_X1 port map( B1 => n21208, B2 => n8530, C1 => n21209, C2 => 
                           n8978, A => n18847, ZN => n18842);
   U15713 : OAI22_X1 port map( A1 => n16043, A2 => n21199, B1 => n16077, B2 => 
                           n21189, ZN => n18847);
   U15714 : AOI221_X1 port map( B1 => n20800, B2 => n8675, C1 => n20840, C2 => 
                           n19801, A => n18836, ZN => n18813);
   U15715 : OAI22_X1 port map( A1 => n16734, A2 => n20848, B1 => n4331, B2 => 
                           n20856, ZN => n18836);
   U15716 : AOI221_X1 port map( B1 => n21208, B2 => n8528, C1 => n21211, C2 => 
                           n8976, A => n18810, ZN => n18805);
   U15717 : OAI22_X1 port map( A1 => n16042, A2 => n21198, B1 => n16076, B2 => 
                           n21190, ZN => n18810);
   U15718 : AOI221_X1 port map( B1 => n20800, B2 => n8664, C1 => n20840, C2 => 
                           n19802, A => n18799, ZN => n18776);
   U15719 : OAI22_X1 port map( A1 => n16733, A2 => n20848, B1 => n4333, B2 => 
                           n20857, ZN => n18799);
   U15720 : AOI221_X1 port map( B1 => n21208, B2 => n8526, C1 => n21210, C2 => 
                           n8974, A => n18773, ZN => n18768);
   U15721 : OAI22_X1 port map( A1 => n16041, A2 => n21199, B1 => n16075, B2 => 
                           n21190, ZN => n18773);
   U15722 : AOI221_X1 port map( B1 => n20800, B2 => n8653, C1 => n20841, C2 => 
                           n19803, A => n18762, ZN => n18739);
   U15723 : OAI22_X1 port map( A1 => n16732, A2 => n20849, B1 => n4335, B2 => 
                           n20857, ZN => n18762);
   U15724 : AOI221_X1 port map( B1 => n21205, B2 => n8524, C1 => n21210, C2 => 
                           n8972, A => n18736, ZN => n18731);
   U15725 : OAI22_X1 port map( A1 => n16040, A2 => n21200, B1 => n16074, B2 => 
                           n21192, ZN => n18736);
   U15726 : AOI221_X1 port map( B1 => n20801, B2 => n8642, C1 => n20839, C2 => 
                           n19804, A => n18725, ZN => n18702);
   U15727 : OAI22_X1 port map( A1 => n16731, A2 => n20849, B1 => n4337, B2 => 
                           n20858, ZN => n18725);
   U15728 : AOI221_X1 port map( B1 => n21208, B2 => n8522, C1 => n21209, C2 => 
                           n8970, A => n18699, ZN => n18694);
   U15729 : OAI22_X1 port map( A1 => n16039, A2 => n21200, B1 => n16073, B2 => 
                           n21191, ZN => n18699);
   U15730 : AOI221_X1 port map( B1 => n20801, B2 => n8631, C1 => n20841, C2 => 
                           n19805, A => n18688, ZN => n18665);
   U15731 : OAI22_X1 port map( A1 => n16730, A2 => n20848, B1 => n4339, B2 => 
                           n20857, ZN => n18688);
   U15732 : AOI221_X1 port map( B1 => n21205, B2 => n8520, C1 => n21211, C2 => 
                           n8968, A => n18662, ZN => n18657);
   U15733 : OAI22_X1 port map( A1 => n16038, A2 => n21199, B1 => n16072, B2 => 
                           n21192, ZN => n18662);
   U15734 : AOI221_X1 port map( B1 => n20805, B2 => n8620, C1 => n20840, C2 => 
                           n19806, A => n18651, ZN => n18628);
   U15735 : OAI22_X1 port map( A1 => n16729, A2 => n20849, B1 => n4341, B2 => 
                           n20858, ZN => n18651);
   U15736 : AOI221_X1 port map( B1 => n21203, B2 => n8518, C1 => n21211, C2 => 
                           n8966, A => n18625, ZN => n18620);
   U15737 : OAI22_X1 port map( A1 => n16037, A2 => n21200, B1 => n16071, B2 => 
                           n21191, ZN => n18625);
   U15738 : AOI221_X1 port map( B1 => n20802, B2 => n8609, C1 => n20841, C2 => 
                           n19807, A => n18614, ZN => n18591);
   U15739 : OAI22_X1 port map( A1 => n16728, A2 => n20848, B1 => n4343, B2 => 
                           n20855, ZN => n18614);
   U15740 : AOI221_X1 port map( B1 => n21204, B2 => n8516, C1 => n21210, C2 => 
                           n8964, A => n18588, ZN => n18583);
   U15741 : OAI22_X1 port map( A1 => n16036, A2 => n21200, B1 => n16070, B2 => 
                           n21192, ZN => n18588);
   U15742 : AOI221_X1 port map( B1 => n20802, B2 => n8598, C1 => n20839, C2 => 
                           n19808, A => n18577, ZN => n18554);
   U15743 : OAI22_X1 port map( A1 => n16727, A2 => n20847, B1 => n4345, B2 => 
                           n20852, ZN => n18577);
   U15744 : AOI221_X1 port map( B1 => n21203, B2 => n8514, C1 => n21209, C2 => 
                           n8962, A => n18551, ZN => n18546);
   U15745 : OAI22_X1 port map( A1 => n16035, A2 => n21195, B1 => n16069, B2 => 
                           n21191, ZN => n18551);
   U15746 : AOI221_X1 port map( B1 => n20804, B2 => n8587, C1 => n20839, C2 => 
                           n19809, A => n18540, ZN => n18517);
   U15747 : OAI22_X1 port map( A1 => n16726, A2 => n20843, B1 => n4347, B2 => 
                           n20852, ZN => n18540);
   U15748 : AOI221_X1 port map( B1 => n21204, B2 => n8512, C1 => n21209, C2 => 
                           n8960, A => n18514, ZN => n18509);
   U15749 : OAI22_X1 port map( A1 => n16034, A2 => n21200, B1 => n16068, B2 => 
                           n21190, ZN => n18514);
   U15750 : AOI221_X1 port map( B1 => n20804, B2 => n8576, C1 => n20840, C2 => 
                           n19810, A => n18497, ZN => n18447);
   U15751 : OAI22_X1 port map( A1 => n16725, A2 => n20843, B1 => n4349, B2 => 
                           n20858, ZN => n18497);
   U15752 : AOI221_X1 port map( B1 => n21205, B2 => n8510, C1 => n21211, C2 => 
                           n8958, A => n18438, ZN => n18422);
   U15753 : OAI22_X1 port map( A1 => n16033, A2 => n21194, B1 => n16067, B2 => 
                           n21189, ZN => n18438);
   U15754 : AOI221_X1 port map( B1 => n21357, B2 => n8906, C1 => n21398, C2 => 
                           n19781, A => n18340, ZN => n18308);
   U15755 : OAI22_X1 port map( A1 => n16755, A2 => n21406, B1 => n4289, B2 => 
                           n21409, ZN => n18340);
   U15756 : AOI221_X1 port map( B1 => n21762, B2 => n8570, C1 => n21767, C2 => 
                           n9018, A => n18305, ZN => n18299);
   U15757 : OAI22_X1 port map( A1 => n16063, A2 => n21756, B1 => n16097, B2 => 
                           n21744, ZN => n18305);
   U15758 : AOI221_X1 port map( B1 => n21357, B2 => n8895, C1 => n21396, C2 => 
                           n19782, A => n18293, ZN => n18261);
   U15759 : OAI22_X1 port map( A1 => n16754, A2 => n21400, B1 => n4291, B2 => 
                           n21410, ZN => n18293);
   U15760 : AOI221_X1 port map( B1 => n21765, B2 => n8568, C1 => n21766, C2 => 
                           n9016, A => n18258, ZN => n18252);
   U15761 : OAI22_X1 port map( A1 => n16062, A2 => n21752, B1 => n16096, B2 => 
                           n21748, ZN => n18258);
   U15762 : AOI221_X1 port map( B1 => n21360, B2 => n8884, C1 => n21396, C2 => 
                           n19783, A => n18246, ZN => n18214);
   U15763 : OAI22_X1 port map( A1 => n16753, A2 => n21401, B1 => n4293, B2 => 
                           n21413, ZN => n18246);
   U15764 : AOI221_X1 port map( B1 => n21764, B2 => n8566, C1 => n21766, C2 => 
                           n9014, A => n18211, ZN => n18205);
   U15765 : OAI22_X1 port map( A1 => n16061, A2 => n21751, B1 => n16095, B2 => 
                           n21745, ZN => n18211);
   U15766 : AOI221_X1 port map( B1 => n21358, B2 => n8873, C1 => n21397, C2 => 
                           n19784, A => n18199, ZN => n18167);
   U15767 : OAI22_X1 port map( A1 => n16752, A2 => n21401, B1 => n4295, B2 => 
                           n21410, ZN => n18199);
   U15768 : AOI221_X1 port map( B1 => n21760, B2 => n8564, C1 => n21768, C2 => 
                           n9012, A => n18164, ZN => n18158);
   U15769 : OAI22_X1 port map( A1 => n16060, A2 => n21755, B1 => n16094, B2 => 
                           n21749, ZN => n18164);
   U15770 : AOI221_X1 port map( B1 => n21358, B2 => n8862, C1 => n21397, C2 => 
                           n19785, A => n18152, ZN => n18120);
   U15771 : OAI22_X1 port map( A1 => n16751, A2 => n21403, B1 => n4297, B2 => 
                           n21411, ZN => n18152);
   U15772 : AOI221_X1 port map( B1 => n21760, B2 => n8562, C1 => n21767, C2 => 
                           n9010, A => n18117, ZN => n18111);
   U15773 : OAI22_X1 port map( A1 => n16059, A2 => n21752, B1 => n16093, B2 => 
                           n21743, ZN => n18117);
   U15774 : AOI221_X1 port map( B1 => n21359, B2 => n8851, C1 => n21398, C2 => 
                           n19786, A => n18105, ZN => n18073);
   U15775 : OAI22_X1 port map( A1 => n16750, A2 => n21402, B1 => n4299, B2 => 
                           n21411, ZN => n18105);
   U15776 : AOI221_X1 port map( B1 => n21760, B2 => n8560, C1 => n21767, C2 => 
                           n9008, A => n18070, ZN => n18064);
   U15777 : OAI22_X1 port map( A1 => n16058, A2 => n21753, B1 => n16092, B2 => 
                           n21744, ZN => n18070);
   U15778 : AOI221_X1 port map( B1 => n21359, B2 => n8840, C1 => n21396, C2 => 
                           n19787, A => n18058, ZN => n18026);
   U15779 : OAI22_X1 port map( A1 => n16749, A2 => n21402, B1 => n4301, B2 => 
                           n21413, ZN => n18058);
   U15780 : AOI221_X1 port map( B1 => n21761, B2 => n8558, C1 => n21766, C2 => 
                           n9006, A => n18023, ZN => n18017);
   U15781 : OAI22_X1 port map( A1 => n16057, A2 => n21753, B1 => n16091, B2 => 
                           n21744, ZN => n18023);
   U15782 : AOI221_X1 port map( B1 => n21359, B2 => n8829, C1 => n21398, C2 => 
                           n19788, A => n18011, ZN => n17979);
   U15783 : OAI22_X1 port map( A1 => n16748, A2 => n21402, B1 => n4303, B2 => 
                           n21410, ZN => n18011);
   U15784 : AOI221_X1 port map( B1 => n21761, B2 => n8556, C1 => n21768, C2 => 
                           n9004, A => n17976, ZN => n17970);
   U15785 : OAI22_X1 port map( A1 => n16056, A2 => n21754, B1 => n16090, B2 => 
                           n21745, ZN => n17976);
   U15786 : AOI221_X1 port map( B1 => n21360, B2 => n8818, C1 => n21397, C2 => 
                           n19789, A => n17964, ZN => n17932);
   U15787 : OAI22_X1 port map( A1 => n16747, A2 => n21401, B1 => n4305, B2 => 
                           n21414, ZN => n17964);
   U15788 : AOI221_X1 port map( B1 => n21762, B2 => n8554, C1 => n21768, C2 => 
                           n9002, A => n17929, ZN => n17923);
   U15789 : OAI22_X1 port map( A1 => n16055, A2 => n21753, B1 => n16089, B2 => 
                           n21743, ZN => n17929);
   U15790 : AOI221_X1 port map( B1 => n21360, B2 => n8807, C1 => n21398, C2 => 
                           n19790, A => n17917, ZN => n17885);
   U15791 : OAI22_X1 port map( A1 => n16746, A2 => n21403, B1 => n4307, B2 => 
                           n21412, ZN => n17917);
   U15792 : AOI221_X1 port map( B1 => n21761, B2 => n8552, C1 => n21767, C2 => 
                           n9000, A => n17882, ZN => n17876);
   U15793 : OAI22_X1 port map( A1 => n16054, A2 => n21752, B1 => n16088, B2 => 
                           n21745, ZN => n17882);
   U15794 : AOI221_X1 port map( B1 => n21361, B2 => n8796, C1 => n21396, C2 => 
                           n19791, A => n17870, ZN => n17838);
   U15795 : OAI22_X1 port map( A1 => n16745, A2 => n21404, B1 => n4309, B2 => 
                           n21413, ZN => n17870);
   U15796 : AOI221_X1 port map( B1 => n21763, B2 => n8550, C1 => n21766, C2 => 
                           n8998, A => n17835, ZN => n17829);
   U15797 : OAI22_X1 port map( A1 => n16053, A2 => n21755, B1 => n16087, B2 => 
                           n21746, ZN => n17835);
   U15798 : AOI221_X1 port map( B1 => n21361, B2 => n8785, C1 => n21396, C2 => 
                           n19792, A => n17823, ZN => n17791);
   U15799 : OAI22_X1 port map( A1 => n16744, A2 => n21401, B1 => n4311, B2 => 
                           n21410, ZN => n17823);
   U15800 : AOI221_X1 port map( B1 => n21763, B2 => n8548, C1 => n21766, C2 => 
                           n8996, A => n17788, ZN => n17782);
   U15801 : OAI22_X1 port map( A1 => n16052, A2 => n21752, B1 => n16086, B2 => 
                           n21743, ZN => n17788);
   U15802 : AOI221_X1 port map( B1 => n21358, B2 => n8774, C1 => n21397, C2 => 
                           n19793, A => n17776, ZN => n17744);
   U15803 : OAI22_X1 port map( A1 => n16743, A2 => n21402, B1 => n4313, B2 => 
                           n21411, ZN => n17776);
   U15804 : AOI221_X1 port map( B1 => n21764, B2 => n8546, C1 => n21768, C2 => 
                           n8994, A => n17741, ZN => n17735);
   U15805 : OAI22_X1 port map( A1 => n16051, A2 => n21754, B1 => n16085, B2 => 
                           n21744, ZN => n17741);
   U15806 : AOI221_X1 port map( B1 => n21360, B2 => n8763, C1 => n21397, C2 => 
                           n19794, A => n17729, ZN => n17697);
   U15807 : OAI22_X1 port map( A1 => n16742, A2 => n21402, B1 => n4315, B2 => 
                           n21411, ZN => n17729);
   U15808 : AOI221_X1 port map( B1 => n21763, B2 => n8544, C1 => n21767, C2 => 
                           n8992, A => n17694, ZN => n17688);
   U15809 : OAI22_X1 port map( A1 => n16050, A2 => n21753, B1 => n16084, B2 => 
                           n21745, ZN => n17694);
   U15810 : AOI221_X1 port map( B1 => n21361, B2 => n8752, C1 => n21398, C2 => 
                           n19795, A => n17682, ZN => n17650);
   U15811 : OAI22_X1 port map( A1 => n16741, A2 => n21405, B1 => n4317, B2 => 
                           n21409, ZN => n17682);
   U15812 : AOI221_X1 port map( B1 => n21763, B2 => n8542, C1 => n21767, C2 => 
                           n8990, A => n17647, ZN => n17641);
   U15813 : OAI22_X1 port map( A1 => n16049, A2 => n21754, B1 => n16083, B2 => 
                           n21745, ZN => n17647);
   U15814 : AOI221_X1 port map( B1 => n21359, B2 => n8741, C1 => n21396, C2 => 
                           n19796, A => n17635, ZN => n17603);
   U15815 : OAI22_X1 port map( A1 => n16740, A2 => n21402, B1 => n4319, B2 => 
                           n21409, ZN => n17635);
   U15816 : AOI221_X1 port map( B1 => n21764, B2 => n8540, C1 => n21766, C2 => 
                           n8988, A => n17600, ZN => n17594);
   U15817 : OAI22_X1 port map( A1 => n16048, A2 => n21754, B1 => n16082, B2 => 
                           n21749, ZN => n17600);
   U15818 : AOI221_X1 port map( B1 => n21360, B2 => n8730, C1 => n21398, C2 => 
                           n19797, A => n17588, ZN => n17556);
   U15819 : OAI22_X1 port map( A1 => n16739, A2 => n21400, B1 => n4321, B2 => 
                           n21411, ZN => n17588);
   U15820 : AOI221_X1 port map( B1 => n21764, B2 => n8538, C1 => n21768, C2 => 
                           n8986, A => n17553, ZN => n17547);
   U15821 : OAI22_X1 port map( A1 => n16047, A2 => n21751, B1 => n16081, B2 => 
                           n21744, ZN => n17553);
   U15822 : AOI221_X1 port map( B1 => n21362, B2 => n8719, C1 => n21397, C2 => 
                           n19798, A => n17541, ZN => n17509);
   U15823 : OAI22_X1 port map( A1 => n16738, A2 => n21403, B1 => n4323, B2 => 
                           n21412, ZN => n17541);
   U15824 : AOI221_X1 port map( B1 => n21762, B2 => n8536, C1 => n21768, C2 => 
                           n8984, A => n17506, ZN => n17500);
   U15825 : OAI22_X1 port map( A1 => n16046, A2 => n21755, B1 => n16080, B2 => 
                           n21746, ZN => n17506);
   U15826 : AOI221_X1 port map( B1 => n21362, B2 => n8708, C1 => n21398, C2 => 
                           n19799, A => n17494, ZN => n17462);
   U15827 : OAI22_X1 port map( A1 => n16737, A2 => n21404, B1 => n4325, B2 => 
                           n21412, ZN => n17494);
   U15828 : AOI221_X1 port map( B1 => n21764, B2 => n8534, C1 => n21767, C2 => 
                           n8982, A => n17459, ZN => n17453);
   U15829 : OAI22_X1 port map( A1 => n16045, A2 => n21756, B1 => n16079, B2 => 
                           n21747, ZN => n17459);
   U15830 : AOI221_X1 port map( B1 => n21362, B2 => n8697, C1 => n21396, C2 => 
                           n19800, A => n17447, ZN => n17415);
   U15831 : OAI22_X1 port map( A1 => n16736, A2 => n21403, B1 => n4327, B2 => 
                           n21413, ZN => n17447);
   U15832 : AOI221_X1 port map( B1 => n21765, B2 => n8532, C1 => n21766, C2 => 
                           n8980, A => n17412, ZN => n17406);
   U15833 : OAI22_X1 port map( A1 => n16044, A2 => n21751, B1 => n16078, B2 => 
                           n21743, ZN => n17412);
   U15834 : AOI221_X1 port map( B1 => n21362, B2 => n8686, C1 => n21396, C2 => 
                           n19686, A => n17400, ZN => n17368);
   U15835 : OAI22_X1 port map( A1 => n16735, A2 => n21404, B1 => n4329, B2 => 
                           n21415, ZN => n17400);
   U15836 : AOI221_X1 port map( B1 => n21765, B2 => n8530, C1 => n21766, C2 => 
                           n8978, A => n17365, ZN => n17359);
   U15837 : OAI22_X1 port map( A1 => n16043, A2 => n21756, B1 => n16077, B2 => 
                           n21746, ZN => n17365);
   U15838 : AOI221_X1 port map( B1 => n21357, B2 => n8675, C1 => n21397, C2 => 
                           n19801, A => n17353, ZN => n17321);
   U15839 : OAI22_X1 port map( A1 => n16734, A2 => n21405, B1 => n4331, B2 => 
                           n21413, ZN => n17353);
   U15840 : AOI221_X1 port map( B1 => n21765, B2 => n8528, C1 => n21768, C2 => 
                           n8976, A => n17318, ZN => n17312);
   U15841 : OAI22_X1 port map( A1 => n16042, A2 => n21755, B1 => n16076, B2 => 
                           n21747, ZN => n17318);
   U15842 : AOI221_X1 port map( B1 => n21357, B2 => n8664, C1 => n21397, C2 => 
                           n19802, A => n17306, ZN => n17274);
   U15843 : OAI22_X1 port map( A1 => n16733, A2 => n21405, B1 => n4333, B2 => 
                           n21414, ZN => n17306);
   U15844 : AOI221_X1 port map( B1 => n21765, B2 => n8526, C1 => n21767, C2 => 
                           n8974, A => n17271, ZN => n17265);
   U15845 : OAI22_X1 port map( A1 => n16041, A2 => n21756, B1 => n16075, B2 => 
                           n21747, ZN => n17271);
   U15846 : AOI221_X1 port map( B1 => n21357, B2 => n8653, C1 => n21398, C2 => 
                           n19803, A => n17259, ZN => n17227);
   U15847 : OAI22_X1 port map( A1 => n16732, A2 => n21406, B1 => n4335, B2 => 
                           n21414, ZN => n17259);
   U15848 : AOI221_X1 port map( B1 => n21762, B2 => n8524, C1 => n21767, C2 => 
                           n8972, A => n17224, ZN => n17218);
   U15849 : OAI22_X1 port map( A1 => n16040, A2 => n21757, B1 => n16074, B2 => 
                           n21749, ZN => n17224);
   U15850 : AOI221_X1 port map( B1 => n21358, B2 => n8642, C1 => n21396, C2 => 
                           n19804, A => n17212, ZN => n17180);
   U15851 : OAI22_X1 port map( A1 => n16731, A2 => n21406, B1 => n4337, B2 => 
                           n21415, ZN => n17212);
   U15852 : AOI221_X1 port map( B1 => n21765, B2 => n8522, C1 => n21766, C2 => 
                           n8970, A => n17177, ZN => n17171);
   U15853 : OAI22_X1 port map( A1 => n16039, A2 => n21757, B1 => n16073, B2 => 
                           n21748, ZN => n17177);
   U15854 : AOI221_X1 port map( B1 => n21358, B2 => n8631, C1 => n21398, C2 => 
                           n19805, A => n17165, ZN => n17133);
   U15855 : OAI22_X1 port map( A1 => n16730, A2 => n21405, B1 => n4339, B2 => 
                           n21414, ZN => n17165);
   U15856 : AOI221_X1 port map( B1 => n21762, B2 => n8520, C1 => n21768, C2 => 
                           n8968, A => n17130, ZN => n17124);
   U15857 : OAI22_X1 port map( A1 => n16038, A2 => n21756, B1 => n16072, B2 => 
                           n21749, ZN => n17130);
   U15858 : AOI221_X1 port map( B1 => n21362, B2 => n8620, C1 => n21397, C2 => 
                           n19806, A => n17118, ZN => n17086);
   U15859 : OAI22_X1 port map( A1 => n16729, A2 => n21406, B1 => n4341, B2 => 
                           n21415, ZN => n17118);
   U15860 : AOI221_X1 port map( B1 => n21760, B2 => n8518, C1 => n21768, C2 => 
                           n8966, A => n17083, ZN => n17077);
   U15861 : OAI22_X1 port map( A1 => n16037, A2 => n21757, B1 => n16071, B2 => 
                           n21748, ZN => n17083);
   U15862 : AOI221_X1 port map( B1 => n21359, B2 => n8609, C1 => n21398, C2 => 
                           n19807, A => n17071, ZN => n17039);
   U15863 : OAI22_X1 port map( A1 => n16728, A2 => n21405, B1 => n4343, B2 => 
                           n21412, ZN => n17071);
   U15864 : AOI221_X1 port map( B1 => n21761, B2 => n8516, C1 => n21767, C2 => 
                           n8964, A => n17036, ZN => n17030);
   U15865 : OAI22_X1 port map( A1 => n16036, A2 => n21757, B1 => n16070, B2 => 
                           n21749, ZN => n17036);
   U15866 : AOI221_X1 port map( B1 => n21359, B2 => n8598, C1 => n21396, C2 => 
                           n19808, A => n17024, ZN => n16992);
   U15867 : OAI22_X1 port map( A1 => n16727, A2 => n21404, B1 => n4345, B2 => 
                           n21409, ZN => n17024);
   U15868 : AOI221_X1 port map( B1 => n21760, B2 => n8514, C1 => n21766, C2 => 
                           n8962, A => n16989, ZN => n16983);
   U15869 : OAI22_X1 port map( A1 => n16035, A2 => n21752, B1 => n16069, B2 => 
                           n21748, ZN => n16989);
   U15870 : AOI221_X1 port map( B1 => n21361, B2 => n8587, C1 => n21396, C2 => 
                           n19809, A => n16977, ZN => n16945);
   U15871 : OAI22_X1 port map( A1 => n16726, A2 => n21400, B1 => n4347, B2 => 
                           n21409, ZN => n16977);
   U15872 : AOI221_X1 port map( B1 => n21761, B2 => n8512, C1 => n21766, C2 => 
                           n8960, A => n16942, ZN => n16936);
   U15873 : OAI22_X1 port map( A1 => n16034, A2 => n21757, B1 => n16068, B2 => 
                           n21747, ZN => n16942);
   U15874 : AOI221_X1 port map( B1 => n21361, B2 => n8576, C1 => n21397, C2 => 
                           n19810, A => n16924, ZN => n16865);
   U15875 : OAI22_X1 port map( A1 => n16725, A2 => n21400, B1 => n4349, B2 => 
                           n21415, ZN => n16924);
   U15876 : AOI221_X1 port map( B1 => n21762, B2 => n8510, C1 => n21768, C2 => 
                           n8958, A => n16856, ZN => n16839);
   U15877 : OAI22_X1 port map( A1 => n16033, A2 => n21751, B1 => n16067, B2 => 
                           n21746, ZN => n16856);
   U15878 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(5), A3 => n19665,
                           ZN => n19663);
   U15879 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(5), A3 => n18399,
                           ZN => n18396);
   U15880 : NOR3_X1 port map( A1 => ADD_RD1(4), A2 => ADD_RD1(5), A3 => 
                           ADD_RD1(3), ZN => n19660);
   U15881 : NOR3_X1 port map( A1 => ADD_RD2(4), A2 => ADD_RD2(5), A3 => 
                           ADD_RD2(3), ZN => n18393);
   U15882 : AOI221_X1 port map( B1 => n21213, B2 => n8571, C1 => n21226, C2 => 
                           n9019, A => n19588, ZN => n19581);
   U15883 : OAI22_X1 port map( A1 => n15502, A2 => n21237, B1 => n15468, B2 => 
                           n21232, ZN => n19588);
   U15884 : AOI221_X1 port map( B1 => n21214, B2 => n8569, C1 => n21223, C2 => 
                           n9017, A => n19551, ZN => n19544);
   U15885 : OAI22_X1 port map( A1 => n15501, A2 => n21242, B1 => n15467, B2 => 
                           n21229, ZN => n19551);
   U15886 : AOI221_X1 port map( B1 => n21214, B2 => n8567, C1 => n21221, C2 => 
                           n9015, A => n19514, ZN => n19507);
   U15887 : OAI22_X1 port map( A1 => n15500, A2 => n21237, B1 => n15466, B2 => 
                           n21229, ZN => n19514);
   U15888 : AOI221_X1 port map( B1 => n21215, B2 => n8563, C1 => n21222, C2 => 
                           n9011, A => n19440, ZN => n19433);
   U15889 : OAI22_X1 port map( A1 => n15498, A2 => n21238, B1 => n15464, B2 => 
                           n21229, ZN => n19440);
   U15890 : AOI221_X1 port map( B1 => n21213, B2 => n8561, C1 => n21222, C2 => 
                           n9009, A => n19403, ZN => n19396);
   U15891 : OAI22_X1 port map( A1 => n15497, A2 => n21240, B1 => n15463, B2 => 
                           n21230, ZN => n19403);
   U15892 : AOI221_X1 port map( B1 => n21215, B2 => n8559, C1 => n21223, C2 => 
                           n9007, A => n19366, ZN => n19359);
   U15893 : OAI22_X1 port map( A1 => n15496, A2 => n21239, B1 => n15462, B2 => 
                           n21231, ZN => n19366);
   U15894 : AOI221_X1 port map( B1 => n21216, B2 => n8557, C1 => n21224, C2 => 
                           n9005, A => n19329, ZN => n19322);
   U15895 : OAI22_X1 port map( A1 => n15495, A2 => n21240, B1 => n15461, B2 => 
                           n21231, ZN => n19329);
   U15896 : AOI221_X1 port map( B1 => n21216, B2 => n8555, C1 => n21224, C2 => 
                           n9003, A => n19292, ZN => n19285);
   U15897 : OAI22_X1 port map( A1 => n15494, A2 => n21240, B1 => n15460, B2 => 
                           n21231, ZN => n19292);
   U15898 : AOI221_X1 port map( B1 => n21217, B2 => n8553, C1 => n21225, C2 => 
                           n9001, A => n19255, ZN => n19248);
   U15899 : OAI22_X1 port map( A1 => n15493, A2 => n21237, B1 => n15459, B2 => 
                           n21235, ZN => n19255);
   U15900 : AOI221_X1 port map( B1 => n21217, B2 => n8551, C1 => n21226, C2 => 
                           n8999, A => n19218, ZN => n19211);
   U15901 : OAI22_X1 port map( A1 => n15492, A2 => n21241, B1 => n15458, B2 => 
                           n21232, ZN => n19218);
   U15902 : AOI221_X1 port map( B1 => n21217, B2 => n8549, C1 => n21226, C2 => 
                           n8997, A => n19181, ZN => n19174);
   U15903 : OAI22_X1 port map( A1 => n15491, A2 => n21238, B1 => n15457, B2 => 
                           n21229, ZN => n19181);
   U15904 : AOI221_X1 port map( B1 => n21218, B2 => n8547, C1 => n21227, C2 => 
                           n8995, A => n19144, ZN => n19137);
   U15905 : OAI22_X1 port map( A1 => n15490, A2 => n21239, B1 => n15456, B2 => 
                           n21230, ZN => n19144);
   U15906 : AOI221_X1 port map( B1 => n21217, B2 => n8545, C1 => n21222, C2 => 
                           n8993, A => n19107, ZN => n19100);
   U15907 : OAI22_X1 port map( A1 => n15489, A2 => n21239, B1 => n15455, B2 => 
                           n21231, ZN => n19107);
   U15908 : AOI221_X1 port map( B1 => n21217, B2 => n8543, C1 => n21224, C2 => 
                           n8991, A => n19070, ZN => n19063);
   U15909 : OAI22_X1 port map( A1 => n15488, A2 => n21240, B1 => n15454, B2 => 
                           n21230, ZN => n19070);
   U15910 : AOI221_X1 port map( B1 => n21218, B2 => n8541, C1 => n21225, C2 => 
                           n8989, A => n19033, ZN => n19026);
   U15911 : OAI22_X1 port map( A1 => n15487, A2 => n21239, B1 => n15453, B2 => 
                           n21233, ZN => n19033);
   U15912 : AOI221_X1 port map( B1 => n21218, B2 => n8539, C1 => n21226, C2 => 
                           n8987, A => n18996, ZN => n18989);
   U15913 : OAI22_X1 port map( A1 => n15486, A2 => n21238, B1 => n15452, B2 => 
                           n21234, ZN => n18996);
   U15914 : AOI221_X1 port map( B1 => n21216, B2 => n8537, C1 => n21226, C2 => 
                           n8985, A => n18959, ZN => n18952);
   U15915 : OAI22_X1 port map( A1 => n15485, A2 => n21241, B1 => n15451, B2 => 
                           n21232, ZN => n18959);
   U15916 : AOI221_X1 port map( B1 => n21218, B2 => n8535, C1 => n21227, C2 => 
                           n8983, A => n18922, ZN => n18915);
   U15917 : OAI22_X1 port map( A1 => n15484, A2 => n21242, B1 => n15450, B2 => 
                           n21233, ZN => n18922);
   U15918 : AOI221_X1 port map( B1 => n21219, B2 => n8533, C1 => n21227, C2 => 
                           n8981, A => n18885, ZN => n18878);
   U15919 : OAI22_X1 port map( A1 => n15483, A2 => n21237, B1 => n15449, B2 => 
                           n21229, ZN => n18885);
   U15920 : AOI221_X1 port map( B1 => n21219, B2 => n8531, C1 => n21227, C2 => 
                           n8979, A => n18848, ZN => n18841);
   U15921 : OAI22_X1 port map( A1 => n15482, A2 => n21242, B1 => n15448, B2 => 
                           n21232, ZN => n18848);
   U15922 : AOI221_X1 port map( B1 => n21215, B2 => n8513, C1 => n21223, C2 => 
                           n8961, A => n18515, ZN => n18508);
   U15923 : OAI22_X1 port map( A1 => n15473, A2 => n21238, B1 => n15439, B2 => 
                           n21233, ZN => n18515);
   U15924 : AOI221_X1 port map( B1 => n21215, B2 => n8511, C1 => n21224, C2 => 
                           n8959, A => n18443, ZN => n18421);
   U15925 : OAI22_X1 port map( A1 => n15472, A2 => n21241, B1 => n15438, B2 => 
                           n21230, ZN => n18443);
   U15926 : AOI221_X1 port map( B1 => n21770, B2 => n8571, C1 => n21783, C2 => 
                           n9019, A => n18306, ZN => n18298);
   U15927 : OAI22_X1 port map( A1 => n15502, A2 => n21794, B1 => n15468, B2 => 
                           n21789, ZN => n18306);
   U15928 : AOI221_X1 port map( B1 => n21771, B2 => n8569, C1 => n21780, C2 => 
                           n9017, A => n18259, ZN => n18251);
   U15929 : OAI22_X1 port map( A1 => n15501, A2 => n21799, B1 => n15467, B2 => 
                           n21786, ZN => n18259);
   U15930 : AOI221_X1 port map( B1 => n21771, B2 => n8567, C1 => n21778, C2 => 
                           n9015, A => n18212, ZN => n18204);
   U15931 : OAI22_X1 port map( A1 => n15500, A2 => n21794, B1 => n15466, B2 => 
                           n21786, ZN => n18212);
   U15932 : AOI221_X1 port map( B1 => n21772, B2 => n8563, C1 => n21779, C2 => 
                           n9011, A => n18118, ZN => n18110);
   U15933 : OAI22_X1 port map( A1 => n15498, A2 => n21795, B1 => n15464, B2 => 
                           n21786, ZN => n18118);
   U15934 : AOI221_X1 port map( B1 => n21770, B2 => n8561, C1 => n21779, C2 => 
                           n9009, A => n18071, ZN => n18063);
   U15935 : OAI22_X1 port map( A1 => n15497, A2 => n21797, B1 => n15463, B2 => 
                           n21787, ZN => n18071);
   U15936 : AOI221_X1 port map( B1 => n21772, B2 => n8559, C1 => n21780, C2 => 
                           n9007, A => n18024, ZN => n18016);
   U15937 : OAI22_X1 port map( A1 => n15496, A2 => n21796, B1 => n15462, B2 => 
                           n21788, ZN => n18024);
   U15938 : AOI221_X1 port map( B1 => n21773, B2 => n8557, C1 => n21781, C2 => 
                           n9005, A => n17977, ZN => n17969);
   U15939 : OAI22_X1 port map( A1 => n15495, A2 => n21797, B1 => n15461, B2 => 
                           n21788, ZN => n17977);
   U15940 : AOI221_X1 port map( B1 => n21773, B2 => n8555, C1 => n21781, C2 => 
                           n9003, A => n17930, ZN => n17922);
   U15941 : OAI22_X1 port map( A1 => n15494, A2 => n21797, B1 => n15460, B2 => 
                           n21788, ZN => n17930);
   U15942 : AOI221_X1 port map( B1 => n21774, B2 => n8553, C1 => n21782, C2 => 
                           n9001, A => n17883, ZN => n17875);
   U15943 : OAI22_X1 port map( A1 => n15493, A2 => n21794, B1 => n15459, B2 => 
                           n21792, ZN => n17883);
   U15944 : AOI221_X1 port map( B1 => n21774, B2 => n8551, C1 => n21783, C2 => 
                           n8999, A => n17836, ZN => n17828);
   U15945 : OAI22_X1 port map( A1 => n15492, A2 => n21798, B1 => n15458, B2 => 
                           n21789, ZN => n17836);
   U15946 : AOI221_X1 port map( B1 => n21774, B2 => n8549, C1 => n21783, C2 => 
                           n8997, A => n17789, ZN => n17781);
   U15947 : OAI22_X1 port map( A1 => n15491, A2 => n21795, B1 => n15457, B2 => 
                           n21786, ZN => n17789);
   U15948 : AOI221_X1 port map( B1 => n21775, B2 => n8547, C1 => n21784, C2 => 
                           n8995, A => n17742, ZN => n17734);
   U15949 : OAI22_X1 port map( A1 => n15490, A2 => n21796, B1 => n15456, B2 => 
                           n21787, ZN => n17742);
   U15950 : AOI221_X1 port map( B1 => n21774, B2 => n8545, C1 => n21779, C2 => 
                           n8993, A => n17695, ZN => n17687);
   U15951 : OAI22_X1 port map( A1 => n15489, A2 => n21796, B1 => n15455, B2 => 
                           n21788, ZN => n17695);
   U15952 : AOI221_X1 port map( B1 => n21774, B2 => n8543, C1 => n21781, C2 => 
                           n8991, A => n17648, ZN => n17640);
   U15953 : OAI22_X1 port map( A1 => n15488, A2 => n21797, B1 => n15454, B2 => 
                           n21787, ZN => n17648);
   U15954 : AOI221_X1 port map( B1 => n21775, B2 => n8541, C1 => n21782, C2 => 
                           n8989, A => n17601, ZN => n17593);
   U15955 : OAI22_X1 port map( A1 => n15487, A2 => n21796, B1 => n15453, B2 => 
                           n21790, ZN => n17601);
   U15956 : AOI221_X1 port map( B1 => n21775, B2 => n8539, C1 => n21783, C2 => 
                           n8987, A => n17554, ZN => n17546);
   U15957 : OAI22_X1 port map( A1 => n15486, A2 => n21795, B1 => n15452, B2 => 
                           n21791, ZN => n17554);
   U15958 : AOI221_X1 port map( B1 => n21773, B2 => n8537, C1 => n21783, C2 => 
                           n8985, A => n17507, ZN => n17499);
   U15959 : OAI22_X1 port map( A1 => n15485, A2 => n21798, B1 => n15451, B2 => 
                           n21789, ZN => n17507);
   U15960 : AOI221_X1 port map( B1 => n21775, B2 => n8535, C1 => n21784, C2 => 
                           n8983, A => n17460, ZN => n17452);
   U15961 : OAI22_X1 port map( A1 => n15484, A2 => n21799, B1 => n15450, B2 => 
                           n21790, ZN => n17460);
   U15962 : AOI221_X1 port map( B1 => n21776, B2 => n8533, C1 => n21784, C2 => 
                           n8981, A => n17413, ZN => n17405);
   U15963 : OAI22_X1 port map( A1 => n15483, A2 => n21794, B1 => n15449, B2 => 
                           n21786, ZN => n17413);
   U15964 : AOI221_X1 port map( B1 => n21776, B2 => n8531, C1 => n21784, C2 => 
                           n8979, A => n17366, ZN => n17358);
   U15965 : OAI22_X1 port map( A1 => n15482, A2 => n21799, B1 => n15448, B2 => 
                           n21789, ZN => n17366);
   U15966 : AOI221_X1 port map( B1 => n21772, B2 => n8513, C1 => n21780, C2 => 
                           n8961, A => n16943, ZN => n16935);
   U15967 : OAI22_X1 port map( A1 => n15473, A2 => n21795, B1 => n15439, B2 => 
                           n21790, ZN => n16943);
   U15968 : AOI221_X1 port map( B1 => n21772, B2 => n8511, C1 => n21781, C2 => 
                           n8959, A => n16861, ZN => n16838);
   U15969 : OAI22_X1 port map( A1 => n15472, A2 => n21798, B1 => n15438, B2 => 
                           n21787, ZN => n16861);
   U15970 : AOI221_X1 port map( B1 => n20722, B2 => n8956, C1 => n20737, C2 => 
                           n8508, A => n19614, ZN => n19589);
   U15971 : OAI22_X1 port map( A1 => n15606, A2 => n20744, B1 => n4351, B2 => 
                           n20785, ZN => n19614);
   U15972 : AOI221_X1 port map( B1 => n20722, B2 => n8955, C1 => n20737, C2 => 
                           n8507, A => n19577, ZN => n19552);
   U15973 : OAI22_X1 port map( A1 => n15605, A2 => n20745, B1 => n4352, B2 => 
                           n20785, ZN => n19577);
   U15974 : AOI221_X1 port map( B1 => n20723, B2 => n8954, C1 => n20738, C2 => 
                           n8506, A => n19540, ZN => n19515);
   U15975 : OAI22_X1 port map( A1 => n15604, A2 => n20745, B1 => n4353, B2 => 
                           n20789, ZN => n19540);
   U15976 : AOI221_X1 port map( B1 => n20724, B2 => n8953, C1 => n20738, C2 => 
                           n8505, A => n19503, ZN => n19478);
   U15977 : OAI22_X1 port map( A1 => n15603, A2 => n20749, B1 => n4354, B2 => 
                           n20786, ZN => n19503);
   U15978 : AOI221_X1 port map( B1 => n21214, B2 => n8565, C1 => n21221, C2 => 
                           n9013, A => n19477, ZN => n19470);
   U15979 : OAI22_X1 port map( A1 => n15499, A2 => n21243, B1 => n15465, B2 => 
                           n21229, ZN => n19477);
   U15980 : AOI221_X1 port map( B1 => n20724, B2 => n8952, C1 => n20738, C2 => 
                           n8504, A => n19466, ZN => n19441);
   U15981 : OAI22_X1 port map( A1 => n15602, A2 => n20748, B1 => n4355, B2 => 
                           n20787, ZN => n19466);
   U15982 : AOI221_X1 port map( B1 => n20725, B2 => n8951, C1 => n20739, C2 => 
                           n8503, A => n19429, ZN => n19404);
   U15983 : OAI22_X1 port map( A1 => n15601, A2 => n20746, B1 => n4356, B2 => 
                           n20787, ZN => n19429);
   U15984 : AOI221_X1 port map( B1 => n20725, B2 => n8950, C1 => n20739, C2 => 
                           n8502, A => n19392, ZN => n19367);
   U15985 : OAI22_X1 port map( A1 => n15600, A2 => n20746, B1 => n4357, B2 => 
                           n20791, ZN => n19392);
   U15986 : AOI221_X1 port map( B1 => n20725, B2 => n8949, C1 => n20739, C2 => 
                           n8501, A => n19355, ZN => n19330);
   U15987 : OAI22_X1 port map( A1 => n15599, A2 => n20746, B1 => n4358, B2 => 
                           n20785, ZN => n19355);
   U15988 : AOI221_X1 port map( B1 => n20726, B2 => n8948, C1 => n20741, C2 => 
                           n8500, A => n19318, ZN => n19293);
   U15989 : OAI22_X1 port map( A1 => n15598, A2 => n20745, B1 => n4359, B2 => 
                           n20786, ZN => n19318);
   U15990 : AOI221_X1 port map( B1 => n20726, B2 => n8947, C1 => n20742, C2 => 
                           n8499, A => n19281, ZN => n19256);
   U15991 : OAI22_X1 port map( A1 => n15597, A2 => n20747, B1 => n4360, B2 => 
                           n20788, ZN => n19281);
   U15992 : AOI221_X1 port map( B1 => n20727, B2 => n8946, C1 => n20740, C2 => 
                           n8498, A => n19244, ZN => n19219);
   U15993 : OAI22_X1 port map( A1 => n15596, A2 => n20748, B1 => n4361, B2 => 
                           n20789, ZN => n19244);
   U15994 : AOI221_X1 port map( B1 => n20727, B2 => n8945, C1 => n20741, C2 => 
                           n8497, A => n19207, ZN => n19182);
   U15995 : OAI22_X1 port map( A1 => n15595, A2 => n20750, B1 => n4362, B2 => 
                           n20786, ZN => n19207);
   U15996 : AOI221_X1 port map( B1 => n20724, B2 => n8944, C1 => n20741, C2 => 
                           n8496, A => n19170, ZN => n19145);
   U15997 : OAI22_X1 port map( A1 => n15594, A2 => n20746, B1 => n4363, B2 => 
                           n20787, ZN => n19170);
   U15998 : AOI221_X1 port map( B1 => n20726, B2 => n8943, C1 => n20742, C2 => 
                           n8495, A => n19133, ZN => n19108);
   U15999 : OAI22_X1 port map( A1 => n15593, A2 => n20746, B1 => n4364, B2 => 
                           n20787, ZN => n19133);
   U16000 : AOI221_X1 port map( B1 => n20727, B2 => n8942, C1 => n20740, C2 => 
                           n8494, A => n19096, ZN => n19071);
   U16001 : OAI22_X1 port map( A1 => n15592, A2 => n20749, B1 => n4365, B2 => 
                           n20790, ZN => n19096);
   U16002 : AOI221_X1 port map( B1 => n20725, B2 => n8941, C1 => n20741, C2 => 
                           n8493, A => n19059, ZN => n19034);
   U16003 : OAI22_X1 port map( A1 => n15591, A2 => n20746, B1 => n4366, B2 => 
                           n20788, ZN => n19059);
   U16004 : AOI221_X1 port map( B1 => n20726, B2 => n8940, C1 => n20741, C2 => 
                           n8492, A => n19022, ZN => n18997);
   U16005 : OAI22_X1 port map( A1 => n15590, A2 => n20744, B1 => n4367, B2 => 
                           n20785, ZN => n19022);
   U16006 : AOI221_X1 port map( B1 => n20728, B2 => n8939, C1 => n20742, C2 => 
                           n8491, A => n18985, ZN => n18960);
   U16007 : OAI22_X1 port map( A1 => n15589, A2 => n20747, B1 => n4368, B2 => 
                           n20788, ZN => n18985);
   U16008 : AOI221_X1 port map( B1 => n20728, B2 => n8938, C1 => n20742, C2 => 
                           n8490, A => n18948, ZN => n18923);
   U16009 : OAI22_X1 port map( A1 => n15588, A2 => n20748, B1 => n4369, B2 => 
                           n20788, ZN => n18948);
   U16010 : AOI221_X1 port map( B1 => n20728, B2 => n8937, C1 => n20742, C2 => 
                           n8489, A => n18911, ZN => n18886);
   U16011 : OAI22_X1 port map( A1 => n15587, A2 => n20748, B1 => n4370, B2 => 
                           n20789, ZN => n18911);
   U16012 : AOI221_X1 port map( B1 => n20728, B2 => n8936, C1 => n20742, C2 => 
                           n8488, A => n18874, ZN => n18849);
   U16013 : OAI22_X1 port map( A1 => n15586, A2 => n20747, B1 => n4371, B2 => 
                           n20791, ZN => n18874);
   U16014 : AOI221_X1 port map( B1 => n20722, B2 => n8935, C1 => n20737, C2 => 
                           n8487, A => n18837, ZN => n18812);
   U16015 : OAI22_X1 port map( A1 => n15585, A2 => n20749, B1 => n4372, B2 => 
                           n20789, ZN => n18837);
   U16016 : AOI221_X1 port map( B1 => n21219, B2 => n8529, C1 => n21221, C2 => 
                           n8977, A => n18811, ZN => n18804);
   U16017 : OAI22_X1 port map( A1 => n15481, A2 => n21241, B1 => n15447, B2 => 
                           n21233, ZN => n18811);
   U16018 : AOI221_X1 port map( B1 => n20722, B2 => n8934, C1 => n20737, C2 => 
                           n8486, A => n18800, ZN => n18775);
   U16019 : OAI22_X1 port map( A1 => n15584, A2 => n20749, B1 => n4373, B2 => 
                           n20790, ZN => n18800);
   U16020 : AOI221_X1 port map( B1 => n21219, B2 => n8527, C1 => n21223, C2 => 
                           n8975, A => n18774, ZN => n18767);
   U16021 : OAI22_X1 port map( A1 => n15480, A2 => n21242, B1 => n15446, B2 => 
                           n21233, ZN => n18774);
   U16022 : AOI221_X1 port map( B1 => n20722, B2 => n8933, C1 => n20740, C2 => 
                           n8485, A => n18763, ZN => n18738);
   U16023 : OAI22_X1 port map( A1 => n15583, A2 => n20750, B1 => n4374, B2 => 
                           n20790, ZN => n18763);
   U16024 : AOI221_X1 port map( B1 => n21213, B2 => n8525, C1 => n21225, C2 => 
                           n8973, A => n18737, ZN => n18730);
   U16025 : OAI22_X1 port map( A1 => n15479, A2 => n21243, B1 => n15445, B2 => 
                           n21234, ZN => n18737);
   U16026 : AOI221_X1 port map( B1 => n20723, B2 => n8932, C1 => n20738, C2 => 
                           n8484, A => n18726, ZN => n18701);
   U16027 : OAI22_X1 port map( A1 => n15582, A2 => n20750, B1 => n4375, B2 => 
                           n20791, ZN => n18726);
   U16028 : AOI221_X1 port map( B1 => n21214, B2 => n8523, C1 => n21225, C2 => 
                           n8971, A => n18700, ZN => n18693);
   U16029 : OAI22_X1 port map( A1 => n15478, A2 => n21243, B1 => n15444, B2 => 
                           n21234, ZN => n18700);
   U16030 : AOI221_X1 port map( B1 => n20724, B2 => n8931, C1 => n20738, C2 => 
                           n8483, A => n18689, ZN => n18664);
   U16031 : OAI22_X1 port map( A1 => n15581, A2 => n20749, B1 => n4376, B2 => 
                           n20790, ZN => n18689);
   U16032 : AOI221_X1 port map( B1 => n21213, B2 => n8521, C1 => n21221, C2 => 
                           n8969, A => n18663, ZN => n18656);
   U16033 : OAI22_X1 port map( A1 => n15477, A2 => n21243, B1 => n15443, B2 => 
                           n21235, ZN => n18663);
   U16034 : AOI221_X1 port map( B1 => n20723, B2 => n8930, C1 => n20740, C2 => 
                           n8482, A => n18652, ZN => n18627);
   U16035 : OAI22_X1 port map( A1 => n15580, A2 => n20750, B1 => n4377, B2 => 
                           n20791, ZN => n18652);
   U16036 : AOI221_X1 port map( B1 => n21214, B2 => n8519, C1 => n21222, C2 => 
                           n8967, A => n18626, ZN => n18619);
   U16037 : OAI22_X1 port map( A1 => n15476, A2 => n21243, B1 => n15442, B2 => 
                           n21235, ZN => n18626);
   U16038 : AOI221_X1 port map( B1 => n20725, B2 => n8929, C1 => n20739, C2 => 
                           n8481, A => n18615, ZN => n18590);
   U16039 : OAI22_X1 port map( A1 => n15579, A2 => n20747, B1 => n4378, B2 => 
                           n20790, ZN => n18615);
   U16040 : AOI221_X1 port map( B1 => n21215, B2 => n8517, C1 => n21223, C2 => 
                           n8965, A => n18589, ZN => n18582);
   U16041 : OAI22_X1 port map( A1 => n15475, A2 => n21241, B1 => n15441, B2 => 
                           n21235, ZN => n18589);
   U16042 : AOI221_X1 port map( B1 => n20725, B2 => n8928, C1 => n20739, C2 => 
                           n8480, A => n18578, ZN => n18553);
   U16043 : OAI22_X1 port map( A1 => n15578, A2 => n20744, B1 => n4379, B2 => 
                           n20785, ZN => n18578);
   U16044 : AOI221_X1 port map( B1 => n21216, B2 => n8515, C1 => n21222, C2 => 
                           n8963, A => n18552, ZN => n18545);
   U16045 : OAI22_X1 port map( A1 => n15474, A2 => n21243, B1 => n15440, B2 => 
                           n21234, ZN => n18552);
   U16046 : AOI221_X1 port map( B1 => n20727, B2 => n8927, C1 => n20737, C2 => 
                           n8479, A => n18541, ZN => n18516);
   U16047 : OAI22_X1 port map( A1 => n15577, A2 => n20745, B1 => n4380, B2 => 
                           n20786, ZN => n18541);
   U16048 : AOI221_X1 port map( B1 => n20727, B2 => n8926, C1 => n20740, C2 => 
                           n8478, A => n18502, ZN => n18446);
   U16049 : OAI22_X1 port map( A1 => n15576, A2 => n20744, B1 => n4381, B2 => 
                           n20791, ZN => n18502);
   U16050 : AOI221_X1 port map( B1 => n21279, B2 => n8956, C1 => n21294, C2 => 
                           n8508, A => n18341, ZN => n18307);
   U16051 : OAI22_X1 port map( A1 => n15606, A2 => n21301, B1 => n4351, B2 => 
                           n21342, ZN => n18341);
   U16052 : AOI221_X1 port map( B1 => n21279, B2 => n8955, C1 => n21294, C2 => 
                           n8507, A => n18294, ZN => n18260);
   U16053 : OAI22_X1 port map( A1 => n15605, A2 => n21302, B1 => n4352, B2 => 
                           n21342, ZN => n18294);
   U16054 : AOI221_X1 port map( B1 => n21280, B2 => n8954, C1 => n21295, C2 => 
                           n8506, A => n18247, ZN => n18213);
   U16055 : OAI22_X1 port map( A1 => n15604, A2 => n21302, B1 => n4353, B2 => 
                           n21346, ZN => n18247);
   U16056 : AOI221_X1 port map( B1 => n21281, B2 => n8953, C1 => n21295, C2 => 
                           n8505, A => n18200, ZN => n18166);
   U16057 : OAI22_X1 port map( A1 => n15603, A2 => n21306, B1 => n4354, B2 => 
                           n21343, ZN => n18200);
   U16058 : AOI221_X1 port map( B1 => n21771, B2 => n8565, C1 => n21778, C2 => 
                           n9013, A => n18165, ZN => n18157);
   U16059 : OAI22_X1 port map( A1 => n15499, A2 => n21800, B1 => n15465, B2 => 
                           n21786, ZN => n18165);
   U16060 : AOI221_X1 port map( B1 => n21281, B2 => n8952, C1 => n21295, C2 => 
                           n8504, A => n18153, ZN => n18119);
   U16061 : OAI22_X1 port map( A1 => n15602, A2 => n21305, B1 => n4355, B2 => 
                           n21344, ZN => n18153);
   U16062 : AOI221_X1 port map( B1 => n21282, B2 => n8951, C1 => n21296, C2 => 
                           n8503, A => n18106, ZN => n18072);
   U16063 : OAI22_X1 port map( A1 => n15601, A2 => n21303, B1 => n4356, B2 => 
                           n21344, ZN => n18106);
   U16064 : AOI221_X1 port map( B1 => n21282, B2 => n8950, C1 => n21296, C2 => 
                           n8502, A => n18059, ZN => n18025);
   U16065 : OAI22_X1 port map( A1 => n15600, A2 => n21303, B1 => n4357, B2 => 
                           n21348, ZN => n18059);
   U16066 : AOI221_X1 port map( B1 => n21282, B2 => n8949, C1 => n21296, C2 => 
                           n8501, A => n18012, ZN => n17978);
   U16067 : OAI22_X1 port map( A1 => n15599, A2 => n21303, B1 => n4358, B2 => 
                           n21342, ZN => n18012);
   U16068 : AOI221_X1 port map( B1 => n21283, B2 => n8948, C1 => n21298, C2 => 
                           n8500, A => n17965, ZN => n17931);
   U16069 : OAI22_X1 port map( A1 => n15598, A2 => n21302, B1 => n4359, B2 => 
                           n21343, ZN => n17965);
   U16070 : AOI221_X1 port map( B1 => n21283, B2 => n8947, C1 => n21299, C2 => 
                           n8499, A => n17918, ZN => n17884);
   U16071 : OAI22_X1 port map( A1 => n15597, A2 => n21304, B1 => n4360, B2 => 
                           n21345, ZN => n17918);
   U16072 : AOI221_X1 port map( B1 => n21284, B2 => n8946, C1 => n21297, C2 => 
                           n8498, A => n17871, ZN => n17837);
   U16073 : OAI22_X1 port map( A1 => n15596, A2 => n21305, B1 => n4361, B2 => 
                           n21346, ZN => n17871);
   U16074 : AOI221_X1 port map( B1 => n21284, B2 => n8945, C1 => n21298, C2 => 
                           n8497, A => n17824, ZN => n17790);
   U16075 : OAI22_X1 port map( A1 => n15595, A2 => n21307, B1 => n4362, B2 => 
                           n21343, ZN => n17824);
   U16076 : AOI221_X1 port map( B1 => n21281, B2 => n8944, C1 => n21298, C2 => 
                           n8496, A => n17777, ZN => n17743);
   U16077 : OAI22_X1 port map( A1 => n15594, A2 => n21303, B1 => n4363, B2 => 
                           n21344, ZN => n17777);
   U16078 : AOI221_X1 port map( B1 => n21283, B2 => n8943, C1 => n21299, C2 => 
                           n8495, A => n17730, ZN => n17696);
   U16079 : OAI22_X1 port map( A1 => n15593, A2 => n21303, B1 => n4364, B2 => 
                           n21344, ZN => n17730);
   U16080 : AOI221_X1 port map( B1 => n21284, B2 => n8942, C1 => n21297, C2 => 
                           n8494, A => n17683, ZN => n17649);
   U16081 : OAI22_X1 port map( A1 => n15592, A2 => n21306, B1 => n4365, B2 => 
                           n21347, ZN => n17683);
   U16082 : AOI221_X1 port map( B1 => n21282, B2 => n8941, C1 => n21298, C2 => 
                           n8493, A => n17636, ZN => n17602);
   U16083 : OAI22_X1 port map( A1 => n15591, A2 => n21303, B1 => n4366, B2 => 
                           n21345, ZN => n17636);
   U16084 : AOI221_X1 port map( B1 => n21283, B2 => n8940, C1 => n21298, C2 => 
                           n8492, A => n17589, ZN => n17555);
   U16085 : OAI22_X1 port map( A1 => n15590, A2 => n21301, B1 => n4367, B2 => 
                           n21342, ZN => n17589);
   U16086 : AOI221_X1 port map( B1 => n21285, B2 => n8939, C1 => n21299, C2 => 
                           n8491, A => n17542, ZN => n17508);
   U16087 : OAI22_X1 port map( A1 => n15589, A2 => n21304, B1 => n4368, B2 => 
                           n21345, ZN => n17542);
   U16088 : AOI221_X1 port map( B1 => n21285, B2 => n8938, C1 => n21299, C2 => 
                           n8490, A => n17495, ZN => n17461);
   U16089 : OAI22_X1 port map( A1 => n15588, A2 => n21305, B1 => n4369, B2 => 
                           n21345, ZN => n17495);
   U16090 : AOI221_X1 port map( B1 => n21285, B2 => n8937, C1 => n21299, C2 => 
                           n8489, A => n17448, ZN => n17414);
   U16091 : OAI22_X1 port map( A1 => n15587, A2 => n21305, B1 => n4370, B2 => 
                           n21346, ZN => n17448);
   U16092 : AOI221_X1 port map( B1 => n21285, B2 => n8936, C1 => n21299, C2 => 
                           n8488, A => n17401, ZN => n17367);
   U16093 : OAI22_X1 port map( A1 => n15586, A2 => n21304, B1 => n4371, B2 => 
                           n21348, ZN => n17401);
   U16094 : AOI221_X1 port map( B1 => n21279, B2 => n8935, C1 => n21294, C2 => 
                           n8487, A => n17354, ZN => n17320);
   U16095 : OAI22_X1 port map( A1 => n15585, A2 => n21306, B1 => n4372, B2 => 
                           n21346, ZN => n17354);
   U16096 : AOI221_X1 port map( B1 => n21776, B2 => n8529, C1 => n21778, C2 => 
                           n8977, A => n17319, ZN => n17311);
   U16097 : OAI22_X1 port map( A1 => n15481, A2 => n21798, B1 => n15447, B2 => 
                           n21790, ZN => n17319);
   U16098 : AOI221_X1 port map( B1 => n21279, B2 => n8934, C1 => n21294, C2 => 
                           n8486, A => n17307, ZN => n17273);
   U16099 : OAI22_X1 port map( A1 => n15584, A2 => n21306, B1 => n4373, B2 => 
                           n21347, ZN => n17307);
   U16100 : AOI221_X1 port map( B1 => n21776, B2 => n8527, C1 => n21780, C2 => 
                           n8975, A => n17272, ZN => n17264);
   U16101 : OAI22_X1 port map( A1 => n15480, A2 => n21799, B1 => n15446, B2 => 
                           n21790, ZN => n17272);
   U16102 : AOI221_X1 port map( B1 => n21279, B2 => n8933, C1 => n21297, C2 => 
                           n8485, A => n17260, ZN => n17226);
   U16103 : OAI22_X1 port map( A1 => n15583, A2 => n21307, B1 => n4374, B2 => 
                           n21347, ZN => n17260);
   U16104 : AOI221_X1 port map( B1 => n21770, B2 => n8525, C1 => n21782, C2 => 
                           n8973, A => n17225, ZN => n17217);
   U16105 : OAI22_X1 port map( A1 => n15479, A2 => n21800, B1 => n15445, B2 => 
                           n21791, ZN => n17225);
   U16106 : AOI221_X1 port map( B1 => n21280, B2 => n8932, C1 => n21295, C2 => 
                           n8484, A => n17213, ZN => n17179);
   U16107 : OAI22_X1 port map( A1 => n15582, A2 => n21307, B1 => n4375, B2 => 
                           n21348, ZN => n17213);
   U16108 : AOI221_X1 port map( B1 => n21771, B2 => n8523, C1 => n21782, C2 => 
                           n8971, A => n17178, ZN => n17170);
   U16109 : OAI22_X1 port map( A1 => n15478, A2 => n21800, B1 => n15444, B2 => 
                           n21791, ZN => n17178);
   U16110 : AOI221_X1 port map( B1 => n21281, B2 => n8931, C1 => n21295, C2 => 
                           n8483, A => n17166, ZN => n17132);
   U16111 : OAI22_X1 port map( A1 => n15581, A2 => n21306, B1 => n4376, B2 => 
                           n21347, ZN => n17166);
   U16112 : AOI221_X1 port map( B1 => n21770, B2 => n8521, C1 => n21778, C2 => 
                           n8969, A => n17131, ZN => n17123);
   U16113 : OAI22_X1 port map( A1 => n15477, A2 => n21800, B1 => n15443, B2 => 
                           n21792, ZN => n17131);
   U16114 : AOI221_X1 port map( B1 => n21280, B2 => n8930, C1 => n21297, C2 => 
                           n8482, A => n17119, ZN => n17085);
   U16115 : OAI22_X1 port map( A1 => n15580, A2 => n21307, B1 => n4377, B2 => 
                           n21348, ZN => n17119);
   U16116 : AOI221_X1 port map( B1 => n21771, B2 => n8519, C1 => n21779, C2 => 
                           n8967, A => n17084, ZN => n17076);
   U16117 : OAI22_X1 port map( A1 => n15476, A2 => n21800, B1 => n15442, B2 => 
                           n21792, ZN => n17084);
   U16118 : AOI221_X1 port map( B1 => n21282, B2 => n8929, C1 => n21296, C2 => 
                           n8481, A => n17072, ZN => n17038);
   U16119 : OAI22_X1 port map( A1 => n15579, A2 => n21304, B1 => n4378, B2 => 
                           n21347, ZN => n17072);
   U16120 : AOI221_X1 port map( B1 => n21772, B2 => n8517, C1 => n21780, C2 => 
                           n8965, A => n17037, ZN => n17029);
   U16121 : OAI22_X1 port map( A1 => n15475, A2 => n21798, B1 => n15441, B2 => 
                           n21792, ZN => n17037);
   U16122 : AOI221_X1 port map( B1 => n21282, B2 => n8928, C1 => n21296, C2 => 
                           n8480, A => n17025, ZN => n16991);
   U16123 : OAI22_X1 port map( A1 => n15578, A2 => n21301, B1 => n4379, B2 => 
                           n21342, ZN => n17025);
   U16124 : AOI221_X1 port map( B1 => n21773, B2 => n8515, C1 => n21779, C2 => 
                           n8963, A => n16990, ZN => n16982);
   U16125 : OAI22_X1 port map( A1 => n15474, A2 => n21800, B1 => n15440, B2 => 
                           n21791, ZN => n16990);
   U16126 : AOI221_X1 port map( B1 => n21284, B2 => n8927, C1 => n21294, C2 => 
                           n8479, A => n16978, ZN => n16944);
   U16127 : OAI22_X1 port map( A1 => n15577, A2 => n21302, B1 => n4380, B2 => 
                           n21343, ZN => n16978);
   U16128 : AOI221_X1 port map( B1 => n21284, B2 => n8926, C1 => n21297, C2 => 
                           n8478, A => n16929, ZN => n16864);
   U16129 : OAI22_X1 port map( A1 => n15576, A2 => n21301, B1 => n4381, B2 => 
                           n21348, ZN => n16929);
   U16130 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n19671,
                           ZN => n19675);
   U16131 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n18406,
                           ZN => n18411);
   U16132 : NOR3_X1 port map( A1 => n19671, A2 => ADD_RD1(3), A3 => n19666, ZN 
                           => n19678);
   U16133 : NOR3_X1 port map( A1 => n18406, A2 => ADD_RD2(3), A3 => n18400, ZN 
                           => n18415);
   U16134 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(5), A3 => n19666,
                           ZN => n19667);
   U16135 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(5), A3 => n18400,
                           ZN => n18401);
   U16136 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n16795, ZN => n15191);
   U16137 : NAND2_X1 port map( A1 => ADD_WR(0), A2 => n16794, ZN => n15156);
   U16138 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), ZN => n15226);
   U16139 : OAI221_X1 port map( B1 => n15400, B2 => n21030, C1 => n15262, C2 =>
                           n21032, A => n19651, ZN => n19650);
   U16140 : AOI22_X1 port map( A1 => n21038, A2 => n9821, B1 => n21078, B2 => 
                           n19937, ZN => n19651);
   U16141 : OAI221_X1 port map( B1 => n15435, B2 => n21029, C1 => n15297, C2 =>
                           n21037, A => n19659, ZN => n19658);
   U16142 : AOI22_X1 port map( A1 => n21068, A2 => n9853, B1 => n21077, B2 => 
                           n19938, ZN => n19659);
   U16143 : OAI221_X1 port map( B1 => n15399, B2 => n21026, C1 => n15261, C2 =>
                           n21034, A => n19600, ZN => n19599);
   U16144 : AOI22_X1 port map( A1 => n21047, A2 => n9820, B1 => n21080, B2 => 
                           n19939, ZN => n19600);
   U16145 : OAI221_X1 port map( B1 => n15434, B2 => n21031, C1 => n15296, C2 =>
                           n21033, A => n19608, ZN => n19607);
   U16146 : AOI22_X1 port map( A1 => n21046, A2 => n9852, B1 => n21079, B2 => 
                           n19940, ZN => n19608);
   U16147 : OAI221_X1 port map( B1 => n15398, B2 => n21026, C1 => n15260, C2 =>
                           n21032, A => n19563, ZN => n19562);
   U16148 : AOI22_X1 port map( A1 => n21049, A2 => n9819, B1 => n21082, B2 => 
                           n19941, ZN => n19563);
   U16149 : OAI221_X1 port map( B1 => n15433, B2 => n21031, C1 => n15295, C2 =>
                           n21035, A => n19571, ZN => n19570);
   U16150 : AOI22_X1 port map( A1 => n21048, A2 => n9851, B1 => n21081, B2 => 
                           n19942, ZN => n19571);
   U16151 : OAI221_X1 port map( B1 => n15397, B2 => n21028, C1 => n15259, C2 =>
                           n21037, A => n19526, ZN => n19525);
   U16152 : AOI22_X1 port map( A1 => n21051, A2 => n9818, B1 => n21084, B2 => 
                           n19943, ZN => n19526);
   U16153 : OAI221_X1 port map( B1 => n15432, B2 => n21027, C1 => n15294, C2 =>
                           n21036, A => n19534, ZN => n19533);
   U16154 : AOI22_X1 port map( A1 => n21050, A2 => n9850, B1 => n21083, B2 => 
                           n19944, ZN => n19534);
   U16155 : OAI221_X1 port map( B1 => n15396, B2 => n21030, C1 => n15258, C2 =>
                           n21033, A => n19489, ZN => n19488);
   U16156 : AOI22_X1 port map( A1 => n21053, A2 => n9817, B1 => n21086, B2 => 
                           n19945, ZN => n19489);
   U16157 : OAI221_X1 port map( B1 => n15431, B2 => n21029, C1 => n15293, C2 =>
                           n21032, A => n19497, ZN => n19496);
   U16158 : AOI22_X1 port map( A1 => n21052, A2 => n9849, B1 => n21085, B2 => 
                           n19946, ZN => n19497);
   U16159 : OAI221_X1 port map( B1 => n15395, B2 => n21027, C1 => n15257, C2 =>
                           n21033, A => n19452, ZN => n19451);
   U16160 : AOI22_X1 port map( A1 => n21055, A2 => n9816, B1 => n21088, B2 => 
                           n19947, ZN => n19452);
   U16161 : OAI221_X1 port map( B1 => n15430, B2 => n21026, C1 => n15292, C2 =>
                           n21034, A => n19460, ZN => n19459);
   U16162 : AOI22_X1 port map( A1 => n21054, A2 => n9848, B1 => n21087, B2 => 
                           n19948, ZN => n19460);
   U16163 : OAI221_X1 port map( B1 => n15394, B2 => n21026, C1 => n15256, C2 =>
                           n21036, A => n19415, ZN => n19414);
   U16164 : AOI22_X1 port map( A1 => n21057, A2 => n9815, B1 => n21090, B2 => 
                           n19949, ZN => n19415);
   U16165 : OAI221_X1 port map( B1 => n15429, B2 => n21031, C1 => n15291, C2 =>
                           n21035, A => n19423, ZN => n19422);
   U16166 : AOI22_X1 port map( A1 => n21056, A2 => n9847, B1 => n21089, B2 => 
                           n19950, ZN => n19423);
   U16167 : OAI221_X1 port map( B1 => n15393, B2 => n21028, C1 => n15255, C2 =>
                           n21032, A => n19378, ZN => n19377);
   U16168 : AOI22_X1 port map( A1 => n21062, A2 => n9814, B1 => n21092, B2 => 
                           n19951, ZN => n19378);
   U16169 : OAI221_X1 port map( B1 => n15428, B2 => n21027, C1 => n15290, C2 =>
                           n21037, A => n19386, ZN => n19385);
   U16170 : AOI22_X1 port map( A1 => n21062, A2 => n9846, B1 => n21091, B2 => 
                           n19952, ZN => n19386);
   U16171 : OAI221_X1 port map( B1 => n15392, B2 => n21028, C1 => n15254, C2 =>
                           n21034, A => n19341, ZN => n19340);
   U16172 : AOI22_X1 port map( A1 => n21063, A2 => n9813, B1 => n21092, B2 => 
                           n19953, ZN => n19341);
   U16173 : OAI221_X1 port map( B1 => n15427, B2 => n21027, C1 => n15289, C2 =>
                           n21033, A => n19349, ZN => n19348);
   U16174 : AOI22_X1 port map( A1 => n21062, A2 => n9845, B1 => n21101, B2 => 
                           n19954, ZN => n19349);
   U16175 : OAI221_X1 port map( B1 => n15391, B2 => n21030, C1 => n15253, C2 =>
                           n21035, A => n19304, ZN => n19303);
   U16176 : AOI22_X1 port map( A1 => n21064, A2 => n9812, B1 => n21096, B2 => 
                           n19955, ZN => n19304);
   U16177 : OAI221_X1 port map( B1 => n15426, B2 => n21029, C1 => n15288, C2 =>
                           n21034, A => n19312, ZN => n19311);
   U16178 : AOI22_X1 port map( A1 => n21063, A2 => n9844, B1 => n21096, B2 => 
                           n19956, ZN => n19312);
   U16179 : OAI221_X1 port map( B1 => n15390, B2 => n21026, C1 => n15252, C2 =>
                           n21037, A => n19267, ZN => n19266);
   U16180 : AOI22_X1 port map( A1 => n21065, A2 => n9811, B1 => n21097, B2 => 
                           n19957, ZN => n19267);
   U16181 : OAI221_X1 port map( B1 => n15425, B2 => n21031, C1 => n15287, C2 =>
                           n21036, A => n19275, ZN => n19274);
   U16182 : AOI22_X1 port map( A1 => n21066, A2 => n9843, B1 => n21096, B2 => 
                           n19958, ZN => n19275);
   U16183 : OAI221_X1 port map( B1 => n15389, B2 => n21029, C1 => n15251, C2 =>
                           n21035, A => n19230, ZN => n19229);
   U16184 : AOI22_X1 port map( A1 => n21067, A2 => n9810, B1 => n21098, B2 => 
                           n19959, ZN => n19230);
   U16185 : OAI221_X1 port map( B1 => n15424, B2 => n21028, C1 => n15286, C2 =>
                           n21032, A => n19238, ZN => n19237);
   U16186 : AOI22_X1 port map( A1 => n21066, A2 => n9842, B1 => n21097, B2 => 
                           n19960, ZN => n19238);
   U16187 : OAI221_X1 port map( B1 => n15388, B2 => n21028, C1 => n15250, C2 =>
                           n21034, A => n19193, ZN => n19192);
   U16188 : AOI22_X1 port map( A1 => n21068, A2 => n9809, B1 => n21099, B2 => 
                           n19961, ZN => n19193);
   U16189 : OAI221_X1 port map( B1 => n15423, B2 => n21027, C1 => n15285, C2 =>
                           n21033, A => n19201, ZN => n19200);
   U16190 : AOI22_X1 port map( A1 => n21068, A2 => n9841, B1 => n21099, B2 => 
                           n19962, ZN => n19201);
   U16191 : OAI221_X1 port map( B1 => n15387, B2 => n21030, C1 => n15249, C2 =>
                           n21036, A => n19156, ZN => n19155);
   U16192 : AOI22_X1 port map( A1 => n21069, A2 => n9808, B1 => n21100, B2 => 
                           n19963, ZN => n19156);
   U16193 : OAI221_X1 port map( B1 => n15422, B2 => n21029, C1 => n15284, C2 =>
                           n21035, A => n19164, ZN => n19163);
   U16194 : AOI22_X1 port map( A1 => n21069, A2 => n9840, B1 => n21099, B2 => 
                           n19964, ZN => n19164);
   U16195 : OAI221_X1 port map( B1 => n15386, B2 => n21030, C1 => n15248, C2 =>
                           n21036, A => n19119, ZN => n19118);
   U16196 : AOI22_X1 port map( A1 => n21065, A2 => n9807, B1 => n21098, B2 => 
                           n19965, ZN => n19119);
   U16197 : OAI221_X1 port map( B1 => n15421, B2 => n21029, C1 => n15283, C2 =>
                           n21037, A => n19127, ZN => n19126);
   U16198 : AOI22_X1 port map( A1 => n21045, A2 => n9839, B1 => n21097, B2 => 
                           n19966, ZN => n19127);
   U16199 : OAI221_X1 port map( B1 => n15385, B2 => n21026, C1 => n15247, C2 =>
                           n21033, A => n19082, ZN => n19081);
   U16200 : AOI22_X1 port map( A1 => n21065, A2 => n9806, B1 => n21099, B2 => 
                           n19967, ZN => n19082);
   U16201 : OAI221_X1 port map( B1 => n15420, B2 => n21031, C1 => n15282, C2 =>
                           n21032, A => n19090, ZN => n19089);
   U16202 : AOI22_X1 port map( A1 => n21066, A2 => n9838, B1 => n21099, B2 => 
                           n19968, ZN => n19090);
   U16203 : OAI221_X1 port map( B1 => n15384, B2 => n21028, C1 => n15246, C2 =>
                           n21035, A => n19045, ZN => n19044);
   U16204 : AOI22_X1 port map( A1 => n21067, A2 => n9805, B1 => n21100, B2 => 
                           n19969, ZN => n19045);
   U16205 : OAI221_X1 port map( B1 => n15419, B2 => n21027, C1 => n15281, C2 =>
                           n21034, A => n19053, ZN => n19052);
   U16206 : AOI22_X1 port map( A1 => n21066, A2 => n9837, B1 => n21099, B2 => 
                           n19970, ZN => n19053);
   U16207 : OAI221_X1 port map( B1 => n15383, B2 => n21031, C1 => n15245, C2 =>
                           n21037, A => n19008, ZN => n19007);
   U16208 : AOI22_X1 port map( A1 => n21068, A2 => n9804, B1 => n21098, B2 => 
                           n19971, ZN => n19008);
   U16209 : OAI221_X1 port map( B1 => n15418, B2 => n21030, C1 => n15280, C2 =>
                           n21036, A => n19016, ZN => n19015);
   U16210 : AOI22_X1 port map( A1 => n21067, A2 => n9836, B1 => n21096, B2 => 
                           n19972, ZN => n19016);
   U16211 : OAI221_X1 port map( B1 => n15417, B2 => n21029, C1 => n15279, C2 =>
                           n21037, A => n18979, ZN => n18978);
   U16212 : AOI22_X1 port map( A1 => n21069, A2 => n9835, B1 => n21101, B2 => 
                           n19973, ZN => n18979);
   U16213 : OAI221_X1 port map( B1 => n15416, B2 => n21031, C1 => n15278, C2 =>
                           n21033, A => n18942, ZN => n18941);
   U16214 : AOI22_X1 port map( A1 => n21070, A2 => n9834, B1 => n21102, B2 => 
                           n19974, ZN => n18942);
   U16215 : OAI221_X1 port map( B1 => n15380, B2 => n21026, C1 => n15242, C2 =>
                           n21032, A => n18897, ZN => n18896);
   U16216 : AOI22_X1 port map( A1 => n21044, A2 => n9801, B1 => n21103, B2 => 
                           n19975, ZN => n18897);
   U16217 : OAI221_X1 port map( B1 => n15415, B2 => n21031, C1 => n15277, C2 =>
                           n21035, A => n18905, ZN => n18904);
   U16218 : AOI22_X1 port map( A1 => n21067, A2 => n9833, B1 => n21102, B2 => 
                           n19976, ZN => n18905);
   U16219 : OAI221_X1 port map( B1 => n15414, B2 => n21027, C1 => n15276, C2 =>
                           n21036, A => n18868, ZN => n18867);
   U16220 : AOI22_X1 port map( A1 => n21045, A2 => n9832, B1 => n21103, B2 => 
                           n19977, ZN => n18868);
   U16221 : OAI221_X1 port map( B1 => n15378, B2 => n21030, C1 => n15240, C2 =>
                           n21033, A => n18823, ZN => n18822);
   U16222 : AOI22_X1 port map( A1 => n21070, A2 => n9799, B1 => n21078, B2 => 
                           n19978, ZN => n18823);
   U16223 : OAI221_X1 port map( B1 => n15413, B2 => n21029, C1 => n15275, C2 =>
                           n21032, A => n18831, ZN => n18830);
   U16224 : AOI22_X1 port map( A1 => n21066, A2 => n9831, B1 => n21077, B2 => 
                           n19979, ZN => n18831);
   U16225 : OAI221_X1 port map( B1 => n15377, B2 => n21027, C1 => n15239, C2 =>
                           n21033, A => n18786, ZN => n18785);
   U16226 : AOI22_X1 port map( A1 => n21047, A2 => n9798, B1 => n21080, B2 => 
                           n19980, ZN => n18786);
   U16227 : OAI221_X1 port map( B1 => n15412, B2 => n21026, C1 => n15274, C2 =>
                           n21034, A => n18794, ZN => n18793);
   U16228 : AOI22_X1 port map( A1 => n21046, A2 => n9830, B1 => n21079, B2 => 
                           n19981, ZN => n18794);
   U16229 : OAI221_X1 port map( B1 => n15376, B2 => n21026, C1 => n15238, C2 =>
                           n21036, A => n18749, ZN => n18748);
   U16230 : AOI22_X1 port map( A1 => n21049, A2 => n9797, B1 => n21082, B2 => 
                           n19982, ZN => n18749);
   U16231 : OAI221_X1 port map( B1 => n15411, B2 => n21031, C1 => n15273, C2 =>
                           n21035, A => n18757, ZN => n18756);
   U16232 : AOI22_X1 port map( A1 => n21048, A2 => n9829, B1 => n21081, B2 => 
                           n19983, ZN => n18757);
   U16233 : OAI221_X1 port map( B1 => n15375, B2 => n21028, C1 => n15237, C2 =>
                           n21032, A => n18712, ZN => n18711);
   U16234 : AOI22_X1 port map( A1 => n21051, A2 => n9796, B1 => n21084, B2 => 
                           n19984, ZN => n18712);
   U16235 : OAI221_X1 port map( B1 => n15410, B2 => n21027, C1 => n15272, C2 =>
                           n21037, A => n18720, ZN => n18719);
   U16236 : AOI22_X1 port map( A1 => n21050, A2 => n9828, B1 => n21083, B2 => 
                           n19985, ZN => n18720);
   U16237 : OAI221_X1 port map( B1 => n15374, B2 => n21028, C1 => n15236, C2 =>
                           n21034, A => n18675, ZN => n18674);
   U16238 : AOI22_X1 port map( A1 => n21053, A2 => n9795, B1 => n21086, B2 => 
                           n19986, ZN => n18675);
   U16239 : OAI221_X1 port map( B1 => n15409, B2 => n21027, C1 => n15271, C2 =>
                           n21033, A => n18683, ZN => n18682);
   U16240 : AOI22_X1 port map( A1 => n21052, A2 => n9827, B1 => n21085, B2 => 
                           n19987, ZN => n18683);
   U16241 : OAI221_X1 port map( B1 => n15373, B2 => n21030, C1 => n15235, C2 =>
                           n21035, A => n18638, ZN => n18637);
   U16242 : AOI22_X1 port map( A1 => n21055, A2 => n9794, B1 => n21088, B2 => 
                           n19988, ZN => n18638);
   U16243 : OAI221_X1 port map( B1 => n15408, B2 => n21029, C1 => n15270, C2 =>
                           n21034, A => n18646, ZN => n18645);
   U16244 : AOI22_X1 port map( A1 => n21054, A2 => n9826, B1 => n21087, B2 => 
                           n19989, ZN => n18646);
   U16245 : OAI221_X1 port map( B1 => n15372, B2 => n21026, C1 => n15234, C2 =>
                           n21037, A => n18601, ZN => n18600);
   U16246 : AOI22_X1 port map( A1 => n21057, A2 => n9793, B1 => n21090, B2 => 
                           n19990, ZN => n18601);
   U16247 : OAI221_X1 port map( B1 => n15407, B2 => n21031, C1 => n15269, C2 =>
                           n21036, A => n18609, ZN => n18608);
   U16248 : AOI22_X1 port map( A1 => n21056, A2 => n9825, B1 => n21089, B2 => 
                           n19991, ZN => n18609);
   U16249 : OAI221_X1 port map( B1 => n15371, B2 => n21029, C1 => n15233, C2 =>
                           n21035, A => n18564, ZN => n18563);
   U16250 : AOI22_X1 port map( A1 => n21062, A2 => n9792, B1 => n21092, B2 => 
                           n19992, ZN => n18564);
   U16251 : OAI221_X1 port map( B1 => n15406, B2 => n21028, C1 => n15268, C2 =>
                           n21032, A => n18572, ZN => n18571);
   U16252 : AOI22_X1 port map( A1 => n21062, A2 => n9824, B1 => n21091, B2 => 
                           n19993, ZN => n18572);
   U16253 : OAI221_X1 port map( B1 => n15370, B2 => n21028, C1 => n15232, C2 =>
                           n21034, A => n18527, ZN => n18526);
   U16254 : AOI22_X1 port map( A1 => n21063, A2 => n9791, B1 => n21101, B2 => 
                           n19994, ZN => n18527);
   U16255 : OAI221_X1 port map( B1 => n15405, B2 => n21027, C1 => n15267, C2 =>
                           n21033, A => n18535, ZN => n18534);
   U16256 : AOI22_X1 port map( A1 => n21062, A2 => n9823, B1 => n21100, B2 => 
                           n19995, ZN => n18535);
   U16257 : OAI221_X1 port map( B1 => n15369, B2 => n21030, C1 => n15231, C2 =>
                           n21036, A => n18464, ZN => n18461);
   U16258 : AOI22_X1 port map( A1 => n21064, A2 => n9790, B1 => n21096, B2 => 
                           n19996, ZN => n18464);
   U16259 : OAI221_X1 port map( B1 => n15404, B2 => n21029, C1 => n15266, C2 =>
                           n21035, A => n18486, ZN => n18485);
   U16260 : AOI22_X1 port map( A1 => n21064, A2 => n9822, B1 => n21096, B2 => 
                           n19997, ZN => n18486);
   U16261 : OAI221_X1 port map( B1 => n15400, B2 => n21587, C1 => n15262, C2 =>
                           n21589, A => n18380, ZN => n18379);
   U16262 : AOI22_X1 port map( A1 => n21595, A2 => n9821, B1 => n21635, B2 => 
                           n19937, ZN => n18380);
   U16263 : OAI221_X1 port map( B1 => n15435, B2 => n21586, C1 => n15297, C2 =>
                           n21594, A => n18391, ZN => n18390);
   U16264 : AOI22_X1 port map( A1 => n21625, A2 => n9853, B1 => n21634, B2 => 
                           n19938, ZN => n18391);
   U16265 : OAI221_X1 port map( B1 => n15399, B2 => n21583, C1 => n15261, C2 =>
                           n21591, A => n18319, ZN => n18318);
   U16266 : AOI22_X1 port map( A1 => n21604, A2 => n9820, B1 => n21637, B2 => 
                           n19939, ZN => n18319);
   U16267 : OAI221_X1 port map( B1 => n15434, B2 => n21588, C1 => n15296, C2 =>
                           n21590, A => n18330, ZN => n18329);
   U16268 : AOI22_X1 port map( A1 => n21603, A2 => n9852, B1 => n21636, B2 => 
                           n19940, ZN => n18330);
   U16269 : OAI221_X1 port map( B1 => n15398, B2 => n21583, C1 => n15260, C2 =>
                           n21589, A => n18272, ZN => n18271);
   U16270 : AOI22_X1 port map( A1 => n21606, A2 => n9819, B1 => n21639, B2 => 
                           n19941, ZN => n18272);
   U16271 : OAI221_X1 port map( B1 => n15433, B2 => n21588, C1 => n15295, C2 =>
                           n21592, A => n18283, ZN => n18282);
   U16272 : AOI22_X1 port map( A1 => n21605, A2 => n9851, B1 => n21638, B2 => 
                           n19942, ZN => n18283);
   U16273 : OAI221_X1 port map( B1 => n15397, B2 => n21585, C1 => n15259, C2 =>
                           n21594, A => n18225, ZN => n18224);
   U16274 : AOI22_X1 port map( A1 => n21608, A2 => n9818, B1 => n21641, B2 => 
                           n19943, ZN => n18225);
   U16275 : OAI221_X1 port map( B1 => n15432, B2 => n21584, C1 => n15294, C2 =>
                           n21593, A => n18236, ZN => n18235);
   U16276 : AOI22_X1 port map( A1 => n21607, A2 => n9850, B1 => n21640, B2 => 
                           n19944, ZN => n18236);
   U16277 : OAI221_X1 port map( B1 => n15396, B2 => n21587, C1 => n15258, C2 =>
                           n21590, A => n18178, ZN => n18177);
   U16278 : AOI22_X1 port map( A1 => n21610, A2 => n9817, B1 => n21643, B2 => 
                           n19945, ZN => n18178);
   U16279 : OAI221_X1 port map( B1 => n15431, B2 => n21586, C1 => n15293, C2 =>
                           n21589, A => n18189, ZN => n18188);
   U16280 : AOI22_X1 port map( A1 => n21609, A2 => n9849, B1 => n21642, B2 => 
                           n19946, ZN => n18189);
   U16281 : OAI221_X1 port map( B1 => n15395, B2 => n21584, C1 => n15257, C2 =>
                           n21590, A => n18131, ZN => n18130);
   U16282 : AOI22_X1 port map( A1 => n21612, A2 => n9816, B1 => n21645, B2 => 
                           n19947, ZN => n18131);
   U16283 : OAI221_X1 port map( B1 => n15430, B2 => n21583, C1 => n15292, C2 =>
                           n21591, A => n18142, ZN => n18141);
   U16284 : AOI22_X1 port map( A1 => n21611, A2 => n9848, B1 => n21644, B2 => 
                           n19948, ZN => n18142);
   U16285 : OAI221_X1 port map( B1 => n15394, B2 => n21583, C1 => n15256, C2 =>
                           n21593, A => n18084, ZN => n18083);
   U16286 : AOI22_X1 port map( A1 => n21614, A2 => n9815, B1 => n21647, B2 => 
                           n19949, ZN => n18084);
   U16287 : OAI221_X1 port map( B1 => n15429, B2 => n21588, C1 => n15291, C2 =>
                           n21592, A => n18095, ZN => n18094);
   U16288 : AOI22_X1 port map( A1 => n21613, A2 => n9847, B1 => n21646, B2 => 
                           n19950, ZN => n18095);
   U16289 : OAI221_X1 port map( B1 => n15393, B2 => n21585, C1 => n15255, C2 =>
                           n21589, A => n18037, ZN => n18036);
   U16290 : AOI22_X1 port map( A1 => n21619, A2 => n9814, B1 => n21649, B2 => 
                           n19951, ZN => n18037);
   U16291 : OAI221_X1 port map( B1 => n15428, B2 => n21584, C1 => n15290, C2 =>
                           n21594, A => n18048, ZN => n18047);
   U16292 : AOI22_X1 port map( A1 => n21619, A2 => n9846, B1 => n21648, B2 => 
                           n19952, ZN => n18048);
   U16293 : OAI221_X1 port map( B1 => n15392, B2 => n21585, C1 => n15254, C2 =>
                           n21591, A => n17990, ZN => n17989);
   U16294 : AOI22_X1 port map( A1 => n21620, A2 => n9813, B1 => n21649, B2 => 
                           n19953, ZN => n17990);
   U16295 : OAI221_X1 port map( B1 => n15427, B2 => n21584, C1 => n15289, C2 =>
                           n21590, A => n18001, ZN => n18000);
   U16296 : AOI22_X1 port map( A1 => n21619, A2 => n9845, B1 => n21658, B2 => 
                           n19954, ZN => n18001);
   U16297 : OAI221_X1 port map( B1 => n15391, B2 => n21587, C1 => n15253, C2 =>
                           n21592, A => n17943, ZN => n17942);
   U16298 : AOI22_X1 port map( A1 => n21621, A2 => n9812, B1 => n21653, B2 => 
                           n19955, ZN => n17943);
   U16299 : OAI221_X1 port map( B1 => n15426, B2 => n21586, C1 => n15288, C2 =>
                           n21591, A => n17954, ZN => n17953);
   U16300 : AOI22_X1 port map( A1 => n21620, A2 => n9844, B1 => n21653, B2 => 
                           n19956, ZN => n17954);
   U16301 : OAI221_X1 port map( B1 => n15390, B2 => n21583, C1 => n15252, C2 =>
                           n21594, A => n17896, ZN => n17895);
   U16302 : AOI22_X1 port map( A1 => n21622, A2 => n9811, B1 => n21654, B2 => 
                           n19957, ZN => n17896);
   U16303 : OAI221_X1 port map( B1 => n15425, B2 => n21588, C1 => n15287, C2 =>
                           n21593, A => n17907, ZN => n17906);
   U16304 : AOI22_X1 port map( A1 => n21623, A2 => n9843, B1 => n21653, B2 => 
                           n19958, ZN => n17907);
   U16305 : OAI221_X1 port map( B1 => n15389, B2 => n21586, C1 => n15251, C2 =>
                           n21592, A => n17849, ZN => n17848);
   U16306 : AOI22_X1 port map( A1 => n21624, A2 => n9810, B1 => n21655, B2 => 
                           n19959, ZN => n17849);
   U16307 : OAI221_X1 port map( B1 => n15424, B2 => n21585, C1 => n15286, C2 =>
                           n21589, A => n17860, ZN => n17859);
   U16308 : AOI22_X1 port map( A1 => n21623, A2 => n9842, B1 => n21654, B2 => 
                           n19960, ZN => n17860);
   U16309 : OAI221_X1 port map( B1 => n15388, B2 => n21585, C1 => n15250, C2 =>
                           n21591, A => n17802, ZN => n17801);
   U16310 : AOI22_X1 port map( A1 => n21625, A2 => n9809, B1 => n21656, B2 => 
                           n19961, ZN => n17802);
   U16311 : OAI221_X1 port map( B1 => n15423, B2 => n21584, C1 => n15285, C2 =>
                           n21590, A => n17813, ZN => n17812);
   U16312 : AOI22_X1 port map( A1 => n21625, A2 => n9841, B1 => n21656, B2 => 
                           n19962, ZN => n17813);
   U16313 : OAI221_X1 port map( B1 => n15387, B2 => n21587, C1 => n15249, C2 =>
                           n21593, A => n17755, ZN => n17754);
   U16314 : AOI22_X1 port map( A1 => n21626, A2 => n9808, B1 => n21657, B2 => 
                           n19963, ZN => n17755);
   U16315 : OAI221_X1 port map( B1 => n15422, B2 => n21586, C1 => n15284, C2 =>
                           n21592, A => n17766, ZN => n17765);
   U16316 : AOI22_X1 port map( A1 => n21626, A2 => n9840, B1 => n21656, B2 => 
                           n19964, ZN => n17766);
   U16317 : OAI221_X1 port map( B1 => n15386, B2 => n21587, C1 => n15248, C2 =>
                           n21593, A => n17708, ZN => n17707);
   U16318 : AOI22_X1 port map( A1 => n21622, A2 => n9807, B1 => n21655, B2 => 
                           n19965, ZN => n17708);
   U16319 : OAI221_X1 port map( B1 => n15421, B2 => n21586, C1 => n15283, C2 =>
                           n21594, A => n17719, ZN => n17718);
   U16320 : AOI22_X1 port map( A1 => n21602, A2 => n9839, B1 => n21654, B2 => 
                           n19966, ZN => n17719);
   U16321 : OAI221_X1 port map( B1 => n15385, B2 => n21583, C1 => n15247, C2 =>
                           n21590, A => n17661, ZN => n17660);
   U16322 : AOI22_X1 port map( A1 => n21622, A2 => n9806, B1 => n21656, B2 => 
                           n19967, ZN => n17661);
   U16323 : OAI221_X1 port map( B1 => n15420, B2 => n21588, C1 => n15282, C2 =>
                           n21589, A => n17672, ZN => n17671);
   U16324 : AOI22_X1 port map( A1 => n21623, A2 => n9838, B1 => n21656, B2 => 
                           n19968, ZN => n17672);
   U16325 : OAI221_X1 port map( B1 => n15384, B2 => n21585, C1 => n15246, C2 =>
                           n21592, A => n17614, ZN => n17613);
   U16326 : AOI22_X1 port map( A1 => n21624, A2 => n9805, B1 => n21657, B2 => 
                           n19969, ZN => n17614);
   U16327 : OAI221_X1 port map( B1 => n15419, B2 => n21584, C1 => n15281, C2 =>
                           n21591, A => n17625, ZN => n17624);
   U16328 : AOI22_X1 port map( A1 => n21623, A2 => n9837, B1 => n21656, B2 => 
                           n19970, ZN => n17625);
   U16329 : OAI221_X1 port map( B1 => n15383, B2 => n21588, C1 => n15245, C2 =>
                           n21594, A => n17567, ZN => n17566);
   U16330 : AOI22_X1 port map( A1 => n21625, A2 => n9804, B1 => n21655, B2 => 
                           n19971, ZN => n17567);
   U16331 : OAI221_X1 port map( B1 => n15418, B2 => n21587, C1 => n15280, C2 =>
                           n21593, A => n17578, ZN => n17577);
   U16332 : AOI22_X1 port map( A1 => n21624, A2 => n9836, B1 => n21653, B2 => 
                           n19972, ZN => n17578);
   U16333 : OAI221_X1 port map( B1 => n15417, B2 => n21586, C1 => n15279, C2 =>
                           n21594, A => n17531, ZN => n17530);
   U16334 : AOI22_X1 port map( A1 => n21626, A2 => n9835, B1 => n21658, B2 => 
                           n19973, ZN => n17531);
   U16335 : OAI221_X1 port map( B1 => n15416, B2 => n21588, C1 => n15278, C2 =>
                           n21590, A => n17484, ZN => n17483);
   U16336 : AOI22_X1 port map( A1 => n21627, A2 => n9834, B1 => n21659, B2 => 
                           n19974, ZN => n17484);
   U16337 : OAI221_X1 port map( B1 => n15380, B2 => n21583, C1 => n15242, C2 =>
                           n21589, A => n17426, ZN => n17425);
   U16338 : AOI22_X1 port map( A1 => n21601, A2 => n9801, B1 => n21660, B2 => 
                           n19975, ZN => n17426);
   U16339 : OAI221_X1 port map( B1 => n15415, B2 => n21588, C1 => n15277, C2 =>
                           n21592, A => n17437, ZN => n17436);
   U16340 : AOI22_X1 port map( A1 => n21624, A2 => n9833, B1 => n21659, B2 => 
                           n19976, ZN => n17437);
   U16341 : OAI221_X1 port map( B1 => n15414, B2 => n21584, C1 => n15276, C2 =>
                           n21593, A => n17390, ZN => n17389);
   U16342 : AOI22_X1 port map( A1 => n21602, A2 => n9832, B1 => n21660, B2 => 
                           n19977, ZN => n17390);
   U16343 : OAI221_X1 port map( B1 => n15378, B2 => n21587, C1 => n15240, C2 =>
                           n21590, A => n17332, ZN => n17331);
   U16344 : AOI22_X1 port map( A1 => n21627, A2 => n9799, B1 => n21635, B2 => 
                           n19978, ZN => n17332);
   U16345 : OAI221_X1 port map( B1 => n15413, B2 => n21586, C1 => n15275, C2 =>
                           n21589, A => n17343, ZN => n17342);
   U16346 : AOI22_X1 port map( A1 => n21623, A2 => n9831, B1 => n21634, B2 => 
                           n19979, ZN => n17343);
   U16347 : OAI221_X1 port map( B1 => n15377, B2 => n21584, C1 => n15239, C2 =>
                           n21590, A => n17285, ZN => n17284);
   U16348 : AOI22_X1 port map( A1 => n21604, A2 => n9798, B1 => n21637, B2 => 
                           n19980, ZN => n17285);
   U16349 : OAI221_X1 port map( B1 => n15412, B2 => n21583, C1 => n15274, C2 =>
                           n21591, A => n17296, ZN => n17295);
   U16350 : AOI22_X1 port map( A1 => n21603, A2 => n9830, B1 => n21636, B2 => 
                           n19981, ZN => n17296);
   U16351 : OAI221_X1 port map( B1 => n15376, B2 => n21583, C1 => n15238, C2 =>
                           n21593, A => n17238, ZN => n17237);
   U16352 : AOI22_X1 port map( A1 => n21606, A2 => n9797, B1 => n21639, B2 => 
                           n19982, ZN => n17238);
   U16353 : OAI221_X1 port map( B1 => n15411, B2 => n21588, C1 => n15273, C2 =>
                           n21592, A => n17249, ZN => n17248);
   U16354 : AOI22_X1 port map( A1 => n21605, A2 => n9829, B1 => n21638, B2 => 
                           n19983, ZN => n17249);
   U16355 : OAI221_X1 port map( B1 => n15375, B2 => n21585, C1 => n15237, C2 =>
                           n21589, A => n17191, ZN => n17190);
   U16356 : AOI22_X1 port map( A1 => n21608, A2 => n9796, B1 => n21641, B2 => 
                           n19984, ZN => n17191);
   U16357 : OAI221_X1 port map( B1 => n15410, B2 => n21584, C1 => n15272, C2 =>
                           n21594, A => n17202, ZN => n17201);
   U16358 : AOI22_X1 port map( A1 => n21607, A2 => n9828, B1 => n21640, B2 => 
                           n19985, ZN => n17202);
   U16359 : OAI221_X1 port map( B1 => n15374, B2 => n21585, C1 => n15236, C2 =>
                           n21591, A => n17144, ZN => n17143);
   U16360 : AOI22_X1 port map( A1 => n21610, A2 => n9795, B1 => n21643, B2 => 
                           n19986, ZN => n17144);
   U16361 : OAI221_X1 port map( B1 => n15409, B2 => n21584, C1 => n15271, C2 =>
                           n21590, A => n17155, ZN => n17154);
   U16362 : AOI22_X1 port map( A1 => n21609, A2 => n9827, B1 => n21642, B2 => 
                           n19987, ZN => n17155);
   U16363 : OAI221_X1 port map( B1 => n15373, B2 => n21587, C1 => n15235, C2 =>
                           n21592, A => n17097, ZN => n17096);
   U16364 : AOI22_X1 port map( A1 => n21612, A2 => n9794, B1 => n21645, B2 => 
                           n19988, ZN => n17097);
   U16365 : OAI221_X1 port map( B1 => n15408, B2 => n21586, C1 => n15270, C2 =>
                           n21591, A => n17108, ZN => n17107);
   U16366 : AOI22_X1 port map( A1 => n21611, A2 => n9826, B1 => n21644, B2 => 
                           n19989, ZN => n17108);
   U16367 : OAI221_X1 port map( B1 => n15372, B2 => n21583, C1 => n15234, C2 =>
                           n21594, A => n17050, ZN => n17049);
   U16368 : AOI22_X1 port map( A1 => n21614, A2 => n9793, B1 => n21647, B2 => 
                           n19990, ZN => n17050);
   U16369 : OAI221_X1 port map( B1 => n15407, B2 => n21588, C1 => n15269, C2 =>
                           n21593, A => n17061, ZN => n17060);
   U16370 : AOI22_X1 port map( A1 => n21613, A2 => n9825, B1 => n21646, B2 => 
                           n19991, ZN => n17061);
   U16371 : OAI221_X1 port map( B1 => n15371, B2 => n21586, C1 => n15233, C2 =>
                           n21592, A => n17003, ZN => n17002);
   U16372 : AOI22_X1 port map( A1 => n21619, A2 => n9792, B1 => n21649, B2 => 
                           n19992, ZN => n17003);
   U16373 : OAI221_X1 port map( B1 => n15406, B2 => n21585, C1 => n15268, C2 =>
                           n21589, A => n17014, ZN => n17013);
   U16374 : AOI22_X1 port map( A1 => n21619, A2 => n9824, B1 => n21648, B2 => 
                           n19993, ZN => n17014);
   U16375 : OAI221_X1 port map( B1 => n15370, B2 => n21585, C1 => n15232, C2 =>
                           n21591, A => n16956, ZN => n16955);
   U16376 : AOI22_X1 port map( A1 => n21620, A2 => n9791, B1 => n21658, B2 => 
                           n19994, ZN => n16956);
   U16377 : OAI221_X1 port map( B1 => n15405, B2 => n21584, C1 => n15267, C2 =>
                           n21590, A => n16967, ZN => n16966);
   U16378 : AOI22_X1 port map( A1 => n21619, A2 => n9823, B1 => n21657, B2 => 
                           n19995, ZN => n16967);
   U16379 : OAI221_X1 port map( B1 => n15369, B2 => n21587, C1 => n15231, C2 =>
                           n21593, A => n16883, ZN => n16880);
   U16380 : AOI22_X1 port map( A1 => n21621, A2 => n9790, B1 => n21653, B2 => 
                           n19996, ZN => n16883);
   U16381 : OAI221_X1 port map( B1 => n15404, B2 => n21586, C1 => n15266, C2 =>
                           n21592, A => n16908, ZN => n16907);
   U16382 : AOI22_X1 port map( A1 => n21621, A2 => n9822, B1 => n21653, B2 => 
                           n19997, ZN => n16908);
   U16383 : OAI221_X1 port map( B1 => n15679, B2 => n20985, C1 => n15785, C2 =>
                           n20987, A => n19652, ZN => n19649);
   U16384 : AOI22_X1 port map( A1 => n21000, A2 => n19813, B1 => n20696, B2 => 
                           n8921, ZN => n19652);
   U16385 : OAI221_X1 port map( B1 => n15714, B2 => n20984, C1 => n15820, C2 =>
                           n20992, A => n19664, ZN => n19657);
   U16386 : AOI22_X1 port map( A1 => n20999, A2 => n19814, B1 => n20695, B2 => 
                           n8925, ZN => n19664);
   U16387 : OAI221_X1 port map( B1 => n15678, B2 => n20981, C1 => n15784, C2 =>
                           n20989, A => n19601, ZN => n19598);
   U16388 : AOI22_X1 port map( A1 => n21002, A2 => n19815, B1 => n20698, B2 => 
                           n8910, ZN => n19601);
   U16389 : OAI221_X1 port map( B1 => n15713, B2 => n20986, C1 => n15819, C2 =>
                           n20988, A => n19609, ZN => n19606);
   U16390 : AOI22_X1 port map( A1 => n21001, A2 => n19816, B1 => n20697, B2 => 
                           n8914, ZN => n19609);
   U16391 : OAI221_X1 port map( B1 => n15677, B2 => n20981, C1 => n15783, C2 =>
                           n20987, A => n19564, ZN => n19561);
   U16392 : AOI22_X1 port map( A1 => n21004, A2 => n19817, B1 => n20700, B2 => 
                           n8899, ZN => n19564);
   U16393 : OAI221_X1 port map( B1 => n15712, B2 => n20986, C1 => n15818, C2 =>
                           n20990, A => n19572, ZN => n19569);
   U16394 : AOI22_X1 port map( A1 => n21003, A2 => n19818, B1 => n20699, B2 => 
                           n8903, ZN => n19572);
   U16395 : OAI221_X1 port map( B1 => n15676, B2 => n20983, C1 => n15782, C2 =>
                           n20992, A => n19527, ZN => n19524);
   U16396 : AOI22_X1 port map( A1 => n21006, A2 => n19819, B1 => n20702, B2 => 
                           n8888, ZN => n19527);
   U16397 : OAI221_X1 port map( B1 => n15711, B2 => n20982, C1 => n15817, C2 =>
                           n20991, A => n19535, ZN => n19532);
   U16398 : AOI22_X1 port map( A1 => n21005, A2 => n19820, B1 => n20701, B2 => 
                           n8892, ZN => n19535);
   U16399 : OAI221_X1 port map( B1 => n15675, B2 => n20985, C1 => n15781, C2 =>
                           n20988, A => n19490, ZN => n19487);
   U16400 : AOI22_X1 port map( A1 => n21008, A2 => n19821, B1 => n20704, B2 => 
                           n8877, ZN => n19490);
   U16401 : OAI221_X1 port map( B1 => n15710, B2 => n20984, C1 => n15816, C2 =>
                           n20987, A => n19498, ZN => n19495);
   U16402 : AOI22_X1 port map( A1 => n21007, A2 => n19822, B1 => n20703, B2 => 
                           n8881, ZN => n19498);
   U16403 : OAI221_X1 port map( B1 => n15674, B2 => n20982, C1 => n15780, C2 =>
                           n20988, A => n19453, ZN => n19450);
   U16404 : AOI22_X1 port map( A1 => n21010, A2 => n19823, B1 => n20706, B2 => 
                           n8866, ZN => n19453);
   U16405 : OAI221_X1 port map( B1 => n15709, B2 => n20981, C1 => n15815, C2 =>
                           n20989, A => n19461, ZN => n19458);
   U16406 : AOI22_X1 port map( A1 => n21009, A2 => n19824, B1 => n20705, B2 => 
                           n8870, ZN => n19461);
   U16407 : OAI221_X1 port map( B1 => n15673, B2 => n20981, C1 => n15779, C2 =>
                           n20991, A => n19416, ZN => n19413);
   U16408 : AOI22_X1 port map( A1 => n21012, A2 => n19825, B1 => n20708, B2 => 
                           n8855, ZN => n19416);
   U16409 : OAI221_X1 port map( B1 => n15708, B2 => n20986, C1 => n15814, C2 =>
                           n20990, A => n19424, ZN => n19421);
   U16410 : AOI22_X1 port map( A1 => n21011, A2 => n19826, B1 => n20707, B2 => 
                           n8859, ZN => n19424);
   U16411 : OAI221_X1 port map( B1 => n15672, B2 => n20983, C1 => n15778, C2 =>
                           n20987, A => n19379, ZN => n19376);
   U16412 : AOI22_X1 port map( A1 => n21012, A2 => n19827, B1 => n20708, B2 => 
                           n8844, ZN => n19379);
   U16413 : OAI221_X1 port map( B1 => n15707, B2 => n20982, C1 => n15813, C2 =>
                           n20992, A => n19387, ZN => n19384);
   U16414 : AOI22_X1 port map( A1 => n21021, A2 => n19828, B1 => n20719, B2 => 
                           n8848, ZN => n19387);
   U16415 : OAI221_X1 port map( B1 => n15671, B2 => n20983, C1 => n15777, C2 =>
                           n20989, A => n19342, ZN => n19339);
   U16416 : AOI22_X1 port map( A1 => n21018, A2 => n19829, B1 => n20712, B2 => 
                           n8833, ZN => n19342);
   U16417 : OAI221_X1 port map( B1 => n15706, B2 => n20982, C1 => n15812, C2 =>
                           n20988, A => n19350, ZN => n19347);
   U16418 : AOI22_X1 port map( A1 => n21017, A2 => n19830, B1 => n20712, B2 => 
                           n8837, ZN => n19350);
   U16419 : OAI221_X1 port map( B1 => n15670, B2 => n20985, C1 => n15776, C2 =>
                           n20990, A => n19305, ZN => n19302);
   U16420 : AOI22_X1 port map( A1 => n21019, A2 => n19831, B1 => n20713, B2 => 
                           n8822, ZN => n19305);
   U16421 : OAI221_X1 port map( B1 => n15705, B2 => n20984, C1 => n15811, C2 =>
                           n20989, A => n19313, ZN => n19310);
   U16422 : AOI22_X1 port map( A1 => n21017, A2 => n19832, B1 => n20712, B2 => 
                           n8826, ZN => n19313);
   U16423 : OAI221_X1 port map( B1 => n15669, B2 => n20981, C1 => n15775, C2 =>
                           n20992, A => n19268, ZN => n19265);
   U16424 : AOI22_X1 port map( A1 => n21020, A2 => n19833, B1 => n20714, B2 => 
                           n8811, ZN => n19268);
   U16425 : OAI221_X1 port map( B1 => n15704, B2 => n20986, C1 => n15810, C2 =>
                           n20991, A => n19276, ZN => n19273);
   U16426 : AOI22_X1 port map( A1 => n21019, A2 => n19834, B1 => n20713, B2 => 
                           n8815, ZN => n19276);
   U16427 : OAI221_X1 port map( B1 => n15668, B2 => n20984, C1 => n15774, C2 =>
                           n20990, A => n19231, ZN => n19228);
   U16428 : AOI22_X1 port map( A1 => n21021, A2 => n19835, B1 => n20715, B2 => 
                           n8800, ZN => n19231);
   U16429 : OAI221_X1 port map( B1 => n15703, B2 => n20983, C1 => n15809, C2 =>
                           n20987, A => n19239, ZN => n19236);
   U16430 : AOI22_X1 port map( A1 => n21022, A2 => n19836, B1 => n20715, B2 => 
                           n8804, ZN => n19239);
   U16431 : OAI221_X1 port map( B1 => n15667, B2 => n20983, C1 => n15773, C2 =>
                           n20989, A => n19194, ZN => n19191);
   U16432 : AOI22_X1 port map( A1 => n21023, A2 => n19837, B1 => n20716, B2 => 
                           n8789, ZN => n19194);
   U16433 : OAI221_X1 port map( B1 => n15702, B2 => n20982, C1 => n15808, C2 =>
                           n20988, A => n19202, ZN => n19199);
   U16434 : AOI22_X1 port map( A1 => n21022, A2 => n19838, B1 => n20715, B2 => 
                           n8793, ZN => n19202);
   U16435 : OAI221_X1 port map( B1 => n15666, B2 => n20985, C1 => n15772, C2 =>
                           n20991, A => n19157, ZN => n19154);
   U16436 : AOI22_X1 port map( A1 => n21018, A2 => n19839, B1 => n20717, B2 => 
                           n8778, ZN => n19157);
   U16437 : OAI221_X1 port map( B1 => n15701, B2 => n20984, C1 => n15807, C2 =>
                           n20990, A => n19165, ZN => n19162);
   U16438 : AOI22_X1 port map( A1 => n21023, A2 => n19840, B1 => n20717, B2 => 
                           n8782, ZN => n19165);
   U16439 : OAI221_X1 port map( B1 => n15665, B2 => n20985, C1 => n15771, C2 =>
                           n20991, A => n19120, ZN => n19117);
   U16440 : AOI22_X1 port map( A1 => n21020, A2 => n19841, B1 => n20714, B2 => 
                           n8767, ZN => n19120);
   U16441 : OAI221_X1 port map( B1 => n15700, B2 => n20984, C1 => n15806, C2 =>
                           n20992, A => n19128, ZN => n19125);
   U16442 : AOI22_X1 port map( A1 => n20999, A2 => n19842, B1 => n20694, B2 => 
                           n8771, ZN => n19128);
   U16443 : OAI221_X1 port map( B1 => n15664, B2 => n20981, C1 => n15770, C2 =>
                           n20988, A => n19083, ZN => n19080);
   U16444 : AOI22_X1 port map( A1 => n21021, A2 => n19843, B1 => n20715, B2 => 
                           n8756, ZN => n19083);
   U16445 : OAI221_X1 port map( B1 => n15699, B2 => n20986, C1 => n15805, C2 =>
                           n20987, A => n19091, ZN => n19088);
   U16446 : AOI22_X1 port map( A1 => n21022, A2 => n19844, B1 => n20715, B2 => 
                           n8760, ZN => n19091);
   U16447 : OAI221_X1 port map( B1 => n15663, B2 => n20983, C1 => n15769, C2 =>
                           n20990, A => n19046, ZN => n19043);
   U16448 : AOI22_X1 port map( A1 => n21023, A2 => n19845, B1 => n20716, B2 => 
                           n8745, ZN => n19046);
   U16449 : OAI221_X1 port map( B1 => n15698, B2 => n20982, C1 => n15804, C2 =>
                           n20989, A => n19054, ZN => n19051);
   U16450 : AOI22_X1 port map( A1 => n21022, A2 => n19846, B1 => n20715, B2 => 
                           n8749, ZN => n19054);
   U16451 : OAI221_X1 port map( B1 => n15662, B2 => n20986, C1 => n15768, C2 =>
                           n20992, A => n19009, ZN => n19006);
   U16452 : AOI22_X1 port map( A1 => n21020, A2 => n19847, B1 => n20713, B2 => 
                           n8734, ZN => n19009);
   U16453 : OAI221_X1 port map( B1 => n15697, B2 => n20985, C1 => n15803, C2 =>
                           n20991, A => n19017, ZN => n19014);
   U16454 : AOI22_X1 port map( A1 => n21023, A2 => n19848, B1 => n20717, B2 => 
                           n8738, ZN => n19017);
   U16455 : OAI221_X1 port map( B1 => n15661, B2 => n20985, C1 => n15767, C2 =>
                           n20987, A => n18972, ZN => n18969);
   U16456 : AOI22_X1 port map( A1 => n21024, A2 => n19849, B1 => n20718, B2 => 
                           n8723, ZN => n18972);
   U16457 : OAI221_X1 port map( B1 => n15696, B2 => n20984, C1 => n15802, C2 =>
                           n20992, A => n18980, ZN => n18977);
   U16458 : AOI22_X1 port map( A1 => n21024, A2 => n19850, B1 => n20718, B2 => 
                           n8727, ZN => n18980);
   U16459 : OAI221_X1 port map( B1 => n15660, B2 => n20981, C1 => n15766, C2 =>
                           n20989, A => n18935, ZN => n18932);
   U16460 : AOI22_X1 port map( A1 => n21025, A2 => n19851, B1 => n20719, B2 => 
                           n8712, ZN => n18935);
   U16461 : OAI221_X1 port map( B1 => n15695, B2 => n20986, C1 => n15801, C2 =>
                           n20988, A => n18943, ZN => n18940);
   U16462 : AOI22_X1 port map( A1 => n21024, A2 => n19852, B1 => n20718, B2 => 
                           n8716, ZN => n18943);
   U16463 : OAI221_X1 port map( B1 => n15694, B2 => n20986, C1 => n15800, C2 =>
                           n20990, A => n18906, ZN => n18903);
   U16464 : AOI22_X1 port map( A1 => n21025, A2 => n19680, B1 => n20719, B2 => 
                           n8705, ZN => n18906);
   U16465 : OAI221_X1 port map( B1 => n15658, B2 => n20983, C1 => n15764, C2 =>
                           n20992, A => n18861, ZN => n18858);
   U16466 : AOI22_X1 port map( A1 => n20999, A2 => n19853, B1 => n20694, B2 => 
                           n8690, ZN => n18861);
   U16467 : OAI221_X1 port map( B1 => n15693, B2 => n20982, C1 => n15799, C2 =>
                           n20991, A => n18869, ZN => n18866);
   U16468 : AOI22_X1 port map( A1 => n21022, A2 => n19854, B1 => n20693, B2 => 
                           n8694, ZN => n18869);
   U16469 : OAI221_X1 port map( B1 => n15657, B2 => n20985, C1 => n15763, C2 =>
                           n20988, A => n18824, ZN => n18821);
   U16470 : AOI22_X1 port map( A1 => n21000, A2 => n19855, B1 => n20696, B2 => 
                           n8679, ZN => n18824);
   U16471 : OAI221_X1 port map( B1 => n15692, B2 => n20984, C1 => n15798, C2 =>
                           n20987, A => n18832, ZN => n18829);
   U16472 : AOI22_X1 port map( A1 => n21025, A2 => n19856, B1 => n20695, B2 => 
                           n8683, ZN => n18832);
   U16473 : OAI221_X1 port map( B1 => n15656, B2 => n20982, C1 => n15762, C2 =>
                           n20988, A => n18787, ZN => n18784);
   U16474 : AOI22_X1 port map( A1 => n21002, A2 => n19857, B1 => n20698, B2 => 
                           n8668, ZN => n18787);
   U16475 : OAI221_X1 port map( B1 => n15691, B2 => n20981, C1 => n15797, C2 =>
                           n20989, A => n18795, ZN => n18792);
   U16476 : AOI22_X1 port map( A1 => n21001, A2 => n19858, B1 => n20697, B2 => 
                           n8672, ZN => n18795);
   U16477 : OAI221_X1 port map( B1 => n15655, B2 => n20981, C1 => n15761, C2 =>
                           n20991, A => n18750, ZN => n18747);
   U16478 : AOI22_X1 port map( A1 => n21004, A2 => n19859, B1 => n20700, B2 => 
                           n8657, ZN => n18750);
   U16479 : OAI221_X1 port map( B1 => n15690, B2 => n20986, C1 => n15796, C2 =>
                           n20990, A => n18758, ZN => n18755);
   U16480 : AOI22_X1 port map( A1 => n21003, A2 => n19860, B1 => n20699, B2 => 
                           n8661, ZN => n18758);
   U16481 : OAI221_X1 port map( B1 => n15654, B2 => n20983, C1 => n15760, C2 =>
                           n20987, A => n18713, ZN => n18710);
   U16482 : AOI22_X1 port map( A1 => n21006, A2 => n19861, B1 => n20702, B2 => 
                           n8646, ZN => n18713);
   U16483 : OAI221_X1 port map( B1 => n15689, B2 => n20982, C1 => n15795, C2 =>
                           n20992, A => n18721, ZN => n18718);
   U16484 : AOI22_X1 port map( A1 => n21005, A2 => n19862, B1 => n20701, B2 => 
                           n8650, ZN => n18721);
   U16485 : OAI221_X1 port map( B1 => n15653, B2 => n20983, C1 => n15759, C2 =>
                           n20989, A => n18676, ZN => n18673);
   U16486 : AOI22_X1 port map( A1 => n21008, A2 => n19863, B1 => n20704, B2 => 
                           n8635, ZN => n18676);
   U16487 : OAI221_X1 port map( B1 => n15688, B2 => n20982, C1 => n15794, C2 =>
                           n20988, A => n18684, ZN => n18681);
   U16488 : AOI22_X1 port map( A1 => n21007, A2 => n19864, B1 => n20703, B2 => 
                           n8639, ZN => n18684);
   U16489 : OAI221_X1 port map( B1 => n15652, B2 => n20985, C1 => n15758, C2 =>
                           n20990, A => n18639, ZN => n18636);
   U16490 : AOI22_X1 port map( A1 => n21010, A2 => n19865, B1 => n20706, B2 => 
                           n8624, ZN => n18639);
   U16491 : OAI221_X1 port map( B1 => n15687, B2 => n20984, C1 => n15793, C2 =>
                           n20989, A => n18647, ZN => n18644);
   U16492 : AOI22_X1 port map( A1 => n21009, A2 => n19866, B1 => n20705, B2 => 
                           n8628, ZN => n18647);
   U16493 : OAI221_X1 port map( B1 => n15651, B2 => n20981, C1 => n15757, C2 =>
                           n20992, A => n18602, ZN => n18599);
   U16494 : AOI22_X1 port map( A1 => n21012, A2 => n19867, B1 => n20708, B2 => 
                           n8613, ZN => n18602);
   U16495 : OAI221_X1 port map( B1 => n15686, B2 => n20986, C1 => n15792, C2 =>
                           n20991, A => n18610, ZN => n18607);
   U16496 : AOI22_X1 port map( A1 => n21011, A2 => n19868, B1 => n20707, B2 => 
                           n8617, ZN => n18610);
   U16497 : OAI221_X1 port map( B1 => n15650, B2 => n20984, C1 => n15756, C2 =>
                           n20990, A => n18565, ZN => n18562);
   U16498 : AOI22_X1 port map( A1 => n21024, A2 => n19869, B1 => n20718, B2 => 
                           n8602, ZN => n18565);
   U16499 : OAI221_X1 port map( B1 => n15685, B2 => n20983, C1 => n15791, C2 =>
                           n20987, A => n18573, ZN => n18570);
   U16500 : AOI22_X1 port map( A1 => n21021, A2 => n19870, B1 => n20718, B2 => 
                           n8606, ZN => n18573);
   U16501 : OAI221_X1 port map( B1 => n15649, B2 => n20983, C1 => n15755, C2 =>
                           n20989, A => n18528, ZN => n18525);
   U16502 : AOI22_X1 port map( A1 => n21018, A2 => n19871, B1 => n20712, B2 => 
                           n8591, ZN => n18528);
   U16503 : OAI221_X1 port map( B1 => n15684, B2 => n20982, C1 => n15790, C2 =>
                           n20988, A => n18536, ZN => n18533);
   U16504 : AOI22_X1 port map( A1 => n21017, A2 => n19872, B1 => n20712, B2 => 
                           n8595, ZN => n18536);
   U16505 : OAI221_X1 port map( B1 => n15648, B2 => n20985, C1 => n15754, C2 =>
                           n20991, A => n18469, ZN => n18460);
   U16506 : AOI22_X1 port map( A1 => n21019, A2 => n19873, B1 => n20714, B2 => 
                           n8580, ZN => n18469);
   U16507 : OAI221_X1 port map( B1 => n15683, B2 => n20984, C1 => n15789, C2 =>
                           n20990, A => n18487, ZN => n18484);
   U16508 : AOI22_X1 port map( A1 => n21017, A2 => n19874, B1 => n20712, B2 => 
                           n8584, ZN => n18487);
   U16509 : OAI221_X1 port map( B1 => n15679, B2 => n21542, C1 => n15785, C2 =>
                           n21544, A => n18382, ZN => n18378);
   U16510 : AOI22_X1 port map( A1 => n21557, A2 => n19813, B1 => n21253, B2 => 
                           n8921, ZN => n18382);
   U16511 : OAI221_X1 port map( B1 => n15714, B2 => n21541, C1 => n15820, C2 =>
                           n21549, A => n18397, ZN => n18389);
   U16512 : AOI22_X1 port map( A1 => n21556, A2 => n19814, B1 => n21252, B2 => 
                           n8925, ZN => n18397);
   U16513 : OAI221_X1 port map( B1 => n15678, B2 => n21538, C1 => n15784, C2 =>
                           n21546, A => n18321, ZN => n18317);
   U16514 : AOI22_X1 port map( A1 => n21559, A2 => n19815, B1 => n21255, B2 => 
                           n8910, ZN => n18321);
   U16515 : OAI221_X1 port map( B1 => n15713, B2 => n21543, C1 => n15819, C2 =>
                           n21545, A => n18332, ZN => n18328);
   U16516 : AOI22_X1 port map( A1 => n21558, A2 => n19816, B1 => n21254, B2 => 
                           n8914, ZN => n18332);
   U16517 : OAI221_X1 port map( B1 => n15677, B2 => n21538, C1 => n15783, C2 =>
                           n21544, A => n18274, ZN => n18270);
   U16518 : AOI22_X1 port map( A1 => n21561, A2 => n19817, B1 => n21257, B2 => 
                           n8899, ZN => n18274);
   U16519 : OAI221_X1 port map( B1 => n15712, B2 => n21543, C1 => n15818, C2 =>
                           n21547, A => n18285, ZN => n18281);
   U16520 : AOI22_X1 port map( A1 => n21560, A2 => n19818, B1 => n21256, B2 => 
                           n8903, ZN => n18285);
   U16521 : OAI221_X1 port map( B1 => n15676, B2 => n21540, C1 => n15782, C2 =>
                           n21549, A => n18227, ZN => n18223);
   U16522 : AOI22_X1 port map( A1 => n21563, A2 => n19819, B1 => n21259, B2 => 
                           n8888, ZN => n18227);
   U16523 : OAI221_X1 port map( B1 => n15711, B2 => n21539, C1 => n15817, C2 =>
                           n21548, A => n18238, ZN => n18234);
   U16524 : AOI22_X1 port map( A1 => n21562, A2 => n19820, B1 => n21258, B2 => 
                           n8892, ZN => n18238);
   U16525 : OAI221_X1 port map( B1 => n15675, B2 => n21542, C1 => n15781, C2 =>
                           n21545, A => n18180, ZN => n18176);
   U16526 : AOI22_X1 port map( A1 => n21565, A2 => n19821, B1 => n21261, B2 => 
                           n8877, ZN => n18180);
   U16527 : OAI221_X1 port map( B1 => n15710, B2 => n21541, C1 => n15816, C2 =>
                           n21544, A => n18191, ZN => n18187);
   U16528 : AOI22_X1 port map( A1 => n21564, A2 => n19822, B1 => n21260, B2 => 
                           n8881, ZN => n18191);
   U16529 : OAI221_X1 port map( B1 => n15674, B2 => n21539, C1 => n15780, C2 =>
                           n21545, A => n18133, ZN => n18129);
   U16530 : AOI22_X1 port map( A1 => n21567, A2 => n19823, B1 => n21263, B2 => 
                           n8866, ZN => n18133);
   U16531 : OAI221_X1 port map( B1 => n15709, B2 => n21538, C1 => n15815, C2 =>
                           n21546, A => n18144, ZN => n18140);
   U16532 : AOI22_X1 port map( A1 => n21566, A2 => n19824, B1 => n21262, B2 => 
                           n8870, ZN => n18144);
   U16533 : OAI221_X1 port map( B1 => n15673, B2 => n21538, C1 => n15779, C2 =>
                           n21548, A => n18086, ZN => n18082);
   U16534 : AOI22_X1 port map( A1 => n21569, A2 => n19825, B1 => n21265, B2 => 
                           n8855, ZN => n18086);
   U16535 : OAI221_X1 port map( B1 => n15708, B2 => n21543, C1 => n15814, C2 =>
                           n21547, A => n18097, ZN => n18093);
   U16536 : AOI22_X1 port map( A1 => n21568, A2 => n19826, B1 => n21264, B2 => 
                           n8859, ZN => n18097);
   U16537 : OAI221_X1 port map( B1 => n15672, B2 => n21540, C1 => n15778, C2 =>
                           n21544, A => n18039, ZN => n18035);
   U16538 : AOI22_X1 port map( A1 => n21569, A2 => n19827, B1 => n21265, B2 => 
                           n8844, ZN => n18039);
   U16539 : OAI221_X1 port map( B1 => n15707, B2 => n21539, C1 => n15813, C2 =>
                           n21549, A => n18050, ZN => n18046);
   U16540 : AOI22_X1 port map( A1 => n21578, A2 => n19828, B1 => n21276, B2 => 
                           n8848, ZN => n18050);
   U16541 : OAI221_X1 port map( B1 => n15671, B2 => n21540, C1 => n15777, C2 =>
                           n21546, A => n17992, ZN => n17988);
   U16542 : AOI22_X1 port map( A1 => n21575, A2 => n19829, B1 => n21269, B2 => 
                           n8833, ZN => n17992);
   U16543 : OAI221_X1 port map( B1 => n15706, B2 => n21539, C1 => n15812, C2 =>
                           n21545, A => n18003, ZN => n17999);
   U16544 : AOI22_X1 port map( A1 => n21574, A2 => n19830, B1 => n21269, B2 => 
                           n8837, ZN => n18003);
   U16545 : OAI221_X1 port map( B1 => n15670, B2 => n21542, C1 => n15776, C2 =>
                           n21547, A => n17945, ZN => n17941);
   U16546 : AOI22_X1 port map( A1 => n21576, A2 => n19831, B1 => n21270, B2 => 
                           n8822, ZN => n17945);
   U16547 : OAI221_X1 port map( B1 => n15705, B2 => n21541, C1 => n15811, C2 =>
                           n21546, A => n17956, ZN => n17952);
   U16548 : AOI22_X1 port map( A1 => n21574, A2 => n19832, B1 => n21269, B2 => 
                           n8826, ZN => n17956);
   U16549 : OAI221_X1 port map( B1 => n15669, B2 => n21538, C1 => n15775, C2 =>
                           n21549, A => n17898, ZN => n17894);
   U16550 : AOI22_X1 port map( A1 => n21577, A2 => n19833, B1 => n21271, B2 => 
                           n8811, ZN => n17898);
   U16551 : OAI221_X1 port map( B1 => n15704, B2 => n21543, C1 => n15810, C2 =>
                           n21548, A => n17909, ZN => n17905);
   U16552 : AOI22_X1 port map( A1 => n21576, A2 => n19834, B1 => n21270, B2 => 
                           n8815, ZN => n17909);
   U16553 : OAI221_X1 port map( B1 => n15668, B2 => n21541, C1 => n15774, C2 =>
                           n21547, A => n17851, ZN => n17847);
   U16554 : AOI22_X1 port map( A1 => n21578, A2 => n19835, B1 => n21272, B2 => 
                           n8800, ZN => n17851);
   U16555 : OAI221_X1 port map( B1 => n15703, B2 => n21540, C1 => n15809, C2 =>
                           n21544, A => n17862, ZN => n17858);
   U16556 : AOI22_X1 port map( A1 => n21579, A2 => n19836, B1 => n21272, B2 => 
                           n8804, ZN => n17862);
   U16557 : OAI221_X1 port map( B1 => n15667, B2 => n21540, C1 => n15773, C2 =>
                           n21546, A => n17804, ZN => n17800);
   U16558 : AOI22_X1 port map( A1 => n21580, A2 => n19837, B1 => n21273, B2 => 
                           n8789, ZN => n17804);
   U16559 : OAI221_X1 port map( B1 => n15702, B2 => n21539, C1 => n15808, C2 =>
                           n21545, A => n17815, ZN => n17811);
   U16560 : AOI22_X1 port map( A1 => n21579, A2 => n19838, B1 => n21272, B2 => 
                           n8793, ZN => n17815);
   U16561 : OAI221_X1 port map( B1 => n15666, B2 => n21542, C1 => n15772, C2 =>
                           n21548, A => n17757, ZN => n17753);
   U16562 : AOI22_X1 port map( A1 => n21575, A2 => n19839, B1 => n21274, B2 => 
                           n8778, ZN => n17757);
   U16563 : OAI221_X1 port map( B1 => n15701, B2 => n21541, C1 => n15807, C2 =>
                           n21547, A => n17768, ZN => n17764);
   U16564 : AOI22_X1 port map( A1 => n21580, A2 => n19840, B1 => n21274, B2 => 
                           n8782, ZN => n17768);
   U16565 : OAI221_X1 port map( B1 => n15665, B2 => n21542, C1 => n15771, C2 =>
                           n21548, A => n17710, ZN => n17706);
   U16566 : AOI22_X1 port map( A1 => n21577, A2 => n19841, B1 => n21271, B2 => 
                           n8767, ZN => n17710);
   U16567 : OAI221_X1 port map( B1 => n15700, B2 => n21541, C1 => n15806, C2 =>
                           n21549, A => n17721, ZN => n17717);
   U16568 : AOI22_X1 port map( A1 => n21556, A2 => n19842, B1 => n21251, B2 => 
                           n8771, ZN => n17721);
   U16569 : OAI221_X1 port map( B1 => n15664, B2 => n21538, C1 => n15770, C2 =>
                           n21545, A => n17663, ZN => n17659);
   U16570 : AOI22_X1 port map( A1 => n21578, A2 => n19843, B1 => n21272, B2 => 
                           n8756, ZN => n17663);
   U16571 : OAI221_X1 port map( B1 => n15699, B2 => n21543, C1 => n15805, C2 =>
                           n21544, A => n17674, ZN => n17670);
   U16572 : AOI22_X1 port map( A1 => n21579, A2 => n19844, B1 => n21272, B2 => 
                           n8760, ZN => n17674);
   U16573 : OAI221_X1 port map( B1 => n15663, B2 => n21540, C1 => n15769, C2 =>
                           n21547, A => n17616, ZN => n17612);
   U16574 : AOI22_X1 port map( A1 => n21580, A2 => n19845, B1 => n21273, B2 => 
                           n8745, ZN => n17616);
   U16575 : OAI221_X1 port map( B1 => n15698, B2 => n21539, C1 => n15804, C2 =>
                           n21546, A => n17627, ZN => n17623);
   U16576 : AOI22_X1 port map( A1 => n21579, A2 => n19846, B1 => n21272, B2 => 
                           n8749, ZN => n17627);
   U16577 : OAI221_X1 port map( B1 => n15662, B2 => n21543, C1 => n15768, C2 =>
                           n21549, A => n17569, ZN => n17565);
   U16578 : AOI22_X1 port map( A1 => n21577, A2 => n19847, B1 => n21270, B2 => 
                           n8734, ZN => n17569);
   U16579 : OAI221_X1 port map( B1 => n15697, B2 => n21542, C1 => n15803, C2 =>
                           n21548, A => n17580, ZN => n17576);
   U16580 : AOI22_X1 port map( A1 => n21580, A2 => n19848, B1 => n21274, B2 => 
                           n8738, ZN => n17580);
   U16581 : OAI221_X1 port map( B1 => n15661, B2 => n21542, C1 => n15767, C2 =>
                           n21544, A => n17522, ZN => n17518);
   U16582 : AOI22_X1 port map( A1 => n21581, A2 => n19849, B1 => n21275, B2 => 
                           n8723, ZN => n17522);
   U16583 : OAI221_X1 port map( B1 => n15696, B2 => n21541, C1 => n15802, C2 =>
                           n21549, A => n17533, ZN => n17529);
   U16584 : AOI22_X1 port map( A1 => n21581, A2 => n19850, B1 => n21275, B2 => 
                           n8727, ZN => n17533);
   U16585 : OAI221_X1 port map( B1 => n15660, B2 => n21538, C1 => n15766, C2 =>
                           n21546, A => n17475, ZN => n17471);
   U16586 : AOI22_X1 port map( A1 => n21582, A2 => n19851, B1 => n21276, B2 => 
                           n8712, ZN => n17475);
   U16587 : OAI221_X1 port map( B1 => n15695, B2 => n21543, C1 => n15801, C2 =>
                           n21545, A => n17486, ZN => n17482);
   U16588 : AOI22_X1 port map( A1 => n21581, A2 => n19852, B1 => n21275, B2 => 
                           n8716, ZN => n17486);
   U16589 : OAI221_X1 port map( B1 => n15694, B2 => n21543, C1 => n15800, C2 =>
                           n21547, A => n17439, ZN => n17435);
   U16590 : AOI22_X1 port map( A1 => n21582, A2 => n19680, B1 => n21276, B2 => 
                           n8705, ZN => n17439);
   U16591 : OAI221_X1 port map( B1 => n15658, B2 => n21540, C1 => n15764, C2 =>
                           n21549, A => n17381, ZN => n17377);
   U16592 : AOI22_X1 port map( A1 => n21556, A2 => n19853, B1 => n21251, B2 => 
                           n8690, ZN => n17381);
   U16593 : OAI221_X1 port map( B1 => n15693, B2 => n21539, C1 => n15799, C2 =>
                           n21548, A => n17392, ZN => n17388);
   U16594 : AOI22_X1 port map( A1 => n21579, A2 => n19854, B1 => n21250, B2 => 
                           n8694, ZN => n17392);
   U16595 : OAI221_X1 port map( B1 => n15657, B2 => n21542, C1 => n15763, C2 =>
                           n21545, A => n17334, ZN => n17330);
   U16596 : AOI22_X1 port map( A1 => n21557, A2 => n19855, B1 => n21253, B2 => 
                           n8679, ZN => n17334);
   U16597 : OAI221_X1 port map( B1 => n15692, B2 => n21541, C1 => n15798, C2 =>
                           n21544, A => n17345, ZN => n17341);
   U16598 : AOI22_X1 port map( A1 => n21582, A2 => n19856, B1 => n21252, B2 => 
                           n8683, ZN => n17345);
   U16599 : OAI221_X1 port map( B1 => n15656, B2 => n21539, C1 => n15762, C2 =>
                           n21545, A => n17287, ZN => n17283);
   U16600 : AOI22_X1 port map( A1 => n21559, A2 => n19857, B1 => n21255, B2 => 
                           n8668, ZN => n17287);
   U16601 : OAI221_X1 port map( B1 => n15691, B2 => n21538, C1 => n15797, C2 =>
                           n21546, A => n17298, ZN => n17294);
   U16602 : AOI22_X1 port map( A1 => n21558, A2 => n19858, B1 => n21254, B2 => 
                           n8672, ZN => n17298);
   U16603 : OAI221_X1 port map( B1 => n15655, B2 => n21538, C1 => n15761, C2 =>
                           n21548, A => n17240, ZN => n17236);
   U16604 : AOI22_X1 port map( A1 => n21561, A2 => n19859, B1 => n21257, B2 => 
                           n8657, ZN => n17240);
   U16605 : OAI221_X1 port map( B1 => n15690, B2 => n21543, C1 => n15796, C2 =>
                           n21547, A => n17251, ZN => n17247);
   U16606 : AOI22_X1 port map( A1 => n21560, A2 => n19860, B1 => n21256, B2 => 
                           n8661, ZN => n17251);
   U16607 : OAI221_X1 port map( B1 => n15654, B2 => n21540, C1 => n15760, C2 =>
                           n21544, A => n17193, ZN => n17189);
   U16608 : AOI22_X1 port map( A1 => n21563, A2 => n19861, B1 => n21259, B2 => 
                           n8646, ZN => n17193);
   U16609 : OAI221_X1 port map( B1 => n15689, B2 => n21539, C1 => n15795, C2 =>
                           n21549, A => n17204, ZN => n17200);
   U16610 : AOI22_X1 port map( A1 => n21562, A2 => n19862, B1 => n21258, B2 => 
                           n8650, ZN => n17204);
   U16611 : OAI221_X1 port map( B1 => n15653, B2 => n21540, C1 => n15759, C2 =>
                           n21546, A => n17146, ZN => n17142);
   U16612 : AOI22_X1 port map( A1 => n21565, A2 => n19863, B1 => n21261, B2 => 
                           n8635, ZN => n17146);
   U16613 : OAI221_X1 port map( B1 => n15688, B2 => n21539, C1 => n15794, C2 =>
                           n21545, A => n17157, ZN => n17153);
   U16614 : AOI22_X1 port map( A1 => n21564, A2 => n19864, B1 => n21260, B2 => 
                           n8639, ZN => n17157);
   U16615 : OAI221_X1 port map( B1 => n15652, B2 => n21542, C1 => n15758, C2 =>
                           n21547, A => n17099, ZN => n17095);
   U16616 : AOI22_X1 port map( A1 => n21567, A2 => n19865, B1 => n21263, B2 => 
                           n8624, ZN => n17099);
   U16617 : OAI221_X1 port map( B1 => n15687, B2 => n21541, C1 => n15793, C2 =>
                           n21546, A => n17110, ZN => n17106);
   U16618 : AOI22_X1 port map( A1 => n21566, A2 => n19866, B1 => n21262, B2 => 
                           n8628, ZN => n17110);
   U16619 : OAI221_X1 port map( B1 => n15651, B2 => n21538, C1 => n15757, C2 =>
                           n21549, A => n17052, ZN => n17048);
   U16620 : AOI22_X1 port map( A1 => n21569, A2 => n19867, B1 => n21265, B2 => 
                           n8613, ZN => n17052);
   U16621 : OAI221_X1 port map( B1 => n15686, B2 => n21543, C1 => n15792, C2 =>
                           n21548, A => n17063, ZN => n17059);
   U16622 : AOI22_X1 port map( A1 => n21568, A2 => n19868, B1 => n21264, B2 => 
                           n8617, ZN => n17063);
   U16623 : OAI221_X1 port map( B1 => n15650, B2 => n21541, C1 => n15756, C2 =>
                           n21547, A => n17005, ZN => n17001);
   U16624 : AOI22_X1 port map( A1 => n21581, A2 => n19869, B1 => n21275, B2 => 
                           n8602, ZN => n17005);
   U16625 : OAI221_X1 port map( B1 => n15685, B2 => n21540, C1 => n15791, C2 =>
                           n21544, A => n17016, ZN => n17012);
   U16626 : AOI22_X1 port map( A1 => n21578, A2 => n19870, B1 => n21275, B2 => 
                           n8606, ZN => n17016);
   U16627 : OAI221_X1 port map( B1 => n15649, B2 => n21540, C1 => n15755, C2 =>
                           n21546, A => n16958, ZN => n16954);
   U16628 : AOI22_X1 port map( A1 => n21575, A2 => n19871, B1 => n21269, B2 => 
                           n8591, ZN => n16958);
   U16629 : OAI221_X1 port map( B1 => n15684, B2 => n21539, C1 => n15790, C2 =>
                           n21545, A => n16969, ZN => n16965);
   U16630 : AOI22_X1 port map( A1 => n21574, A2 => n19872, B1 => n21269, B2 => 
                           n8595, ZN => n16969);
   U16631 : OAI221_X1 port map( B1 => n15648, B2 => n21542, C1 => n15754, C2 =>
                           n21548, A => n16889, ZN => n16879);
   U16632 : AOI22_X1 port map( A1 => n21576, A2 => n19873, B1 => n21271, B2 => 
                           n8580, ZN => n16889);
   U16633 : OAI221_X1 port map( B1 => n15683, B2 => n21541, C1 => n15789, C2 =>
                           n21547, A => n16910, ZN => n16906);
   U16634 : AOI22_X1 port map( A1 => n21574, A2 => n19874, B1 => n21269, B2 => 
                           n8584, ZN => n16910);
   U16635 : OAI221_X1 port map( B1 => n7457, B2 => n20796, C1 => n16553, C2 => 
                           n20729, A => n19653, ZN => n19648);
   U16636 : AOI22_X1 port map( A1 => n20751, A2 => n9367, B1 => n20813, B2 => 
                           n8919, ZN => n19653);
   U16637 : OAI221_X1 port map( B1 => n7456, B2 => n20795, C1 => n7454, C2 => 
                           n20734, A => n19668, ZN => n19656);
   U16638 : AOI22_X1 port map( A1 => n20780, A2 => n9371, B1 => n20812, B2 => 
                           n8923, ZN => n19668);
   U16639 : OAI221_X1 port map( B1 => n7489, B2 => n20792, C1 => n16552, C2 => 
                           n20731, A => n19602, ZN => n19597);
   U16640 : AOI22_X1 port map( A1 => n20760, A2 => n9356, B1 => n20815, B2 => 
                           n8908, ZN => n19602);
   U16641 : OAI221_X1 port map( B1 => n7488, B2 => n20797, C1 => n7486, C2 => 
                           n20730, A => n19610, ZN => n19605);
   U16642 : AOI22_X1 port map( A1 => n20759, A2 => n9360, B1 => n20814, B2 => 
                           n8912, ZN => n19610);
   U16643 : OAI221_X1 port map( B1 => n7521, B2 => n20792, C1 => n16551, C2 => 
                           n20729, A => n19565, ZN => n19560);
   U16644 : AOI22_X1 port map( A1 => n20762, A2 => n9345, B1 => n20817, B2 => 
                           n8897, ZN => n19565);
   U16645 : OAI221_X1 port map( B1 => n7520, B2 => n20797, C1 => n7518, C2 => 
                           n20732, A => n19573, ZN => n19568);
   U16646 : AOI22_X1 port map( A1 => n20761, A2 => n9349, B1 => n20816, B2 => 
                           n8901, ZN => n19573);
   U16647 : OAI221_X1 port map( B1 => n7553, B2 => n20794, C1 => n16550, C2 => 
                           n20734, A => n19528, ZN => n19523);
   U16648 : AOI22_X1 port map( A1 => n20764, A2 => n9334, B1 => n20819, B2 => 
                           n8886, ZN => n19528);
   U16649 : OAI221_X1 port map( B1 => n7552, B2 => n20793, C1 => n7550, C2 => 
                           n20733, A => n19536, ZN => n19531);
   U16650 : AOI22_X1 port map( A1 => n20763, A2 => n9338, B1 => n20818, B2 => 
                           n8890, ZN => n19536);
   U16651 : OAI221_X1 port map( B1 => n7585, B2 => n20796, C1 => n16549, C2 => 
                           n20730, A => n19491, ZN => n19486);
   U16652 : AOI22_X1 port map( A1 => n20766, A2 => n9323, B1 => n20821, B2 => 
                           n8875, ZN => n19491);
   U16653 : OAI221_X1 port map( B1 => n7584, B2 => n20795, C1 => n7582, C2 => 
                           n20729, A => n19499, ZN => n19494);
   U16654 : AOI22_X1 port map( A1 => n20765, A2 => n9327, B1 => n20820, B2 => 
                           n8879, ZN => n19499);
   U16655 : OAI221_X1 port map( B1 => n7617, B2 => n20793, C1 => n16548, C2 => 
                           n20730, A => n19454, ZN => n19449);
   U16656 : AOI22_X1 port map( A1 => n20768, A2 => n9312, B1 => n20823, B2 => 
                           n8864, ZN => n19454);
   U16657 : OAI221_X1 port map( B1 => n7616, B2 => n20792, C1 => n7614, C2 => 
                           n20731, A => n19462, ZN => n19457);
   U16658 : AOI22_X1 port map( A1 => n20767, A2 => n9316, B1 => n20822, B2 => 
                           n8868, ZN => n19462);
   U16659 : OAI221_X1 port map( B1 => n7649, B2 => n20792, C1 => n16547, C2 => 
                           n20733, A => n19417, ZN => n19412);
   U16660 : AOI22_X1 port map( A1 => n20770, A2 => n9301, B1 => n20825, B2 => 
                           n8853, ZN => n19417);
   U16661 : OAI221_X1 port map( B1 => n7648, B2 => n20797, C1 => n7646, C2 => 
                           n20732, A => n19425, ZN => n19420);
   U16662 : AOI22_X1 port map( A1 => n20769, A2 => n9305, B1 => n20824, B2 => 
                           n8857, ZN => n19425);
   U16663 : OAI221_X1 port map( B1 => n7681, B2 => n20794, C1 => n16546, C2 => 
                           n20729, A => n19380, ZN => n19375);
   U16664 : AOI22_X1 port map( A1 => n20775, A2 => n9290, B1 => n20827, B2 => 
                           n8842, ZN => n19380);
   U16665 : OAI221_X1 port map( B1 => n7680, B2 => n20793, C1 => n7678, C2 => 
                           n20734, A => n19388, ZN => n19383);
   U16666 : AOI22_X1 port map( A1 => n20775, A2 => n9294, B1 => n20826, B2 => 
                           n8846, ZN => n19388);
   U16667 : OAI221_X1 port map( B1 => n7713, B2 => n20794, C1 => n16545, C2 => 
                           n20731, A => n19343, ZN => n19338);
   U16668 : AOI22_X1 port map( A1 => n20776, A2 => n9279, B1 => n20831, B2 => 
                           n8831, ZN => n19343);
   U16669 : OAI221_X1 port map( B1 => n7712, B2 => n20793, C1 => n7710, C2 => 
                           n20730, A => n19351, ZN => n19346);
   U16670 : AOI22_X1 port map( A1 => n20775, A2 => n9283, B1 => n20831, B2 => 
                           n8835, ZN => n19351);
   U16671 : OAI221_X1 port map( B1 => n7745, B2 => n20796, C1 => n16544, C2 => 
                           n20732, A => n19306, ZN => n19301);
   U16672 : AOI22_X1 port map( A1 => n20777, A2 => n9268, B1 => n20832, B2 => 
                           n8820, ZN => n19306);
   U16673 : OAI221_X1 port map( B1 => n7744, B2 => n20795, C1 => n7742, C2 => 
                           n20731, A => n19314, ZN => n19309);
   U16674 : AOI22_X1 port map( A1 => n20776, A2 => n9272, B1 => n20831, B2 => 
                           n8824, ZN => n19314);
   U16675 : OAI221_X1 port map( B1 => n7777, B2 => n20792, C1 => n16543, C2 => 
                           n20734, A => n19269, ZN => n19264);
   U16676 : AOI22_X1 port map( A1 => n20778, A2 => n9257, B1 => n20833, B2 => 
                           n8809, ZN => n19269);
   U16677 : OAI221_X1 port map( B1 => n7776, B2 => n20797, C1 => n7774, C2 => 
                           n20733, A => n19277, ZN => n19272);
   U16678 : AOI22_X1 port map( A1 => n20779, A2 => n9261, B1 => n20832, B2 => 
                           n8813, ZN => n19277);
   U16679 : OAI221_X1 port map( B1 => n7809, B2 => n20795, C1 => n16542, C2 => 
                           n20732, A => n19232, ZN => n19227);
   U16680 : AOI22_X1 port map( A1 => n20780, A2 => n9246, B1 => n20834, B2 => 
                           n8798, ZN => n19232);
   U16681 : OAI221_X1 port map( B1 => n7808, B2 => n20794, C1 => n7806, C2 => 
                           n20729, A => n19240, ZN => n19235);
   U16682 : AOI22_X1 port map( A1 => n20779, A2 => n9250, B1 => n20834, B2 => 
                           n8802, ZN => n19240);
   U16683 : OAI221_X1 port map( B1 => n7841, B2 => n20794, C1 => n16541, C2 => 
                           n20731, A => n19195, ZN => n19190);
   U16684 : AOI22_X1 port map( A1 => n20781, A2 => n9235, B1 => n20835, B2 => 
                           n8787, ZN => n19195);
   U16685 : OAI221_X1 port map( B1 => n7840, B2 => n20793, C1 => n7838, C2 => 
                           n20730, A => n19203, ZN => n19198);
   U16686 : AOI22_X1 port map( A1 => n20781, A2 => n9239, B1 => n20834, B2 => 
                           n8791, ZN => n19203);
   U16687 : OAI221_X1 port map( B1 => n7873, B2 => n20796, C1 => n16540, C2 => 
                           n20733, A => n19158, ZN => n19153);
   U16688 : AOI22_X1 port map( A1 => n20782, A2 => n9224, B1 => n20836, B2 => 
                           n8776, ZN => n19158);
   U16689 : OAI221_X1 port map( B1 => n7872, B2 => n20795, C1 => n7870, C2 => 
                           n20732, A => n19166, ZN => n19161);
   U16690 : AOI22_X1 port map( A1 => n20782, A2 => n9228, B1 => n20836, B2 => 
                           n8780, ZN => n19166);
   U16691 : OAI221_X1 port map( B1 => n7905, B2 => n20796, C1 => n16539, C2 => 
                           n20733, A => n19121, ZN => n19116);
   U16692 : AOI22_X1 port map( A1 => n20778, A2 => n9213, B1 => n20833, B2 => 
                           n8765, ZN => n19121);
   U16693 : OAI221_X1 port map( B1 => n7904, B2 => n20795, C1 => n16574, C2 => 
                           n20734, A => n19129, ZN => n19124);
   U16694 : AOI22_X1 port map( A1 => n20758, A2 => n9217, B1 => n20838, B2 => 
                           n8769, ZN => n19129);
   U16695 : OAI221_X1 port map( B1 => n7937, B2 => n20792, C1 => n16538, C2 => 
                           n20730, A => n19084, ZN => n19079);
   U16696 : AOI22_X1 port map( A1 => n20778, A2 => n9202, B1 => n20834, B2 => 
                           n8754, ZN => n19084);
   U16697 : OAI221_X1 port map( B1 => n7936, B2 => n20797, C1 => n16573, C2 => 
                           n20729, A => n19092, ZN => n19087);
   U16698 : AOI22_X1 port map( A1 => n20779, A2 => n9206, B1 => n20834, B2 => 
                           n8758, ZN => n19092);
   U16699 : OAI221_X1 port map( B1 => n7969, B2 => n20794, C1 => n16537, C2 => 
                           n20732, A => n19047, ZN => n19042);
   U16700 : AOI22_X1 port map( A1 => n20780, A2 => n9191, B1 => n20835, B2 => 
                           n8743, ZN => n19047);
   U16701 : OAI221_X1 port map( B1 => n7968, B2 => n20793, C1 => n16572, C2 => 
                           n20731, A => n19055, ZN => n19050);
   U16702 : AOI22_X1 port map( A1 => n20779, A2 => n9195, B1 => n20834, B2 => 
                           n8747, ZN => n19055);
   U16703 : OAI221_X1 port map( B1 => n8001, B2 => n20797, C1 => n16536, C2 => 
                           n20734, A => n19010, ZN => n19005);
   U16704 : AOI22_X1 port map( A1 => n20781, A2 => n9180, B1 => n20832, B2 => 
                           n8732, ZN => n19010);
   U16705 : OAI221_X1 port map( B1 => n8000, B2 => n20796, C1 => n16571, C2 => 
                           n20733, A => n19018, ZN => n19013);
   U16706 : AOI22_X1 port map( A1 => n20780, A2 => n9184, B1 => n20836, B2 => 
                           n8736, ZN => n19018);
   U16707 : OAI221_X1 port map( B1 => n8032, B2 => n20795, C1 => n16570, C2 => 
                           n20734, A => n18981, ZN => n18976);
   U16708 : AOI22_X1 port map( A1 => n20782, A2 => n9173, B1 => n20837, B2 => 
                           n8725, ZN => n18981);
   U16709 : OAI221_X1 port map( B1 => n8064, B2 => n20797, C1 => n16569, C2 => 
                           n20730, A => n18944, ZN => n18939);
   U16710 : AOI22_X1 port map( A1 => n20783, A2 => n9162, B1 => n20837, B2 => 
                           n8714, ZN => n18944);
   U16711 : OAI221_X1 port map( B1 => n8096, B2 => n20797, C1 => n16568, C2 => 
                           n20732, A => n18907, ZN => n18902);
   U16712 : AOI22_X1 port map( A1 => n20757, A2 => n9151, B1 => n20838, B2 => 
                           n8703, ZN => n18907);
   U16713 : OAI221_X1 port map( B1 => n8128, B2 => n20793, C1 => n16567, C2 => 
                           n20733, A => n18870, ZN => n18865);
   U16714 : AOI22_X1 port map( A1 => n20758, A2 => n9140, B1 => n20812, B2 => 
                           n8692, ZN => n18870);
   U16715 : OAI221_X1 port map( B1 => n8161, B2 => n20796, C1 => n16531, C2 => 
                           n20730, A => n18825, ZN => n18820);
   U16716 : AOI22_X1 port map( A1 => n20783, A2 => n9125, B1 => n20813, B2 => 
                           n8677, ZN => n18825);
   U16717 : OAI221_X1 port map( B1 => n8160, B2 => n20795, C1 => n16566, C2 => 
                           n20729, A => n18833, ZN => n18828);
   U16718 : AOI22_X1 port map( A1 => n20779, A2 => n9129, B1 => n20837, B2 => 
                           n8681, ZN => n18833);
   U16719 : OAI221_X1 port map( B1 => n8193, B2 => n20793, C1 => n16530, C2 => 
                           n20730, A => n18788, ZN => n18783);
   U16720 : AOI22_X1 port map( A1 => n20760, A2 => n9114, B1 => n20815, B2 => 
                           n8666, ZN => n18788);
   U16721 : OAI221_X1 port map( B1 => n8192, B2 => n20792, C1 => n16565, C2 => 
                           n20731, A => n18796, ZN => n18791);
   U16722 : AOI22_X1 port map( A1 => n20759, A2 => n9118, B1 => n20814, B2 => 
                           n8670, ZN => n18796);
   U16723 : OAI221_X1 port map( B1 => n8225, B2 => n20792, C1 => n16529, C2 => 
                           n20733, A => n18751, ZN => n18746);
   U16724 : AOI22_X1 port map( A1 => n20762, A2 => n9103, B1 => n20817, B2 => 
                           n8655, ZN => n18751);
   U16725 : OAI221_X1 port map( B1 => n8224, B2 => n20797, C1 => n16564, C2 => 
                           n20732, A => n18759, ZN => n18754);
   U16726 : AOI22_X1 port map( A1 => n20761, A2 => n9107, B1 => n20816, B2 => 
                           n8659, ZN => n18759);
   U16727 : OAI221_X1 port map( B1 => n8257, B2 => n20794, C1 => n16528, C2 => 
                           n20729, A => n18714, ZN => n18709);
   U16728 : AOI22_X1 port map( A1 => n20764, A2 => n9092, B1 => n20819, B2 => 
                           n8644, ZN => n18714);
   U16729 : OAI221_X1 port map( B1 => n8256, B2 => n20793, C1 => n16563, C2 => 
                           n20734, A => n18722, ZN => n18717);
   U16730 : AOI22_X1 port map( A1 => n20763, A2 => n9096, B1 => n20818, B2 => 
                           n8648, ZN => n18722);
   U16731 : OAI221_X1 port map( B1 => n8289, B2 => n20794, C1 => n16527, C2 => 
                           n20731, A => n18677, ZN => n18672);
   U16732 : AOI22_X1 port map( A1 => n20766, A2 => n9081, B1 => n20821, B2 => 
                           n8633, ZN => n18677);
   U16733 : OAI221_X1 port map( B1 => n8288, B2 => n20793, C1 => n16562, C2 => 
                           n20730, A => n18685, ZN => n18680);
   U16734 : AOI22_X1 port map( A1 => n20765, A2 => n9085, B1 => n20820, B2 => 
                           n8637, ZN => n18685);
   U16735 : OAI221_X1 port map( B1 => n8321, B2 => n20796, C1 => n16526, C2 => 
                           n20732, A => n18640, ZN => n18635);
   U16736 : AOI22_X1 port map( A1 => n20768, A2 => n9070, B1 => n20823, B2 => 
                           n8622, ZN => n18640);
   U16737 : OAI221_X1 port map( B1 => n8320, B2 => n20795, C1 => n16561, C2 => 
                           n20731, A => n18648, ZN => n18643);
   U16738 : AOI22_X1 port map( A1 => n20767, A2 => n9074, B1 => n20822, B2 => 
                           n8626, ZN => n18648);
   U16739 : OAI221_X1 port map( B1 => n8353, B2 => n20792, C1 => n16525, C2 => 
                           n20734, A => n18603, ZN => n18598);
   U16740 : AOI22_X1 port map( A1 => n20770, A2 => n9059, B1 => n20825, B2 => 
                           n8611, ZN => n18603);
   U16741 : OAI221_X1 port map( B1 => n8352, B2 => n20797, C1 => n16560, C2 => 
                           n20733, A => n18611, ZN => n18606);
   U16742 : AOI22_X1 port map( A1 => n20769, A2 => n9063, B1 => n20824, B2 => 
                           n8615, ZN => n18611);
   U16743 : OAI221_X1 port map( B1 => n8385, B2 => n20795, C1 => n16524, C2 => 
                           n20732, A => n18566, ZN => n18561);
   U16744 : AOI22_X1 port map( A1 => n20775, A2 => n9048, B1 => n20827, B2 => 
                           n8600, ZN => n18566);
   U16745 : OAI221_X1 port map( B1 => n8384, B2 => n20794, C1 => n16559, C2 => 
                           n20729, A => n18574, ZN => n18569);
   U16746 : AOI22_X1 port map( A1 => n20775, A2 => n9052, B1 => n20826, B2 => 
                           n8604, ZN => n18574);
   U16747 : OAI221_X1 port map( B1 => n8417, B2 => n20794, C1 => n16523, C2 => 
                           n20731, A => n18529, ZN => n18524);
   U16748 : AOI22_X1 port map( A1 => n20776, A2 => n9037, B1 => n20831, B2 => 
                           n8589, ZN => n18529);
   U16749 : OAI221_X1 port map( B1 => n8416, B2 => n20793, C1 => n16558, C2 => 
                           n20730, A => n18537, ZN => n18532);
   U16750 : AOI22_X1 port map( A1 => n20775, A2 => n9041, B1 => n20831, B2 => 
                           n8593, ZN => n18537);
   U16751 : OAI221_X1 port map( B1 => n8449, B2 => n20796, C1 => n16522, C2 => 
                           n20733, A => n18474, ZN => n18459);
   U16752 : AOI22_X1 port map( A1 => n20777, A2 => n9026, B1 => n20833, B2 => 
                           n8578, ZN => n18474);
   U16753 : OAI221_X1 port map( B1 => n8448, B2 => n20795, C1 => n16557, C2 => 
                           n20732, A => n18488, ZN => n18483);
   U16754 : AOI22_X1 port map( A1 => n20777, A2 => n9030, B1 => n20831, B2 => 
                           n8582, ZN => n18488);
   U16755 : OAI221_X1 port map( B1 => n7457, B2 => n21353, C1 => n16553, C2 => 
                           n21286, A => n18384, ZN => n18377);
   U16756 : AOI22_X1 port map( A1 => n21308, A2 => n9367, B1 => n21370, B2 => 
                           n8919, ZN => n18384);
   U16757 : OAI221_X1 port map( B1 => n7456, B2 => n21352, C1 => n7454, C2 => 
                           n21291, A => n18402, ZN => n18388);
   U16758 : AOI22_X1 port map( A1 => n21337, A2 => n9371, B1 => n21369, B2 => 
                           n8923, ZN => n18402);
   U16759 : OAI221_X1 port map( B1 => n7489, B2 => n21349, C1 => n16552, C2 => 
                           n21288, A => n18323, ZN => n18316);
   U16760 : AOI22_X1 port map( A1 => n21317, A2 => n9356, B1 => n21372, B2 => 
                           n8908, ZN => n18323);
   U16761 : OAI221_X1 port map( B1 => n7488, B2 => n21354, C1 => n7486, C2 => 
                           n21287, A => n18334, ZN => n18327);
   U16762 : AOI22_X1 port map( A1 => n21316, A2 => n9360, B1 => n21371, B2 => 
                           n8912, ZN => n18334);
   U16763 : OAI221_X1 port map( B1 => n7521, B2 => n21349, C1 => n16551, C2 => 
                           n21286, A => n18276, ZN => n18269);
   U16764 : AOI22_X1 port map( A1 => n21319, A2 => n9345, B1 => n21374, B2 => 
                           n8897, ZN => n18276);
   U16765 : OAI221_X1 port map( B1 => n7520, B2 => n21354, C1 => n7518, C2 => 
                           n21289, A => n18287, ZN => n18280);
   U16766 : AOI22_X1 port map( A1 => n21318, A2 => n9349, B1 => n21373, B2 => 
                           n8901, ZN => n18287);
   U16767 : OAI221_X1 port map( B1 => n7553, B2 => n21351, C1 => n16550, C2 => 
                           n21291, A => n18229, ZN => n18222);
   U16768 : AOI22_X1 port map( A1 => n21321, A2 => n9334, B1 => n21376, B2 => 
                           n8886, ZN => n18229);
   U16769 : OAI221_X1 port map( B1 => n7552, B2 => n21350, C1 => n7550, C2 => 
                           n21290, A => n18240, ZN => n18233);
   U16770 : AOI22_X1 port map( A1 => n21320, A2 => n9338, B1 => n21375, B2 => 
                           n8890, ZN => n18240);
   U16771 : OAI221_X1 port map( B1 => n7585, B2 => n21353, C1 => n16549, C2 => 
                           n21287, A => n18182, ZN => n18175);
   U16772 : AOI22_X1 port map( A1 => n21323, A2 => n9323, B1 => n21378, B2 => 
                           n8875, ZN => n18182);
   U16773 : OAI221_X1 port map( B1 => n7584, B2 => n21352, C1 => n7582, C2 => 
                           n21286, A => n18193, ZN => n18186);
   U16774 : AOI22_X1 port map( A1 => n21322, A2 => n9327, B1 => n21377, B2 => 
                           n8879, ZN => n18193);
   U16775 : OAI221_X1 port map( B1 => n7617, B2 => n21350, C1 => n16548, C2 => 
                           n21287, A => n18135, ZN => n18128);
   U16776 : AOI22_X1 port map( A1 => n21325, A2 => n9312, B1 => n21380, B2 => 
                           n8864, ZN => n18135);
   U16777 : OAI221_X1 port map( B1 => n7616, B2 => n21349, C1 => n7614, C2 => 
                           n21288, A => n18146, ZN => n18139);
   U16778 : AOI22_X1 port map( A1 => n21324, A2 => n9316, B1 => n21379, B2 => 
                           n8868, ZN => n18146);
   U16779 : OAI221_X1 port map( B1 => n7649, B2 => n21349, C1 => n16547, C2 => 
                           n21290, A => n18088, ZN => n18081);
   U16780 : AOI22_X1 port map( A1 => n21327, A2 => n9301, B1 => n21382, B2 => 
                           n8853, ZN => n18088);
   U16781 : OAI221_X1 port map( B1 => n7648, B2 => n21354, C1 => n7646, C2 => 
                           n21289, A => n18099, ZN => n18092);
   U16782 : AOI22_X1 port map( A1 => n21326, A2 => n9305, B1 => n21381, B2 => 
                           n8857, ZN => n18099);
   U16783 : OAI221_X1 port map( B1 => n7681, B2 => n21351, C1 => n16546, C2 => 
                           n21286, A => n18041, ZN => n18034);
   U16784 : AOI22_X1 port map( A1 => n21332, A2 => n9290, B1 => n21384, B2 => 
                           n8842, ZN => n18041);
   U16785 : OAI221_X1 port map( B1 => n7680, B2 => n21350, C1 => n7678, C2 => 
                           n21291, A => n18052, ZN => n18045);
   U16786 : AOI22_X1 port map( A1 => n21332, A2 => n9294, B1 => n21383, B2 => 
                           n8846, ZN => n18052);
   U16787 : OAI221_X1 port map( B1 => n7713, B2 => n21351, C1 => n16545, C2 => 
                           n21288, A => n17994, ZN => n17987);
   U16788 : AOI22_X1 port map( A1 => n21333, A2 => n9279, B1 => n21388, B2 => 
                           n8831, ZN => n17994);
   U16789 : OAI221_X1 port map( B1 => n7712, B2 => n21350, C1 => n7710, C2 => 
                           n21287, A => n18005, ZN => n17998);
   U16790 : AOI22_X1 port map( A1 => n21332, A2 => n9283, B1 => n21388, B2 => 
                           n8835, ZN => n18005);
   U16791 : OAI221_X1 port map( B1 => n7745, B2 => n21353, C1 => n16544, C2 => 
                           n21289, A => n17947, ZN => n17940);
   U16792 : AOI22_X1 port map( A1 => n21334, A2 => n9268, B1 => n21389, B2 => 
                           n8820, ZN => n17947);
   U16793 : OAI221_X1 port map( B1 => n7744, B2 => n21352, C1 => n7742, C2 => 
                           n21288, A => n17958, ZN => n17951);
   U16794 : AOI22_X1 port map( A1 => n21333, A2 => n9272, B1 => n21388, B2 => 
                           n8824, ZN => n17958);
   U16795 : OAI221_X1 port map( B1 => n7777, B2 => n21349, C1 => n16543, C2 => 
                           n21291, A => n17900, ZN => n17893);
   U16796 : AOI22_X1 port map( A1 => n21335, A2 => n9257, B1 => n21390, B2 => 
                           n8809, ZN => n17900);
   U16797 : OAI221_X1 port map( B1 => n7776, B2 => n21354, C1 => n7774, C2 => 
                           n21290, A => n17911, ZN => n17904);
   U16798 : AOI22_X1 port map( A1 => n21336, A2 => n9261, B1 => n21389, B2 => 
                           n8813, ZN => n17911);
   U16799 : OAI221_X1 port map( B1 => n7809, B2 => n21352, C1 => n16542, C2 => 
                           n21289, A => n17853, ZN => n17846);
   U16800 : AOI22_X1 port map( A1 => n21337, A2 => n9246, B1 => n21391, B2 => 
                           n8798, ZN => n17853);
   U16801 : OAI221_X1 port map( B1 => n7808, B2 => n21351, C1 => n7806, C2 => 
                           n21286, A => n17864, ZN => n17857);
   U16802 : AOI22_X1 port map( A1 => n21336, A2 => n9250, B1 => n21391, B2 => 
                           n8802, ZN => n17864);
   U16803 : OAI221_X1 port map( B1 => n7841, B2 => n21351, C1 => n16541, C2 => 
                           n21288, A => n17806, ZN => n17799);
   U16804 : AOI22_X1 port map( A1 => n21338, A2 => n9235, B1 => n21392, B2 => 
                           n8787, ZN => n17806);
   U16805 : OAI221_X1 port map( B1 => n7840, B2 => n21350, C1 => n7838, C2 => 
                           n21287, A => n17817, ZN => n17810);
   U16806 : AOI22_X1 port map( A1 => n21338, A2 => n9239, B1 => n21391, B2 => 
                           n8791, ZN => n17817);
   U16807 : OAI221_X1 port map( B1 => n7873, B2 => n21353, C1 => n16540, C2 => 
                           n21290, A => n17759, ZN => n17752);
   U16808 : AOI22_X1 port map( A1 => n21339, A2 => n9224, B1 => n21393, B2 => 
                           n8776, ZN => n17759);
   U16809 : OAI221_X1 port map( B1 => n7872, B2 => n21352, C1 => n7870, C2 => 
                           n21289, A => n17770, ZN => n17763);
   U16810 : AOI22_X1 port map( A1 => n21339, A2 => n9228, B1 => n21393, B2 => 
                           n8780, ZN => n17770);
   U16811 : OAI221_X1 port map( B1 => n7905, B2 => n21353, C1 => n16539, C2 => 
                           n21290, A => n17712, ZN => n17705);
   U16812 : AOI22_X1 port map( A1 => n21335, A2 => n9213, B1 => n21390, B2 => 
                           n8765, ZN => n17712);
   U16813 : OAI221_X1 port map( B1 => n7904, B2 => n21352, C1 => n16574, C2 => 
                           n21291, A => n17723, ZN => n17716);
   U16814 : AOI22_X1 port map( A1 => n21315, A2 => n9217, B1 => n21395, B2 => 
                           n8769, ZN => n17723);
   U16815 : OAI221_X1 port map( B1 => n7937, B2 => n21349, C1 => n16538, C2 => 
                           n21287, A => n17665, ZN => n17658);
   U16816 : AOI22_X1 port map( A1 => n21335, A2 => n9202, B1 => n21391, B2 => 
                           n8754, ZN => n17665);
   U16817 : OAI221_X1 port map( B1 => n7936, B2 => n21354, C1 => n16573, C2 => 
                           n21286, A => n17676, ZN => n17669);
   U16818 : AOI22_X1 port map( A1 => n21336, A2 => n9206, B1 => n21391, B2 => 
                           n8758, ZN => n17676);
   U16819 : OAI221_X1 port map( B1 => n7969, B2 => n21351, C1 => n16537, C2 => 
                           n21289, A => n17618, ZN => n17611);
   U16820 : AOI22_X1 port map( A1 => n21337, A2 => n9191, B1 => n21392, B2 => 
                           n8743, ZN => n17618);
   U16821 : OAI221_X1 port map( B1 => n7968, B2 => n21350, C1 => n16572, C2 => 
                           n21288, A => n17629, ZN => n17622);
   U16822 : AOI22_X1 port map( A1 => n21336, A2 => n9195, B1 => n21391, B2 => 
                           n8747, ZN => n17629);
   U16823 : OAI221_X1 port map( B1 => n8001, B2 => n21354, C1 => n16536, C2 => 
                           n21291, A => n17571, ZN => n17564);
   U16824 : AOI22_X1 port map( A1 => n21338, A2 => n9180, B1 => n21389, B2 => 
                           n8732, ZN => n17571);
   U16825 : OAI221_X1 port map( B1 => n8000, B2 => n21353, C1 => n16571, C2 => 
                           n21290, A => n17582, ZN => n17575);
   U16826 : AOI22_X1 port map( A1 => n21337, A2 => n9184, B1 => n21393, B2 => 
                           n8736, ZN => n17582);
   U16827 : OAI221_X1 port map( B1 => n8032, B2 => n21352, C1 => n16570, C2 => 
                           n21291, A => n17535, ZN => n17528);
   U16828 : AOI22_X1 port map( A1 => n21339, A2 => n9173, B1 => n21394, B2 => 
                           n8725, ZN => n17535);
   U16829 : OAI221_X1 port map( B1 => n8064, B2 => n21354, C1 => n16569, C2 => 
                           n21287, A => n17488, ZN => n17481);
   U16830 : AOI22_X1 port map( A1 => n21340, A2 => n9162, B1 => n21394, B2 => 
                           n8714, ZN => n17488);
   U16831 : OAI221_X1 port map( B1 => n8096, B2 => n21354, C1 => n16568, C2 => 
                           n21289, A => n17441, ZN => n17434);
   U16832 : AOI22_X1 port map( A1 => n21314, A2 => n9151, B1 => n21395, B2 => 
                           n8703, ZN => n17441);
   U16833 : OAI221_X1 port map( B1 => n8128, B2 => n21350, C1 => n16567, C2 => 
                           n21290, A => n17394, ZN => n17387);
   U16834 : AOI22_X1 port map( A1 => n21315, A2 => n9140, B1 => n21369, B2 => 
                           n8692, ZN => n17394);
   U16835 : OAI221_X1 port map( B1 => n8161, B2 => n21353, C1 => n16531, C2 => 
                           n21287, A => n17336, ZN => n17329);
   U16836 : AOI22_X1 port map( A1 => n21340, A2 => n9125, B1 => n21370, B2 => 
                           n8677, ZN => n17336);
   U16837 : OAI221_X1 port map( B1 => n8160, B2 => n21352, C1 => n16566, C2 => 
                           n21286, A => n17347, ZN => n17340);
   U16838 : AOI22_X1 port map( A1 => n21336, A2 => n9129, B1 => n21394, B2 => 
                           n8681, ZN => n17347);
   U16839 : OAI221_X1 port map( B1 => n8193, B2 => n21350, C1 => n16530, C2 => 
                           n21287, A => n17289, ZN => n17282);
   U16840 : AOI22_X1 port map( A1 => n21317, A2 => n9114, B1 => n21372, B2 => 
                           n8666, ZN => n17289);
   U16841 : OAI221_X1 port map( B1 => n8192, B2 => n21349, C1 => n16565, C2 => 
                           n21288, A => n17300, ZN => n17293);
   U16842 : AOI22_X1 port map( A1 => n21316, A2 => n9118, B1 => n21371, B2 => 
                           n8670, ZN => n17300);
   U16843 : OAI221_X1 port map( B1 => n8225, B2 => n21349, C1 => n16529, C2 => 
                           n21290, A => n17242, ZN => n17235);
   U16844 : AOI22_X1 port map( A1 => n21319, A2 => n9103, B1 => n21374, B2 => 
                           n8655, ZN => n17242);
   U16845 : OAI221_X1 port map( B1 => n8224, B2 => n21354, C1 => n16564, C2 => 
                           n21289, A => n17253, ZN => n17246);
   U16846 : AOI22_X1 port map( A1 => n21318, A2 => n9107, B1 => n21373, B2 => 
                           n8659, ZN => n17253);
   U16847 : OAI221_X1 port map( B1 => n8257, B2 => n21351, C1 => n16528, C2 => 
                           n21286, A => n17195, ZN => n17188);
   U16848 : AOI22_X1 port map( A1 => n21321, A2 => n9092, B1 => n21376, B2 => 
                           n8644, ZN => n17195);
   U16849 : OAI221_X1 port map( B1 => n8256, B2 => n21350, C1 => n16563, C2 => 
                           n21291, A => n17206, ZN => n17199);
   U16850 : AOI22_X1 port map( A1 => n21320, A2 => n9096, B1 => n21375, B2 => 
                           n8648, ZN => n17206);
   U16851 : OAI221_X1 port map( B1 => n8289, B2 => n21351, C1 => n16527, C2 => 
                           n21288, A => n17148, ZN => n17141);
   U16852 : AOI22_X1 port map( A1 => n21323, A2 => n9081, B1 => n21378, B2 => 
                           n8633, ZN => n17148);
   U16853 : OAI221_X1 port map( B1 => n8288, B2 => n21350, C1 => n16562, C2 => 
                           n21287, A => n17159, ZN => n17152);
   U16854 : AOI22_X1 port map( A1 => n21322, A2 => n9085, B1 => n21377, B2 => 
                           n8637, ZN => n17159);
   U16855 : OAI221_X1 port map( B1 => n8321, B2 => n21353, C1 => n16526, C2 => 
                           n21289, A => n17101, ZN => n17094);
   U16856 : AOI22_X1 port map( A1 => n21325, A2 => n9070, B1 => n21380, B2 => 
                           n8622, ZN => n17101);
   U16857 : OAI221_X1 port map( B1 => n8320, B2 => n21352, C1 => n16561, C2 => 
                           n21288, A => n17112, ZN => n17105);
   U16858 : AOI22_X1 port map( A1 => n21324, A2 => n9074, B1 => n21379, B2 => 
                           n8626, ZN => n17112);
   U16859 : OAI221_X1 port map( B1 => n8353, B2 => n21349, C1 => n16525, C2 => 
                           n21291, A => n17054, ZN => n17047);
   U16860 : AOI22_X1 port map( A1 => n21327, A2 => n9059, B1 => n21382, B2 => 
                           n8611, ZN => n17054);
   U16861 : OAI221_X1 port map( B1 => n8352, B2 => n21354, C1 => n16560, C2 => 
                           n21290, A => n17065, ZN => n17058);
   U16862 : AOI22_X1 port map( A1 => n21326, A2 => n9063, B1 => n21381, B2 => 
                           n8615, ZN => n17065);
   U16863 : OAI221_X1 port map( B1 => n8385, B2 => n21352, C1 => n16524, C2 => 
                           n21289, A => n17007, ZN => n17000);
   U16864 : AOI22_X1 port map( A1 => n21332, A2 => n9048, B1 => n21384, B2 => 
                           n8600, ZN => n17007);
   U16865 : OAI221_X1 port map( B1 => n8384, B2 => n21351, C1 => n16559, C2 => 
                           n21286, A => n17018, ZN => n17011);
   U16866 : AOI22_X1 port map( A1 => n21332, A2 => n9052, B1 => n21383, B2 => 
                           n8604, ZN => n17018);
   U16867 : OAI221_X1 port map( B1 => n8417, B2 => n21351, C1 => n16523, C2 => 
                           n21288, A => n16960, ZN => n16953);
   U16868 : AOI22_X1 port map( A1 => n21333, A2 => n9037, B1 => n21388, B2 => 
                           n8589, ZN => n16960);
   U16869 : OAI221_X1 port map( B1 => n8416, B2 => n21350, C1 => n16558, C2 => 
                           n21287, A => n16971, ZN => n16964);
   U16870 : AOI22_X1 port map( A1 => n21332, A2 => n9041, B1 => n21388, B2 => 
                           n8593, ZN => n16971);
   U16871 : OAI221_X1 port map( B1 => n8449, B2 => n21353, C1 => n16522, C2 => 
                           n21290, A => n16895, ZN => n16878);
   U16872 : AOI22_X1 port map( A1 => n21334, A2 => n9026, B1 => n21390, B2 => 
                           n8578, ZN => n16895);
   U16873 : OAI221_X1 port map( B1 => n8448, B2 => n21352, C1 => n16557, C2 => 
                           n21289, A => n16912, ZN => n16905);
   U16874 : AOI22_X1 port map( A1 => n21334, A2 => n9030, B1 => n21388, B2 => 
                           n8582, ZN => n16912);
   U16875 : OAI221_X1 port map( B1 => n16238, B2 => n20863, C1 => n16132, C2 =>
                           n20873, A => n19654, ZN => n19647);
   U16876 : AOI22_X1 port map( A1 => n20952, A2 => n19875, B1 => n20910, B2 => 
                           n9917, ZN => n19654);
   U16877 : OAI221_X1 port map( B1 => n16273, B2 => n20862, C1 => n16167, C2 =>
                           n20878, A => n19669, ZN => n19655);
   U16878 : AOI22_X1 port map( A1 => n20951, A2 => n19876, B1 => n20909, B2 => 
                           n9949, ZN => n19669);
   U16879 : OAI221_X1 port map( B1 => n16237, B2 => n20859, C1 => n16131, C2 =>
                           n20875, A => n19603, ZN => n19596);
   U16880 : AOI22_X1 port map( A1 => n20954, A2 => n19877, B1 => n20912, B2 => 
                           n9916, ZN => n19603);
   U16881 : OAI221_X1 port map( B1 => n16272, B2 => n20864, C1 => n16166, C2 =>
                           n20874, A => n19611, ZN => n19604);
   U16882 : AOI22_X1 port map( A1 => n20953, A2 => n19878, B1 => n20911, B2 => 
                           n9948, ZN => n19611);
   U16883 : OAI221_X1 port map( B1 => n16236, B2 => n20859, C1 => n16130, C2 =>
                           n20873, A => n19566, ZN => n19559);
   U16884 : AOI22_X1 port map( A1 => n20956, A2 => n19879, B1 => n20914, B2 => 
                           n9915, ZN => n19566);
   U16885 : OAI221_X1 port map( B1 => n16271, B2 => n20864, C1 => n16165, C2 =>
                           n20876, A => n19574, ZN => n19567);
   U16886 : AOI22_X1 port map( A1 => n20955, A2 => n19880, B1 => n20913, B2 => 
                           n9947, ZN => n19574);
   U16887 : OAI221_X1 port map( B1 => n16235, B2 => n20861, C1 => n16129, C2 =>
                           n20878, A => n19529, ZN => n19522);
   U16888 : AOI22_X1 port map( A1 => n20958, A2 => n19881, B1 => n20916, B2 => 
                           n9914, ZN => n19529);
   U16889 : OAI221_X1 port map( B1 => n16270, B2 => n20860, C1 => n16164, C2 =>
                           n20877, A => n19537, ZN => n19530);
   U16890 : AOI22_X1 port map( A1 => n20957, A2 => n19882, B1 => n20915, B2 => 
                           n9946, ZN => n19537);
   U16891 : OAI221_X1 port map( B1 => n16234, B2 => n20863, C1 => n16128, C2 =>
                           n20874, A => n19492, ZN => n19485);
   U16892 : AOI22_X1 port map( A1 => n20960, A2 => n19883, B1 => n20918, B2 => 
                           n9913, ZN => n19492);
   U16893 : OAI221_X1 port map( B1 => n16269, B2 => n20862, C1 => n16163, C2 =>
                           n20873, A => n19500, ZN => n19493);
   U16894 : AOI22_X1 port map( A1 => n20959, A2 => n19884, B1 => n20917, B2 => 
                           n9945, ZN => n19500);
   U16895 : OAI221_X1 port map( B1 => n16233, B2 => n20860, C1 => n16127, C2 =>
                           n20874, A => n19455, ZN => n19448);
   U16896 : AOI22_X1 port map( A1 => n20962, A2 => n19885, B1 => n20920, B2 => 
                           n9912, ZN => n19455);
   U16897 : OAI221_X1 port map( B1 => n16268, B2 => n20859, C1 => n16162, C2 =>
                           n20875, A => n19463, ZN => n19456);
   U16898 : AOI22_X1 port map( A1 => n20961, A2 => n19886, B1 => n20919, B2 => 
                           n9944, ZN => n19463);
   U16899 : OAI221_X1 port map( B1 => n16232, B2 => n20859, C1 => n16126, C2 =>
                           n20877, A => n19418, ZN => n19411);
   U16900 : AOI22_X1 port map( A1 => n20964, A2 => n19887, B1 => n20922, B2 => 
                           n9911, ZN => n19418);
   U16901 : OAI221_X1 port map( B1 => n16267, B2 => n20864, C1 => n16161, C2 =>
                           n20876, A => n19426, ZN => n19419);
   U16902 : AOI22_X1 port map( A1 => n20963, A2 => n19888, B1 => n20921, B2 => 
                           n9943, ZN => n19426);
   U16903 : OAI221_X1 port map( B1 => n16231, B2 => n20861, C1 => n16125, C2 =>
                           n20873, A => n19381, ZN => n19374);
   U16904 : AOI22_X1 port map( A1 => n20964, A2 => n19889, B1 => n20924, B2 => 
                           n9910, ZN => n19381);
   U16905 : OAI221_X1 port map( B1 => n16266, B2 => n20860, C1 => n16160, C2 =>
                           n20878, A => n19389, ZN => n19382);
   U16906 : AOI22_X1 port map( A1 => n20977, A2 => n19890, B1 => n20923, B2 => 
                           n9942, ZN => n19389);
   U16907 : OAI221_X1 port map( B1 => n16230, B2 => n20861, C1 => n16124, C2 =>
                           n20875, A => n19344, ZN => n19337);
   U16908 : AOI22_X1 port map( A1 => n20969, A2 => n19891, B1 => n20928, B2 => 
                           n9909, ZN => n19344);
   U16909 : OAI221_X1 port map( B1 => n16265, B2 => n20860, C1 => n16159, C2 =>
                           n20874, A => n19352, ZN => n19345);
   U16910 : AOI22_X1 port map( A1 => n20969, A2 => n19892, B1 => n20928, B2 => 
                           n9941, ZN => n19352);
   U16911 : OAI221_X1 port map( B1 => n16229, B2 => n20863, C1 => n16123, C2 =>
                           n20876, A => n19307, ZN => n19300);
   U16912 : AOI22_X1 port map( A1 => n20970, A2 => n19893, B1 => n20929, B2 => 
                           n9908, ZN => n19307);
   U16913 : OAI221_X1 port map( B1 => n16264, B2 => n20862, C1 => n16158, C2 =>
                           n20875, A => n19315, ZN => n19308);
   U16914 : AOI22_X1 port map( A1 => n20969, A2 => n19894, B1 => n20928, B2 => 
                           n9940, ZN => n19315);
   U16915 : OAI221_X1 port map( B1 => n16228, B2 => n20859, C1 => n16122, C2 =>
                           n20878, A => n19270, ZN => n19263);
   U16916 : AOI22_X1 port map( A1 => n20971, A2 => n19895, B1 => n20930, B2 => 
                           n9907, ZN => n19270);
   U16917 : OAI221_X1 port map( B1 => n16263, B2 => n20864, C1 => n16157, C2 =>
                           n20877, A => n19278, ZN => n19271);
   U16918 : AOI22_X1 port map( A1 => n20970, A2 => n19896, B1 => n20929, B2 => 
                           n9939, ZN => n19278);
   U16919 : OAI221_X1 port map( B1 => n16227, B2 => n20862, C1 => n16121, C2 =>
                           n20876, A => n19233, ZN => n19226);
   U16920 : AOI22_X1 port map( A1 => n20972, A2 => n19897, B1 => n20931, B2 => 
                           n9906, ZN => n19233);
   U16921 : OAI221_X1 port map( B1 => n16262, B2 => n20861, C1 => n16156, C2 =>
                           n20873, A => n19241, ZN => n19234);
   U16922 : AOI22_X1 port map( A1 => n20973, A2 => n19898, B1 => n20931, B2 => 
                           n9938, ZN => n19241);
   U16923 : OAI221_X1 port map( B1 => n16226, B2 => n20861, C1 => n16120, C2 =>
                           n20875, A => n19196, ZN => n19189);
   U16924 : AOI22_X1 port map( A1 => n20974, A2 => n19899, B1 => n20932, B2 => 
                           n9905, ZN => n19196);
   U16925 : OAI221_X1 port map( B1 => n16261, B2 => n20860, C1 => n16155, C2 =>
                           n20874, A => n19204, ZN => n19197);
   U16926 : AOI22_X1 port map( A1 => n20973, A2 => n19900, B1 => n20931, B2 => 
                           n9937, ZN => n19204);
   U16927 : OAI221_X1 port map( B1 => n16225, B2 => n20863, C1 => n16119, C2 =>
                           n20877, A => n19159, ZN => n19152);
   U16928 : AOI22_X1 port map( A1 => n20975, A2 => n19901, B1 => n20933, B2 => 
                           n9904, ZN => n19159);
   U16929 : OAI221_X1 port map( B1 => n16260, B2 => n20862, C1 => n16154, C2 =>
                           n20876, A => n19167, ZN => n19160);
   U16930 : AOI22_X1 port map( A1 => n20975, A2 => n19902, B1 => n20933, B2 => 
                           n9936, ZN => n19167);
   U16931 : OAI221_X1 port map( B1 => n16224, B2 => n20863, C1 => n16118, C2 =>
                           n20877, A => n19122, ZN => n19115);
   U16932 : AOI22_X1 port map( A1 => n20971, A2 => n19903, B1 => n20930, B2 => 
                           n9903, ZN => n19122);
   U16933 : OAI221_X1 port map( B1 => n16259, B2 => n20862, C1 => n16153, C2 =>
                           n20878, A => n19130, ZN => n19123);
   U16934 : AOI22_X1 port map( A1 => n20973, A2 => n19904, B1 => n20935, B2 => 
                           n9935, ZN => n19130);
   U16935 : OAI221_X1 port map( B1 => n16223, B2 => n20859, C1 => n16117, C2 =>
                           n20874, A => n19085, ZN => n19078);
   U16936 : AOI22_X1 port map( A1 => n20972, A2 => n19905, B1 => n20931, B2 => 
                           n9902, ZN => n19085);
   U16937 : OAI221_X1 port map( B1 => n16258, B2 => n20864, C1 => n16152, C2 =>
                           n20873, A => n19093, ZN => n19086);
   U16938 : AOI22_X1 port map( A1 => n20973, A2 => n19906, B1 => n20931, B2 => 
                           n9934, ZN => n19093);
   U16939 : OAI221_X1 port map( B1 => n16222, B2 => n20861, C1 => n16116, C2 =>
                           n20876, A => n19048, ZN => n19041);
   U16940 : AOI22_X1 port map( A1 => n20974, A2 => n19907, B1 => n20932, B2 => 
                           n9901, ZN => n19048);
   U16941 : OAI221_X1 port map( B1 => n16257, B2 => n20860, C1 => n16151, C2 =>
                           n20875, A => n19056, ZN => n19049);
   U16942 : AOI22_X1 port map( A1 => n20973, A2 => n19908, B1 => n20931, B2 => 
                           n9933, ZN => n19056);
   U16943 : OAI221_X1 port map( B1 => n16221, B2 => n20864, C1 => n16115, C2 =>
                           n20878, A => n19011, ZN => n19004);
   U16944 : AOI22_X1 port map( A1 => n20970, A2 => n19909, B1 => n20929, B2 => 
                           n9900, ZN => n19011);
   U16945 : OAI221_X1 port map( B1 => n16256, B2 => n20863, C1 => n16150, C2 =>
                           n20877, A => n19019, ZN => n19012);
   U16946 : AOI22_X1 port map( A1 => n20975, A2 => n19910, B1 => n20933, B2 => 
                           n9932, ZN => n19019);
   U16947 : OAI221_X1 port map( B1 => n16255, B2 => n20862, C1 => n16149, C2 =>
                           n20878, A => n18982, ZN => n18975);
   U16948 : AOI22_X1 port map( A1 => n20976, A2 => n19911, B1 => n20934, B2 => 
                           n9931, ZN => n18982);
   U16949 : OAI221_X1 port map( B1 => n16254, B2 => n20864, C1 => n16148, C2 =>
                           n20874, A => n18945, ZN => n18938);
   U16950 : AOI22_X1 port map( A1 => n20977, A2 => n19912, B1 => n20934, B2 => 
                           n9930, ZN => n18945);
   U16951 : OAI221_X1 port map( B1 => n16253, B2 => n20864, C1 => n16147, C2 =>
                           n20876, A => n18908, ZN => n18901);
   U16952 : AOI22_X1 port map( A1 => n20977, A2 => n19913, B1 => n20935, B2 => 
                           n9929, ZN => n18908);
   U16953 : OAI221_X1 port map( B1 => n16252, B2 => n20860, C1 => n16146, C2 =>
                           n20877, A => n18871, ZN => n18864);
   U16954 : AOI22_X1 port map( A1 => n20972, A2 => n19914, B1 => n20909, B2 => 
                           n9928, ZN => n18871);
   U16955 : OAI221_X1 port map( B1 => n16216, B2 => n20863, C1 => n16110, C2 =>
                           n20874, A => n18826, ZN => n18819);
   U16956 : AOI22_X1 port map( A1 => n20952, A2 => n19915, B1 => n20910, B2 => 
                           n9895, ZN => n18826);
   U16957 : OAI221_X1 port map( B1 => n16251, B2 => n20862, C1 => n16145, C2 =>
                           n20873, A => n18834, ZN => n18827);
   U16958 : AOI22_X1 port map( A1 => n20951, A2 => n19916, B1 => n20934, B2 => 
                           n9927, ZN => n18834);
   U16959 : OAI221_X1 port map( B1 => n16215, B2 => n20860, C1 => n16109, C2 =>
                           n20874, A => n18789, ZN => n18782);
   U16960 : AOI22_X1 port map( A1 => n20954, A2 => n19917, B1 => n20912, B2 => 
                           n9894, ZN => n18789);
   U16961 : OAI221_X1 port map( B1 => n16250, B2 => n20859, C1 => n16144, C2 =>
                           n20875, A => n18797, ZN => n18790);
   U16962 : AOI22_X1 port map( A1 => n20953, A2 => n19918, B1 => n20911, B2 => 
                           n9926, ZN => n18797);
   U16963 : OAI221_X1 port map( B1 => n16214, B2 => n20859, C1 => n16108, C2 =>
                           n20877, A => n18752, ZN => n18745);
   U16964 : AOI22_X1 port map( A1 => n20956, A2 => n19919, B1 => n20914, B2 => 
                           n9893, ZN => n18752);
   U16965 : OAI221_X1 port map( B1 => n16249, B2 => n20864, C1 => n16143, C2 =>
                           n20876, A => n18760, ZN => n18753);
   U16966 : AOI22_X1 port map( A1 => n20955, A2 => n19920, B1 => n20913, B2 => 
                           n9925, ZN => n18760);
   U16967 : OAI221_X1 port map( B1 => n16213, B2 => n20861, C1 => n16107, C2 =>
                           n20873, A => n18715, ZN => n18708);
   U16968 : AOI22_X1 port map( A1 => n20958, A2 => n19921, B1 => n20916, B2 => 
                           n9892, ZN => n18715);
   U16969 : OAI221_X1 port map( B1 => n16248, B2 => n20860, C1 => n16142, C2 =>
                           n20878, A => n18723, ZN => n18716);
   U16970 : AOI22_X1 port map( A1 => n20957, A2 => n19922, B1 => n20915, B2 => 
                           n9924, ZN => n18723);
   U16971 : OAI221_X1 port map( B1 => n16212, B2 => n20861, C1 => n16106, C2 =>
                           n20875, A => n18678, ZN => n18671);
   U16972 : AOI22_X1 port map( A1 => n20960, A2 => n19923, B1 => n20918, B2 => 
                           n9891, ZN => n18678);
   U16973 : OAI221_X1 port map( B1 => n16247, B2 => n20860, C1 => n16141, C2 =>
                           n20874, A => n18686, ZN => n18679);
   U16974 : AOI22_X1 port map( A1 => n20959, A2 => n19924, B1 => n20917, B2 => 
                           n9923, ZN => n18686);
   U16975 : OAI221_X1 port map( B1 => n16211, B2 => n20863, C1 => n16105, C2 =>
                           n20876, A => n18641, ZN => n18634);
   U16976 : AOI22_X1 port map( A1 => n20962, A2 => n19925, B1 => n20920, B2 => 
                           n9890, ZN => n18641);
   U16977 : OAI221_X1 port map( B1 => n16246, B2 => n20862, C1 => n16140, C2 =>
                           n20875, A => n18649, ZN => n18642);
   U16978 : AOI22_X1 port map( A1 => n20961, A2 => n19926, B1 => n20919, B2 => 
                           n9922, ZN => n18649);
   U16979 : OAI221_X1 port map( B1 => n16210, B2 => n20859, C1 => n16104, C2 =>
                           n20878, A => n18604, ZN => n18597);
   U16980 : AOI22_X1 port map( A1 => n20964, A2 => n19927, B1 => n20922, B2 => 
                           n9889, ZN => n18604);
   U16981 : OAI221_X1 port map( B1 => n16245, B2 => n20864, C1 => n16139, C2 =>
                           n20877, A => n18612, ZN => n18605);
   U16982 : AOI22_X1 port map( A1 => n20963, A2 => n19928, B1 => n20921, B2 => 
                           n9921, ZN => n18612);
   U16983 : OAI221_X1 port map( B1 => n16209, B2 => n20862, C1 => n16103, C2 =>
                           n20876, A => n18567, ZN => n18560);
   U16984 : AOI22_X1 port map( A1 => n20964, A2 => n19929, B1 => n20924, B2 => 
                           n9888, ZN => n18567);
   U16985 : OAI221_X1 port map( B1 => n16244, B2 => n20861, C1 => n16138, C2 =>
                           n20873, A => n18575, ZN => n18568);
   U16986 : AOI22_X1 port map( A1 => n20976, A2 => n19930, B1 => n20923, B2 => 
                           n9920, ZN => n18575);
   U16987 : OAI221_X1 port map( B1 => n16208, B2 => n20861, C1 => n16102, C2 =>
                           n20875, A => n18530, ZN => n18523);
   U16988 : AOI22_X1 port map( A1 => n20969, A2 => n19931, B1 => n20928, B2 => 
                           n9887, ZN => n18530);
   U16989 : OAI221_X1 port map( B1 => n16243, B2 => n20860, C1 => n16137, C2 =>
                           n20874, A => n18538, ZN => n18531);
   U16990 : AOI22_X1 port map( A1 => n20969, A2 => n19932, B1 => n20928, B2 => 
                           n9919, ZN => n18538);
   U16991 : OAI221_X1 port map( B1 => n16207, B2 => n20863, C1 => n16101, C2 =>
                           n20877, A => n18479, ZN => n18458);
   U16992 : AOI22_X1 port map( A1 => n20971, A2 => n19933, B1 => n20930, B2 => 
                           n9886, ZN => n18479);
   U16993 : OAI221_X1 port map( B1 => n16242, B2 => n20862, C1 => n16136, C2 =>
                           n20876, A => n18489, ZN => n18482);
   U16994 : AOI22_X1 port map( A1 => n20969, A2 => n19934, B1 => n20928, B2 => 
                           n9918, ZN => n18489);
   U16995 : OAI221_X1 port map( B1 => n16238, B2 => n21420, C1 => n16132, C2 =>
                           n21430, A => n18385, ZN => n18376);
   U16996 : AOI22_X1 port map( A1 => n21509, A2 => n19875, B1 => n21467, B2 => 
                           n9917, ZN => n18385);
   U16997 : OAI221_X1 port map( B1 => n16273, B2 => n21419, C1 => n16167, C2 =>
                           n21435, A => n18403, ZN => n18387);
   U16998 : AOI22_X1 port map( A1 => n21508, A2 => n19876, B1 => n21466, B2 => 
                           n9949, ZN => n18403);
   U16999 : OAI221_X1 port map( B1 => n16237, B2 => n21416, C1 => n16131, C2 =>
                           n21432, A => n18324, ZN => n18315);
   U17000 : AOI22_X1 port map( A1 => n21511, A2 => n19877, B1 => n21469, B2 => 
                           n9916, ZN => n18324);
   U17001 : OAI221_X1 port map( B1 => n16272, B2 => n21421, C1 => n16166, C2 =>
                           n21431, A => n18335, ZN => n18326);
   U17002 : AOI22_X1 port map( A1 => n21510, A2 => n19878, B1 => n21468, B2 => 
                           n9948, ZN => n18335);
   U17003 : OAI221_X1 port map( B1 => n16236, B2 => n21416, C1 => n16130, C2 =>
                           n21430, A => n18277, ZN => n18268);
   U17004 : AOI22_X1 port map( A1 => n21513, A2 => n19879, B1 => n21471, B2 => 
                           n9915, ZN => n18277);
   U17005 : OAI221_X1 port map( B1 => n16271, B2 => n21421, C1 => n16165, C2 =>
                           n21433, A => n18288, ZN => n18279);
   U17006 : AOI22_X1 port map( A1 => n21512, A2 => n19880, B1 => n21470, B2 => 
                           n9947, ZN => n18288);
   U17007 : OAI221_X1 port map( B1 => n16235, B2 => n21418, C1 => n16129, C2 =>
                           n21435, A => n18230, ZN => n18221);
   U17008 : AOI22_X1 port map( A1 => n21515, A2 => n19881, B1 => n21473, B2 => 
                           n9914, ZN => n18230);
   U17009 : OAI221_X1 port map( B1 => n16270, B2 => n21417, C1 => n16164, C2 =>
                           n21434, A => n18241, ZN => n18232);
   U17010 : AOI22_X1 port map( A1 => n21514, A2 => n19882, B1 => n21472, B2 => 
                           n9946, ZN => n18241);
   U17011 : OAI221_X1 port map( B1 => n16234, B2 => n21420, C1 => n16128, C2 =>
                           n21431, A => n18183, ZN => n18174);
   U17012 : AOI22_X1 port map( A1 => n21517, A2 => n19883, B1 => n21475, B2 => 
                           n9913, ZN => n18183);
   U17013 : OAI221_X1 port map( B1 => n16269, B2 => n21419, C1 => n16163, C2 =>
                           n21430, A => n18194, ZN => n18185);
   U17014 : AOI22_X1 port map( A1 => n21516, A2 => n19884, B1 => n21474, B2 => 
                           n9945, ZN => n18194);
   U17015 : OAI221_X1 port map( B1 => n16233, B2 => n21417, C1 => n16127, C2 =>
                           n21431, A => n18136, ZN => n18127);
   U17016 : AOI22_X1 port map( A1 => n21519, A2 => n19885, B1 => n21477, B2 => 
                           n9912, ZN => n18136);
   U17017 : OAI221_X1 port map( B1 => n16268, B2 => n21416, C1 => n16162, C2 =>
                           n21432, A => n18147, ZN => n18138);
   U17018 : AOI22_X1 port map( A1 => n21518, A2 => n19886, B1 => n21476, B2 => 
                           n9944, ZN => n18147);
   U17019 : OAI221_X1 port map( B1 => n16232, B2 => n21416, C1 => n16126, C2 =>
                           n21434, A => n18089, ZN => n18080);
   U17020 : AOI22_X1 port map( A1 => n21521, A2 => n19887, B1 => n21479, B2 => 
                           n9911, ZN => n18089);
   U17021 : OAI221_X1 port map( B1 => n16267, B2 => n21421, C1 => n16161, C2 =>
                           n21433, A => n18100, ZN => n18091);
   U17022 : AOI22_X1 port map( A1 => n21520, A2 => n19888, B1 => n21478, B2 => 
                           n9943, ZN => n18100);
   U17023 : OAI221_X1 port map( B1 => n16231, B2 => n21418, C1 => n16125, C2 =>
                           n21430, A => n18042, ZN => n18033);
   U17024 : AOI22_X1 port map( A1 => n21521, A2 => n19889, B1 => n21481, B2 => 
                           n9910, ZN => n18042);
   U17025 : OAI221_X1 port map( B1 => n16266, B2 => n21417, C1 => n16160, C2 =>
                           n21435, A => n18053, ZN => n18044);
   U17026 : AOI22_X1 port map( A1 => n21534, A2 => n19890, B1 => n21480, B2 => 
                           n9942, ZN => n18053);
   U17027 : OAI221_X1 port map( B1 => n16230, B2 => n21418, C1 => n16124, C2 =>
                           n21432, A => n17995, ZN => n17986);
   U17028 : AOI22_X1 port map( A1 => n21526, A2 => n19891, B1 => n21485, B2 => 
                           n9909, ZN => n17995);
   U17029 : OAI221_X1 port map( B1 => n16265, B2 => n21417, C1 => n16159, C2 =>
                           n21431, A => n18006, ZN => n17997);
   U17030 : AOI22_X1 port map( A1 => n21526, A2 => n19892, B1 => n21485, B2 => 
                           n9941, ZN => n18006);
   U17031 : OAI221_X1 port map( B1 => n16229, B2 => n21420, C1 => n16123, C2 =>
                           n21433, A => n17948, ZN => n17939);
   U17032 : AOI22_X1 port map( A1 => n21527, A2 => n19893, B1 => n21486, B2 => 
                           n9908, ZN => n17948);
   U17033 : OAI221_X1 port map( B1 => n16264, B2 => n21419, C1 => n16158, C2 =>
                           n21432, A => n17959, ZN => n17950);
   U17034 : AOI22_X1 port map( A1 => n21526, A2 => n19894, B1 => n21485, B2 => 
                           n9940, ZN => n17959);
   U17035 : OAI221_X1 port map( B1 => n16228, B2 => n21416, C1 => n16122, C2 =>
                           n21435, A => n17901, ZN => n17892);
   U17036 : AOI22_X1 port map( A1 => n21528, A2 => n19895, B1 => n21487, B2 => 
                           n9907, ZN => n17901);
   U17037 : OAI221_X1 port map( B1 => n16263, B2 => n21421, C1 => n16157, C2 =>
                           n21434, A => n17912, ZN => n17903);
   U17038 : AOI22_X1 port map( A1 => n21527, A2 => n19896, B1 => n21486, B2 => 
                           n9939, ZN => n17912);
   U17039 : OAI221_X1 port map( B1 => n16227, B2 => n21419, C1 => n16121, C2 =>
                           n21433, A => n17854, ZN => n17845);
   U17040 : AOI22_X1 port map( A1 => n21529, A2 => n19897, B1 => n21488, B2 => 
                           n9906, ZN => n17854);
   U17041 : OAI221_X1 port map( B1 => n16262, B2 => n21418, C1 => n16156, C2 =>
                           n21430, A => n17865, ZN => n17856);
   U17042 : AOI22_X1 port map( A1 => n21530, A2 => n19898, B1 => n21488, B2 => 
                           n9938, ZN => n17865);
   U17043 : OAI221_X1 port map( B1 => n16226, B2 => n21418, C1 => n16120, C2 =>
                           n21432, A => n17807, ZN => n17798);
   U17044 : AOI22_X1 port map( A1 => n21531, A2 => n19899, B1 => n21489, B2 => 
                           n9905, ZN => n17807);
   U17045 : OAI221_X1 port map( B1 => n16261, B2 => n21417, C1 => n16155, C2 =>
                           n21431, A => n17818, ZN => n17809);
   U17046 : AOI22_X1 port map( A1 => n21530, A2 => n19900, B1 => n21488, B2 => 
                           n9937, ZN => n17818);
   U17047 : OAI221_X1 port map( B1 => n16225, B2 => n21420, C1 => n16119, C2 =>
                           n21434, A => n17760, ZN => n17751);
   U17048 : AOI22_X1 port map( A1 => n21532, A2 => n19901, B1 => n21490, B2 => 
                           n9904, ZN => n17760);
   U17049 : OAI221_X1 port map( B1 => n16260, B2 => n21419, C1 => n16154, C2 =>
                           n21433, A => n17771, ZN => n17762);
   U17050 : AOI22_X1 port map( A1 => n21532, A2 => n19902, B1 => n21490, B2 => 
                           n9936, ZN => n17771);
   U17051 : OAI221_X1 port map( B1 => n16224, B2 => n21420, C1 => n16118, C2 =>
                           n21434, A => n17713, ZN => n17704);
   U17052 : AOI22_X1 port map( A1 => n21528, A2 => n19903, B1 => n21487, B2 => 
                           n9903, ZN => n17713);
   U17053 : OAI221_X1 port map( B1 => n16259, B2 => n21419, C1 => n16153, C2 =>
                           n21435, A => n17724, ZN => n17715);
   U17054 : AOI22_X1 port map( A1 => n21530, A2 => n19904, B1 => n21492, B2 => 
                           n9935, ZN => n17724);
   U17055 : OAI221_X1 port map( B1 => n16223, B2 => n21416, C1 => n16117, C2 =>
                           n21431, A => n17666, ZN => n17657);
   U17056 : AOI22_X1 port map( A1 => n21529, A2 => n19905, B1 => n21488, B2 => 
                           n9902, ZN => n17666);
   U17057 : OAI221_X1 port map( B1 => n16258, B2 => n21421, C1 => n16152, C2 =>
                           n21430, A => n17677, ZN => n17668);
   U17058 : AOI22_X1 port map( A1 => n21530, A2 => n19906, B1 => n21488, B2 => 
                           n9934, ZN => n17677);
   U17059 : OAI221_X1 port map( B1 => n16222, B2 => n21418, C1 => n16116, C2 =>
                           n21433, A => n17619, ZN => n17610);
   U17060 : AOI22_X1 port map( A1 => n21531, A2 => n19907, B1 => n21489, B2 => 
                           n9901, ZN => n17619);
   U17061 : OAI221_X1 port map( B1 => n16257, B2 => n21417, C1 => n16151, C2 =>
                           n21432, A => n17630, ZN => n17621);
   U17062 : AOI22_X1 port map( A1 => n21530, A2 => n19908, B1 => n21488, B2 => 
                           n9933, ZN => n17630);
   U17063 : OAI221_X1 port map( B1 => n16221, B2 => n21421, C1 => n16115, C2 =>
                           n21435, A => n17572, ZN => n17563);
   U17064 : AOI22_X1 port map( A1 => n21527, A2 => n19909, B1 => n21486, B2 => 
                           n9900, ZN => n17572);
   U17065 : OAI221_X1 port map( B1 => n16256, B2 => n21420, C1 => n16150, C2 =>
                           n21434, A => n17583, ZN => n17574);
   U17066 : AOI22_X1 port map( A1 => n21532, A2 => n19910, B1 => n21490, B2 => 
                           n9932, ZN => n17583);
   U17067 : OAI221_X1 port map( B1 => n16255, B2 => n21419, C1 => n16149, C2 =>
                           n21435, A => n17536, ZN => n17527);
   U17068 : AOI22_X1 port map( A1 => n21533, A2 => n19911, B1 => n21491, B2 => 
                           n9931, ZN => n17536);
   U17069 : OAI221_X1 port map( B1 => n16254, B2 => n21421, C1 => n16148, C2 =>
                           n21431, A => n17489, ZN => n17480);
   U17070 : AOI22_X1 port map( A1 => n21534, A2 => n19912, B1 => n21491, B2 => 
                           n9930, ZN => n17489);
   U17071 : OAI221_X1 port map( B1 => n16253, B2 => n21421, C1 => n16147, C2 =>
                           n21433, A => n17442, ZN => n17433);
   U17072 : AOI22_X1 port map( A1 => n21534, A2 => n19913, B1 => n21492, B2 => 
                           n9929, ZN => n17442);
   U17073 : OAI221_X1 port map( B1 => n16252, B2 => n21417, C1 => n16146, C2 =>
                           n21434, A => n17395, ZN => n17386);
   U17074 : AOI22_X1 port map( A1 => n21529, A2 => n19914, B1 => n21466, B2 => 
                           n9928, ZN => n17395);
   U17075 : OAI221_X1 port map( B1 => n16216, B2 => n21420, C1 => n16110, C2 =>
                           n21431, A => n17337, ZN => n17328);
   U17076 : AOI22_X1 port map( A1 => n21509, A2 => n19915, B1 => n21467, B2 => 
                           n9895, ZN => n17337);
   U17077 : OAI221_X1 port map( B1 => n16251, B2 => n21419, C1 => n16145, C2 =>
                           n21430, A => n17348, ZN => n17339);
   U17078 : AOI22_X1 port map( A1 => n21508, A2 => n19916, B1 => n21491, B2 => 
                           n9927, ZN => n17348);
   U17079 : OAI221_X1 port map( B1 => n16215, B2 => n21417, C1 => n16109, C2 =>
                           n21431, A => n17290, ZN => n17281);
   U17080 : AOI22_X1 port map( A1 => n21511, A2 => n19917, B1 => n21469, B2 => 
                           n9894, ZN => n17290);
   U17081 : OAI221_X1 port map( B1 => n16250, B2 => n21416, C1 => n16144, C2 =>
                           n21432, A => n17301, ZN => n17292);
   U17082 : AOI22_X1 port map( A1 => n21510, A2 => n19918, B1 => n21468, B2 => 
                           n9926, ZN => n17301);
   U17083 : OAI221_X1 port map( B1 => n16214, B2 => n21416, C1 => n16108, C2 =>
                           n21434, A => n17243, ZN => n17234);
   U17084 : AOI22_X1 port map( A1 => n21513, A2 => n19919, B1 => n21471, B2 => 
                           n9893, ZN => n17243);
   U17085 : OAI221_X1 port map( B1 => n16249, B2 => n21421, C1 => n16143, C2 =>
                           n21433, A => n17254, ZN => n17245);
   U17086 : AOI22_X1 port map( A1 => n21512, A2 => n19920, B1 => n21470, B2 => 
                           n9925, ZN => n17254);
   U17087 : OAI221_X1 port map( B1 => n16213, B2 => n21418, C1 => n16107, C2 =>
                           n21430, A => n17196, ZN => n17187);
   U17088 : AOI22_X1 port map( A1 => n21515, A2 => n19921, B1 => n21473, B2 => 
                           n9892, ZN => n17196);
   U17089 : OAI221_X1 port map( B1 => n16248, B2 => n21417, C1 => n16142, C2 =>
                           n21435, A => n17207, ZN => n17198);
   U17090 : AOI22_X1 port map( A1 => n21514, A2 => n19922, B1 => n21472, B2 => 
                           n9924, ZN => n17207);
   U17091 : OAI221_X1 port map( B1 => n16212, B2 => n21418, C1 => n16106, C2 =>
                           n21432, A => n17149, ZN => n17140);
   U17092 : AOI22_X1 port map( A1 => n21517, A2 => n19923, B1 => n21475, B2 => 
                           n9891, ZN => n17149);
   U17093 : OAI221_X1 port map( B1 => n16247, B2 => n21417, C1 => n16141, C2 =>
                           n21431, A => n17160, ZN => n17151);
   U17094 : AOI22_X1 port map( A1 => n21516, A2 => n19924, B1 => n21474, B2 => 
                           n9923, ZN => n17160);
   U17095 : OAI221_X1 port map( B1 => n16211, B2 => n21420, C1 => n16105, C2 =>
                           n21433, A => n17102, ZN => n17093);
   U17096 : AOI22_X1 port map( A1 => n21519, A2 => n19925, B1 => n21477, B2 => 
                           n9890, ZN => n17102);
   U17097 : OAI221_X1 port map( B1 => n16246, B2 => n21419, C1 => n16140, C2 =>
                           n21432, A => n17113, ZN => n17104);
   U17098 : AOI22_X1 port map( A1 => n21518, A2 => n19926, B1 => n21476, B2 => 
                           n9922, ZN => n17113);
   U17099 : OAI221_X1 port map( B1 => n16210, B2 => n21416, C1 => n16104, C2 =>
                           n21435, A => n17055, ZN => n17046);
   U17100 : AOI22_X1 port map( A1 => n21521, A2 => n19927, B1 => n21479, B2 => 
                           n9889, ZN => n17055);
   U17101 : OAI221_X1 port map( B1 => n16245, B2 => n21421, C1 => n16139, C2 =>
                           n21434, A => n17066, ZN => n17057);
   U17102 : AOI22_X1 port map( A1 => n21520, A2 => n19928, B1 => n21478, B2 => 
                           n9921, ZN => n17066);
   U17103 : OAI221_X1 port map( B1 => n16209, B2 => n21419, C1 => n16103, C2 =>
                           n21433, A => n17008, ZN => n16999);
   U17104 : AOI22_X1 port map( A1 => n21521, A2 => n19929, B1 => n21481, B2 => 
                           n9888, ZN => n17008);
   U17105 : OAI221_X1 port map( B1 => n16244, B2 => n21418, C1 => n16138, C2 =>
                           n21430, A => n17019, ZN => n17010);
   U17106 : AOI22_X1 port map( A1 => n21533, A2 => n19930, B1 => n21480, B2 => 
                           n9920, ZN => n17019);
   U17107 : OAI221_X1 port map( B1 => n16208, B2 => n21418, C1 => n16102, C2 =>
                           n21432, A => n16961, ZN => n16952);
   U17108 : AOI22_X1 port map( A1 => n21526, A2 => n19931, B1 => n21485, B2 => 
                           n9887, ZN => n16961);
   U17109 : OAI221_X1 port map( B1 => n16243, B2 => n21417, C1 => n16137, C2 =>
                           n21431, A => n16972, ZN => n16963);
   U17110 : AOI22_X1 port map( A1 => n21526, A2 => n19932, B1 => n21485, B2 => 
                           n9919, ZN => n16972);
   U17111 : OAI221_X1 port map( B1 => n16207, B2 => n21420, C1 => n16101, C2 =>
                           n21434, A => n16900, ZN => n16877);
   U17112 : AOI22_X1 port map( A1 => n21528, A2 => n19933, B1 => n21487, B2 => 
                           n9886, ZN => n16900);
   U17113 : OAI221_X1 port map( B1 => n16242, B2 => n21419, C1 => n16136, C2 =>
                           n21433, A => n16913, ZN => n16904);
   U17114 : AOI22_X1 port map( A1 => n21526, A2 => n19934, B1 => n21485, B2 => 
                           n9918, ZN => n16913);
   U17115 : INV_X1 port map( A => ADD_RD1(1), ZN => n19645);
   U17116 : INV_X1 port map( A => ADD_RD2(1), ZN => n18374);
   U17117 : NAND2_X1 port map( A1 => n19667, A2 => ADD_RD1(2), ZN => n18468);
   U17118 : NAND2_X1 port map( A1 => n18401, A2 => ADD_RD2(2), ZN => n16888);
   U17119 : NAND2_X1 port map( A1 => n19678, A2 => ADD_RD1(2), ZN => n18472);
   U17120 : NAND2_X1 port map( A1 => n18415, A2 => ADD_RD2(2), ZN => n16893);
   U17121 : NAND2_X1 port map( A1 => n19660, A2 => ADD_RD1(2), ZN => n18463);
   U17122 : NAND2_X1 port map( A1 => n18393, A2 => ADD_RD2(2), ZN => n16882);
   U17123 : NAND2_X1 port map( A1 => ADD_RD1(2), A2 => n19675, ZN => n18477);
   U17124 : NAND2_X1 port map( A1 => ADD_RD2(2), A2 => n18411, ZN => n16898);
   U17125 : OAI22_X1 port map( A1 => n16756, A2 => n18498, B1 => n4287, B2 => 
                           n18499, ZN => n19676);
   U17126 : OAI22_X1 port map( A1 => n15607, A2 => n18503, B1 => n4350, B2 => 
                           n18504, ZN => n19679);
   U17127 : OAI22_X1 port map( A1 => n16756, A2 => n16925, B1 => n4287, B2 => 
                           n16926, ZN => n18413);
   U17128 : OAI22_X1 port map( A1 => n15607, A2 => n16930, B1 => n4350, B2 => 
                           n16931, ZN => n18416);
   U17129 : NAND2_X1 port map( A1 => DATAIN(0), A2 => n22373, ZN => n15150);
   U17130 : NAND2_X1 port map( A1 => DATAIN(1), A2 => n22373, ZN => n15149);
   U17131 : NAND2_X1 port map( A1 => DATAIN(2), A2 => n22373, ZN => n15148);
   U17132 : NAND2_X1 port map( A1 => DATAIN(3), A2 => n22373, ZN => n15147);
   U17133 : NAND2_X1 port map( A1 => DATAIN(4), A2 => n22373, ZN => n15146);
   U17134 : NAND2_X1 port map( A1 => DATAIN(5), A2 => n22373, ZN => n15145);
   U17135 : NAND2_X1 port map( A1 => DATAIN(6), A2 => n22373, ZN => n15144);
   U17136 : NAND2_X1 port map( A1 => DATAIN(7), A2 => n22373, ZN => n15143);
   U17137 : NAND2_X1 port map( A1 => DATAIN(8), A2 => n22373, ZN => n15142);
   U17138 : NAND2_X1 port map( A1 => DATAIN(9), A2 => n22373, ZN => n15141);
   U17139 : NAND2_X1 port map( A1 => DATAIN(10), A2 => n22373, ZN => n15140);
   U17140 : NAND2_X1 port map( A1 => DATAIN(11), A2 => n22373, ZN => n15139);
   U17141 : NAND2_X1 port map( A1 => DATAIN(12), A2 => n22374, ZN => n15138);
   U17142 : NAND2_X1 port map( A1 => DATAIN(13), A2 => n22374, ZN => n15137);
   U17143 : NAND2_X1 port map( A1 => DATAIN(14), A2 => n22374, ZN => n15136);
   U17144 : NAND2_X1 port map( A1 => DATAIN(15), A2 => n22374, ZN => n15135);
   U17145 : NAND2_X1 port map( A1 => DATAIN(16), A2 => n22374, ZN => n15134);
   U17146 : NAND2_X1 port map( A1 => DATAIN(17), A2 => n22374, ZN => n15133);
   U17147 : NAND2_X1 port map( A1 => DATAIN(18), A2 => n22374, ZN => n15132);
   U17148 : NAND2_X1 port map( A1 => DATAIN(19), A2 => n22374, ZN => n15131);
   U17149 : NAND2_X1 port map( A1 => DATAIN(20), A2 => n22374, ZN => n15130);
   U17150 : NAND2_X1 port map( A1 => DATAIN(21), A2 => n22374, ZN => n15129);
   U17151 : NAND2_X1 port map( A1 => DATAIN(22), A2 => n22374, ZN => n15128);
   U17152 : NAND2_X1 port map( A1 => DATAIN(23), A2 => n22374, ZN => n15127);
   U17153 : NAND2_X1 port map( A1 => DATAIN(24), A2 => n22375, ZN => n15126);
   U17154 : NAND2_X1 port map( A1 => DATAIN(25), A2 => n22375, ZN => n15125);
   U17155 : NAND2_X1 port map( A1 => DATAIN(26), A2 => n22375, ZN => n15124);
   U17156 : NAND2_X1 port map( A1 => DATAIN(27), A2 => n22375, ZN => n15123);
   U17157 : NAND2_X1 port map( A1 => DATAIN(28), A2 => n22375, ZN => n15122);
   U17158 : NAND2_X1 port map( A1 => DATAIN(29), A2 => n22375, ZN => n15121);
   U17159 : NAND2_X1 port map( A1 => DATAIN(30), A2 => n22375, ZN => n15120);
   U17160 : NAND2_X1 port map( A1 => DATAIN(31), A2 => n22375, ZN => n15118);
   U17161 : OAI22_X1 port map( A1 => n21826, A2 => n22530, B1 => n16797, B2 => 
                           n16805, ZN => n5494);
   U17162 : OAI22_X1 port map( A1 => n21827, A2 => n22536, B1 => n16797, B2 => 
                           n16804, ZN => n5495);
   U17163 : OAI22_X1 port map( A1 => n21827, A2 => n22542, B1 => n16797, B2 => 
                           n16803, ZN => n5496);
   U17164 : OAI22_X1 port map( A1 => n21827, A2 => n22548, B1 => n21821, B2 => 
                           n16802, ZN => n5497);
   U17165 : OAI22_X1 port map( A1 => n21827, A2 => n22554, B1 => n21821, B2 => 
                           n16801, ZN => n5498);
   U17166 : OAI22_X1 port map( A1 => n21827, A2 => n22560, B1 => n21821, B2 => 
                           n16800, ZN => n5499);
   U17167 : OAI22_X1 port map( A1 => n21828, A2 => n22566, B1 => n21821, B2 => 
                           n16799, ZN => n5500);
   U17168 : OAI22_X1 port map( A1 => n21828, A2 => n22581, B1 => n16797, B2 => 
                           n16798, ZN => n5501);
   U17169 : OAI22_X1 port map( A1 => n21835, A2 => n22530, B1 => n16760, B2 => 
                           n16768, ZN => n5526);
   U17170 : OAI22_X1 port map( A1 => n21836, A2 => n22536, B1 => n16760, B2 => 
                           n16767, ZN => n5527);
   U17171 : OAI22_X1 port map( A1 => n21836, A2 => n22542, B1 => n16760, B2 => 
                           n16766, ZN => n5528);
   U17172 : OAI22_X1 port map( A1 => n21836, A2 => n22548, B1 => n21830, B2 => 
                           n16765, ZN => n5529);
   U17173 : OAI22_X1 port map( A1 => n21836, A2 => n22554, B1 => n21830, B2 => 
                           n16764, ZN => n5530);
   U17174 : OAI22_X1 port map( A1 => n21836, A2 => n22560, B1 => n21830, B2 => 
                           n16763, ZN => n5531);
   U17175 : OAI22_X1 port map( A1 => n21837, A2 => n22566, B1 => n21830, B2 => 
                           n16762, ZN => n5532);
   U17176 : OAI22_X1 port map( A1 => n21837, A2 => n22581, B1 => n16760, B2 => 
                           n16761, ZN => n5533);
   U17177 : OAI22_X1 port map( A1 => n21862, A2 => n22529, B1 => n16690, B2 => 
                           n16698, ZN => n5622);
   U17178 : OAI22_X1 port map( A1 => n21863, A2 => n22535, B1 => n16690, B2 => 
                           n16697, ZN => n5623);
   U17179 : OAI22_X1 port map( A1 => n21863, A2 => n22541, B1 => n16690, B2 => 
                           n16696, ZN => n5624);
   U17180 : OAI22_X1 port map( A1 => n21863, A2 => n22547, B1 => n21857, B2 => 
                           n16695, ZN => n5625);
   U17181 : OAI22_X1 port map( A1 => n21863, A2 => n22553, B1 => n21857, B2 => 
                           n16694, ZN => n5626);
   U17182 : OAI22_X1 port map( A1 => n21863, A2 => n22559, B1 => n21857, B2 => 
                           n16693, ZN => n5627);
   U17183 : OAI22_X1 port map( A1 => n21864, A2 => n22565, B1 => n21857, B2 => 
                           n16692, ZN => n5628);
   U17184 : OAI22_X1 port map( A1 => n21864, A2 => n22580, B1 => n16690, B2 => 
                           n16691, ZN => n5629);
   U17185 : OAI22_X1 port map( A1 => n21871, A2 => n22529, B1 => n16655, B2 => 
                           n16663, ZN => n5654);
   U17186 : OAI22_X1 port map( A1 => n21872, A2 => n22535, B1 => n16655, B2 => 
                           n16662, ZN => n5655);
   U17187 : OAI22_X1 port map( A1 => n21872, A2 => n22541, B1 => n16655, B2 => 
                           n16661, ZN => n5656);
   U17188 : OAI22_X1 port map( A1 => n21872, A2 => n22547, B1 => n21866, B2 => 
                           n16660, ZN => n5657);
   U17189 : OAI22_X1 port map( A1 => n21872, A2 => n22553, B1 => n21866, B2 => 
                           n16659, ZN => n5658);
   U17190 : OAI22_X1 port map( A1 => n21872, A2 => n22559, B1 => n21866, B2 => 
                           n16658, ZN => n5659);
   U17191 : OAI22_X1 port map( A1 => n21873, A2 => n22565, B1 => n21866, B2 => 
                           n16657, ZN => n5660);
   U17192 : OAI22_X1 port map( A1 => n21873, A2 => n22580, B1 => n16655, B2 => 
                           n16656, ZN => n5661);
   U17193 : OAI22_X1 port map( A1 => n21880, A2 => n22529, B1 => n16620, B2 => 
                           n16628, ZN => n5686);
   U17194 : OAI22_X1 port map( A1 => n21881, A2 => n22535, B1 => n16620, B2 => 
                           n16627, ZN => n5687);
   U17195 : OAI22_X1 port map( A1 => n21881, A2 => n22541, B1 => n16620, B2 => 
                           n16626, ZN => n5688);
   U17196 : OAI22_X1 port map( A1 => n21881, A2 => n22547, B1 => n21875, B2 => 
                           n16625, ZN => n5689);
   U17197 : OAI22_X1 port map( A1 => n21881, A2 => n22553, B1 => n21875, B2 => 
                           n16624, ZN => n5690);
   U17198 : OAI22_X1 port map( A1 => n21881, A2 => n22559, B1 => n21875, B2 => 
                           n16623, ZN => n5691);
   U17199 : OAI22_X1 port map( A1 => n21882, A2 => n22565, B1 => n21875, B2 => 
                           n16622, ZN => n5692);
   U17200 : OAI22_X1 port map( A1 => n21882, A2 => n22580, B1 => n16620, B2 => 
                           n16621, ZN => n5693);
   U17201 : OAI22_X1 port map( A1 => n21925, A2 => n22529, B1 => n16576, B2 => 
                           n16584, ZN => n5846);
   U17202 : OAI22_X1 port map( A1 => n21926, A2 => n22535, B1 => n16576, B2 => 
                           n16583, ZN => n5847);
   U17203 : OAI22_X1 port map( A1 => n21926, A2 => n22541, B1 => n16576, B2 => 
                           n16582, ZN => n5848);
   U17204 : OAI22_X1 port map( A1 => n21926, A2 => n22547, B1 => n21920, B2 => 
                           n16581, ZN => n5849);
   U17205 : OAI22_X1 port map( A1 => n21926, A2 => n22553, B1 => n21920, B2 => 
                           n16580, ZN => n5850);
   U17206 : OAI22_X1 port map( A1 => n21926, A2 => n22559, B1 => n21920, B2 => 
                           n16579, ZN => n5851);
   U17207 : OAI22_X1 port map( A1 => n21927, A2 => n22565, B1 => n21920, B2 => 
                           n16578, ZN => n5852);
   U17208 : OAI22_X1 port map( A1 => n21927, A2 => n22580, B1 => n16576, B2 => 
                           n16577, ZN => n5853);
   U17209 : OAI22_X1 port map( A1 => n21961, A2 => n22528, B1 => n16453, B2 => 
                           n16461, ZN => n5974);
   U17210 : OAI22_X1 port map( A1 => n21962, A2 => n22534, B1 => n16453, B2 => 
                           n16460, ZN => n5975);
   U17211 : OAI22_X1 port map( A1 => n21962, A2 => n22540, B1 => n16453, B2 => 
                           n16459, ZN => n5976);
   U17212 : OAI22_X1 port map( A1 => n21962, A2 => n22546, B1 => n21956, B2 => 
                           n16458, ZN => n5977);
   U17213 : OAI22_X1 port map( A1 => n21962, A2 => n22552, B1 => n21956, B2 => 
                           n16457, ZN => n5978);
   U17214 : OAI22_X1 port map( A1 => n21962, A2 => n22558, B1 => n21956, B2 => 
                           n16456, ZN => n5979);
   U17215 : OAI22_X1 port map( A1 => n21963, A2 => n22564, B1 => n21956, B2 => 
                           n16455, ZN => n5980);
   U17216 : OAI22_X1 port map( A1 => n21963, A2 => n22579, B1 => n16453, B2 => 
                           n16454, ZN => n5981);
   U17217 : OAI22_X1 port map( A1 => n21970, A2 => n22528, B1 => n16419, B2 => 
                           n16427, ZN => n6006);
   U17218 : OAI22_X1 port map( A1 => n21971, A2 => n22534, B1 => n16419, B2 => 
                           n16426, ZN => n6007);
   U17219 : OAI22_X1 port map( A1 => n21971, A2 => n22540, B1 => n16419, B2 => 
                           n16425, ZN => n6008);
   U17220 : OAI22_X1 port map( A1 => n21971, A2 => n22546, B1 => n21965, B2 => 
                           n16424, ZN => n6009);
   U17221 : OAI22_X1 port map( A1 => n21971, A2 => n22552, B1 => n21965, B2 => 
                           n16423, ZN => n6010);
   U17222 : OAI22_X1 port map( A1 => n21971, A2 => n22558, B1 => n21965, B2 => 
                           n16422, ZN => n6011);
   U17223 : OAI22_X1 port map( A1 => n21972, A2 => n22564, B1 => n21965, B2 => 
                           n16421, ZN => n6012);
   U17224 : OAI22_X1 port map( A1 => n21972, A2 => n22579, B1 => n16419, B2 => 
                           n16420, ZN => n6013);
   U17225 : OAI22_X1 port map( A1 => n21979, A2 => n22528, B1 => n16384, B2 => 
                           n16392, ZN => n6038);
   U17226 : OAI22_X1 port map( A1 => n21980, A2 => n22534, B1 => n16384, B2 => 
                           n16391, ZN => n6039);
   U17227 : OAI22_X1 port map( A1 => n21980, A2 => n22540, B1 => n16384, B2 => 
                           n16390, ZN => n6040);
   U17228 : OAI22_X1 port map( A1 => n21980, A2 => n22546, B1 => n21974, B2 => 
                           n16389, ZN => n6041);
   U17229 : OAI22_X1 port map( A1 => n21980, A2 => n22552, B1 => n21974, B2 => 
                           n16388, ZN => n6042);
   U17230 : OAI22_X1 port map( A1 => n21980, A2 => n22558, B1 => n21974, B2 => 
                           n16387, ZN => n6043);
   U17231 : OAI22_X1 port map( A1 => n21981, A2 => n22564, B1 => n21974, B2 => 
                           n16386, ZN => n6044);
   U17232 : OAI22_X1 port map( A1 => n21981, A2 => n22579, B1 => n16384, B2 => 
                           n16385, ZN => n6045);
   U17233 : OAI22_X1 port map( A1 => n22033, A2 => n22528, B1 => n16275, B2 => 
                           n16283, ZN => n6230);
   U17234 : OAI22_X1 port map( A1 => n22034, A2 => n22534, B1 => n16275, B2 => 
                           n16282, ZN => n6231);
   U17235 : OAI22_X1 port map( A1 => n22034, A2 => n22540, B1 => n16275, B2 => 
                           n16281, ZN => n6232);
   U17236 : OAI22_X1 port map( A1 => n22034, A2 => n22546, B1 => n22028, B2 => 
                           n16280, ZN => n6233);
   U17237 : OAI22_X1 port map( A1 => n22034, A2 => n22552, B1 => n22028, B2 => 
                           n16279, ZN => n6234);
   U17238 : OAI22_X1 port map( A1 => n22034, A2 => n22558, B1 => n22028, B2 => 
                           n16278, ZN => n6235);
   U17239 : OAI22_X1 port map( A1 => n22035, A2 => n22564, B1 => n22028, B2 => 
                           n16277, ZN => n6236);
   U17240 : OAI22_X1 port map( A1 => n22035, A2 => n22579, B1 => n16275, B2 => 
                           n16276, ZN => n6237);
   U17241 : OAI22_X1 port map( A1 => n22114, A2 => n22527, B1 => n15998, B2 => 
                           n16006, ZN => n6518);
   U17242 : OAI22_X1 port map( A1 => n22115, A2 => n22533, B1 => n15998, B2 => 
                           n16005, ZN => n6519);
   U17243 : OAI22_X1 port map( A1 => n22115, A2 => n22539, B1 => n15998, B2 => 
                           n16004, ZN => n6520);
   U17244 : OAI22_X1 port map( A1 => n22115, A2 => n22545, B1 => n22109, B2 => 
                           n16003, ZN => n6521);
   U17245 : OAI22_X1 port map( A1 => n22115, A2 => n22551, B1 => n22109, B2 => 
                           n16002, ZN => n6522);
   U17246 : OAI22_X1 port map( A1 => n22115, A2 => n22557, B1 => n22109, B2 => 
                           n16001, ZN => n6523);
   U17247 : OAI22_X1 port map( A1 => n22116, A2 => n22563, B1 => n22109, B2 => 
                           n16000, ZN => n6524);
   U17248 : OAI22_X1 port map( A1 => n22116, A2 => n22578, B1 => n15998, B2 => 
                           n15999, ZN => n6525);
   U17249 : OAI22_X1 port map( A1 => n22123, A2 => n22527, B1 => n15963, B2 => 
                           n15971, ZN => n6550);
   U17250 : OAI22_X1 port map( A1 => n22124, A2 => n22533, B1 => n15963, B2 => 
                           n15970, ZN => n6551);
   U17251 : OAI22_X1 port map( A1 => n22124, A2 => n22539, B1 => n15963, B2 => 
                           n15969, ZN => n6552);
   U17252 : OAI22_X1 port map( A1 => n22124, A2 => n22545, B1 => n22118, B2 => 
                           n15968, ZN => n6553);
   U17253 : OAI22_X1 port map( A1 => n22124, A2 => n22551, B1 => n22118, B2 => 
                           n15967, ZN => n6554);
   U17254 : OAI22_X1 port map( A1 => n22124, A2 => n22557, B1 => n22118, B2 => 
                           n15966, ZN => n6555);
   U17255 : OAI22_X1 port map( A1 => n22125, A2 => n22563, B1 => n22118, B2 => 
                           n15965, ZN => n6556);
   U17256 : OAI22_X1 port map( A1 => n22125, A2 => n22578, B1 => n15963, B2 => 
                           n15964, ZN => n6557);
   U17257 : OAI22_X1 port map( A1 => n22132, A2 => n22527, B1 => n15929, B2 => 
                           n15937, ZN => n6582);
   U17258 : OAI22_X1 port map( A1 => n22133, A2 => n22533, B1 => n15929, B2 => 
                           n15936, ZN => n6583);
   U17259 : OAI22_X1 port map( A1 => n22133, A2 => n22539, B1 => n15929, B2 => 
                           n15935, ZN => n6584);
   U17260 : OAI22_X1 port map( A1 => n22133, A2 => n22545, B1 => n22127, B2 => 
                           n15934, ZN => n6585);
   U17261 : OAI22_X1 port map( A1 => n22133, A2 => n22551, B1 => n22127, B2 => 
                           n15933, ZN => n6586);
   U17262 : OAI22_X1 port map( A1 => n22133, A2 => n22557, B1 => n22127, B2 => 
                           n15932, ZN => n6587);
   U17263 : OAI22_X1 port map( A1 => n22134, A2 => n22563, B1 => n22127, B2 => 
                           n15931, ZN => n6588);
   U17264 : OAI22_X1 port map( A1 => n22134, A2 => n22578, B1 => n15929, B2 => 
                           n15930, ZN => n6589);
   U17265 : OAI22_X1 port map( A1 => n22168, A2 => n22526, B1 => n15856, B2 => 
                           n15864, ZN => n6710);
   U17266 : OAI22_X1 port map( A1 => n22169, A2 => n22532, B1 => n15856, B2 => 
                           n15863, ZN => n6711);
   U17267 : OAI22_X1 port map( A1 => n22169, A2 => n22538, B1 => n15856, B2 => 
                           n15862, ZN => n6712);
   U17268 : OAI22_X1 port map( A1 => n22169, A2 => n22544, B1 => n22163, B2 => 
                           n15861, ZN => n6713);
   U17269 : OAI22_X1 port map( A1 => n22169, A2 => n22550, B1 => n22163, B2 => 
                           n15860, ZN => n6714);
   U17270 : OAI22_X1 port map( A1 => n22169, A2 => n22556, B1 => n22163, B2 => 
                           n15859, ZN => n6715);
   U17271 : OAI22_X1 port map( A1 => n22170, A2 => n22562, B1 => n22163, B2 => 
                           n15858, ZN => n6716);
   U17272 : OAI22_X1 port map( A1 => n22170, A2 => n22577, B1 => n15856, B2 => 
                           n15857, ZN => n6717);
   U17273 : OAI22_X1 port map( A1 => n22213, A2 => n22526, B1 => n15716, B2 => 
                           n15724, ZN => n6870);
   U17274 : OAI22_X1 port map( A1 => n22214, A2 => n22532, B1 => n15716, B2 => 
                           n15723, ZN => n6871);
   U17275 : OAI22_X1 port map( A1 => n22214, A2 => n22538, B1 => n15716, B2 => 
                           n15722, ZN => n6872);
   U17276 : OAI22_X1 port map( A1 => n22214, A2 => n22544, B1 => n22208, B2 => 
                           n15721, ZN => n6873);
   U17277 : OAI22_X1 port map( A1 => n22214, A2 => n22550, B1 => n22208, B2 => 
                           n15720, ZN => n6874);
   U17278 : OAI22_X1 port map( A1 => n22214, A2 => n22556, B1 => n22208, B2 => 
                           n15719, ZN => n6875);
   U17279 : OAI22_X1 port map( A1 => n22215, A2 => n22562, B1 => n22208, B2 => 
                           n15718, ZN => n6876);
   U17280 : OAI22_X1 port map( A1 => n22215, A2 => n22577, B1 => n15716, B2 => 
                           n15717, ZN => n6877);
   U17281 : OAI22_X1 port map( A1 => n22240, A2 => n22526, B1 => n15609, B2 => 
                           n15617, ZN => n6966);
   U17282 : OAI22_X1 port map( A1 => n22241, A2 => n22532, B1 => n15609, B2 => 
                           n15616, ZN => n6967);
   U17283 : OAI22_X1 port map( A1 => n22241, A2 => n22538, B1 => n15609, B2 => 
                           n15615, ZN => n6968);
   U17284 : OAI22_X1 port map( A1 => n22241, A2 => n22544, B1 => n22235, B2 => 
                           n15614, ZN => n6969);
   U17285 : OAI22_X1 port map( A1 => n22241, A2 => n22550, B1 => n22235, B2 => 
                           n15613, ZN => n6970);
   U17286 : OAI22_X1 port map( A1 => n22241, A2 => n22556, B1 => n22235, B2 => 
                           n15612, ZN => n6971);
   U17287 : OAI22_X1 port map( A1 => n22242, A2 => n22562, B1 => n22235, B2 => 
                           n15611, ZN => n6972);
   U17288 : OAI22_X1 port map( A1 => n22242, A2 => n22577, B1 => n15609, B2 => 
                           n15610, ZN => n6973);
   U17289 : OAI22_X1 port map( A1 => n22258, A2 => n22526, B1 => n15541, B2 => 
                           n15549, ZN => n7030);
   U17290 : OAI22_X1 port map( A1 => n22259, A2 => n22532, B1 => n15541, B2 => 
                           n15548, ZN => n7031);
   U17291 : OAI22_X1 port map( A1 => n22259, A2 => n22538, B1 => n15541, B2 => 
                           n15547, ZN => n7032);
   U17292 : OAI22_X1 port map( A1 => n22259, A2 => n22544, B1 => n22253, B2 => 
                           n15546, ZN => n7033);
   U17293 : OAI22_X1 port map( A1 => n22259, A2 => n22550, B1 => n22253, B2 => 
                           n15545, ZN => n7034);
   U17294 : OAI22_X1 port map( A1 => n22259, A2 => n22556, B1 => n22253, B2 => 
                           n15544, ZN => n7035);
   U17295 : OAI22_X1 port map( A1 => n22260, A2 => n22562, B1 => n22253, B2 => 
                           n15543, ZN => n7036);
   U17296 : OAI22_X1 port map( A1 => n22260, A2 => n22577, B1 => n15541, B2 => 
                           n15542, ZN => n7037);
   U17297 : OAI22_X1 port map( A1 => n22267, A2 => n22526, B1 => n15506, B2 => 
                           n15514, ZN => n7062);
   U17298 : OAI22_X1 port map( A1 => n22268, A2 => n22532, B1 => n15506, B2 => 
                           n15513, ZN => n7063);
   U17299 : OAI22_X1 port map( A1 => n22268, A2 => n22538, B1 => n15506, B2 => 
                           n15512, ZN => n7064);
   U17300 : OAI22_X1 port map( A1 => n22268, A2 => n22544, B1 => n22262, B2 => 
                           n15511, ZN => n7065);
   U17301 : OAI22_X1 port map( A1 => n22268, A2 => n22550, B1 => n22262, B2 => 
                           n15510, ZN => n7066);
   U17302 : OAI22_X1 port map( A1 => n22268, A2 => n22556, B1 => n22262, B2 => 
                           n15509, ZN => n7067);
   U17303 : OAI22_X1 port map( A1 => n22269, A2 => n22562, B1 => n22262, B2 => 
                           n15508, ZN => n7068);
   U17304 : OAI22_X1 port map( A1 => n22269, A2 => n22577, B1 => n15506, B2 => 
                           n15507, ZN => n7069);
   U17305 : OAI22_X1 port map( A1 => n22312, A2 => n22525, B1 => n15333, B2 => 
                           n15341, ZN => n7222);
   U17306 : OAI22_X1 port map( A1 => n22313, A2 => n22531, B1 => n15333, B2 => 
                           n15340, ZN => n7223);
   U17307 : OAI22_X1 port map( A1 => n22313, A2 => n22537, B1 => n15333, B2 => 
                           n15339, ZN => n7224);
   U17308 : OAI22_X1 port map( A1 => n22313, A2 => n22543, B1 => n22307, B2 => 
                           n15338, ZN => n7225);
   U17309 : OAI22_X1 port map( A1 => n22313, A2 => n22549, B1 => n22307, B2 => 
                           n15337, ZN => n7226);
   U17310 : OAI22_X1 port map( A1 => n22313, A2 => n22555, B1 => n22307, B2 => 
                           n15336, ZN => n7227);
   U17311 : OAI22_X1 port map( A1 => n22314, A2 => n22561, B1 => n22307, B2 => 
                           n15335, ZN => n7228);
   U17312 : OAI22_X1 port map( A1 => n22314, A2 => n22576, B1 => n15333, B2 => 
                           n15334, ZN => n7229);
   U17313 : OAI22_X1 port map( A1 => n22321, A2 => n22525, B1 => n15299, B2 => 
                           n15307, ZN => n7254);
   U17314 : OAI22_X1 port map( A1 => n22322, A2 => n22531, B1 => n15299, B2 => 
                           n15306, ZN => n7255);
   U17315 : OAI22_X1 port map( A1 => n22322, A2 => n22537, B1 => n15299, B2 => 
                           n15305, ZN => n7256);
   U17316 : OAI22_X1 port map( A1 => n22322, A2 => n22543, B1 => n22316, B2 => 
                           n15304, ZN => n7257);
   U17317 : OAI22_X1 port map( A1 => n22322, A2 => n22549, B1 => n22316, B2 => 
                           n15303, ZN => n7258);
   U17318 : OAI22_X1 port map( A1 => n22322, A2 => n22555, B1 => n22316, B2 => 
                           n15302, ZN => n7259);
   U17319 : OAI22_X1 port map( A1 => n22323, A2 => n22561, B1 => n22316, B2 => 
                           n15301, ZN => n7260);
   U17320 : OAI22_X1 port map( A1 => n22323, A2 => n22576, B1 => n15299, B2 => 
                           n15300, ZN => n7261);
   U17321 : OAI22_X1 port map( A1 => n22348, A2 => n22525, B1 => n15193, B2 => 
                           n15201, ZN => n7350);
   U17322 : OAI22_X1 port map( A1 => n22349, A2 => n22531, B1 => n15193, B2 => 
                           n15200, ZN => n7351);
   U17323 : OAI22_X1 port map( A1 => n22349, A2 => n22537, B1 => n15193, B2 => 
                           n15199, ZN => n7352);
   U17324 : OAI22_X1 port map( A1 => n22349, A2 => n22543, B1 => n22343, B2 => 
                           n15198, ZN => n7353);
   U17325 : OAI22_X1 port map( A1 => n22349, A2 => n22549, B1 => n22343, B2 => 
                           n15197, ZN => n7354);
   U17326 : OAI22_X1 port map( A1 => n22349, A2 => n22555, B1 => n22343, B2 => 
                           n15196, ZN => n7355);
   U17327 : OAI22_X1 port map( A1 => n22350, A2 => n22561, B1 => n22343, B2 => 
                           n15195, ZN => n7356);
   U17328 : OAI22_X1 port map( A1 => n22350, A2 => n22576, B1 => n15193, B2 => 
                           n15194, ZN => n7357);
   U17329 : OAI22_X1 port map( A1 => n22357, A2 => n22525, B1 => n15158, B2 => 
                           n15166, ZN => n7382);
   U17330 : OAI22_X1 port map( A1 => n22358, A2 => n22531, B1 => n15158, B2 => 
                           n15165, ZN => n7383);
   U17331 : OAI22_X1 port map( A1 => n22358, A2 => n22537, B1 => n15158, B2 => 
                           n15164, ZN => n7384);
   U17332 : OAI22_X1 port map( A1 => n22358, A2 => n22543, B1 => n22352, B2 => 
                           n15163, ZN => n7385);
   U17333 : OAI22_X1 port map( A1 => n22358, A2 => n22549, B1 => n22352, B2 => 
                           n15162, ZN => n7386);
   U17334 : OAI22_X1 port map( A1 => n22358, A2 => n22555, B1 => n22352, B2 => 
                           n15161, ZN => n7387);
   U17335 : OAI22_X1 port map( A1 => n22359, A2 => n22561, B1 => n22352, B2 => 
                           n15160, ZN => n7388);
   U17336 : OAI22_X1 port map( A1 => n22359, A2 => n22576, B1 => n15158, B2 => 
                           n15159, ZN => n7389);
   U17337 : OAI22_X1 port map( A1 => n4289, A2 => n21801, B1 => n21809, B2 => 
                           n22392, ZN => n5377);
   U17338 : OAI22_X1 port map( A1 => n4291, A2 => n16832, B1 => n21809, B2 => 
                           n22398, ZN => n5379);
   U17339 : OAI22_X1 port map( A1 => n4293, A2 => n16832, B1 => n21809, B2 => 
                           n22404, ZN => n5381);
   U17340 : OAI22_X1 port map( A1 => n4295, A2 => n21801, B1 => n21808, B2 => 
                           n22410, ZN => n5383);
   U17341 : OAI22_X1 port map( A1 => n4297, A2 => n16832, B1 => n21808, B2 => 
                           n22416, ZN => n5385);
   U17342 : OAI22_X1 port map( A1 => n4299, A2 => n21801, B1 => n21808, B2 => 
                           n22422, ZN => n5387);
   U17343 : OAI22_X1 port map( A1 => n4301, A2 => n16832, B1 => n21808, B2 => 
                           n22428, ZN => n5389);
   U17344 : OAI22_X1 port map( A1 => n4303, A2 => n21801, B1 => n21807, B2 => 
                           n22434, ZN => n5391);
   U17345 : OAI22_X1 port map( A1 => n4305, A2 => n21801, B1 => n21807, B2 => 
                           n22440, ZN => n5393);
   U17346 : OAI22_X1 port map( A1 => n4307, A2 => n21801, B1 => n21807, B2 => 
                           n22446, ZN => n5395);
   U17347 : OAI22_X1 port map( A1 => n4309, A2 => n21801, B1 => n21807, B2 => 
                           n22452, ZN => n5397);
   U17348 : OAI22_X1 port map( A1 => n4311, A2 => n21801, B1 => n21806, B2 => 
                           n22458, ZN => n5399);
   U17349 : OAI22_X1 port map( A1 => n4313, A2 => n21801, B1 => n21806, B2 => 
                           n22464, ZN => n5401);
   U17350 : OAI22_X1 port map( A1 => n4315, A2 => n21801, B1 => n21806, B2 => 
                           n22470, ZN => n5403);
   U17351 : OAI22_X1 port map( A1 => n4317, A2 => n21801, B1 => n21806, B2 => 
                           n22476, ZN => n5405);
   U17352 : OAI22_X1 port map( A1 => n4319, A2 => n21801, B1 => n21805, B2 => 
                           n22482, ZN => n5407);
   U17353 : OAI22_X1 port map( A1 => n4321, A2 => n21801, B1 => n21805, B2 => 
                           n22488, ZN => n5409);
   U17354 : OAI22_X1 port map( A1 => n4323, A2 => n21801, B1 => n21805, B2 => 
                           n22494, ZN => n5411);
   U17355 : OAI22_X1 port map( A1 => n4325, A2 => n21801, B1 => n21805, B2 => 
                           n22500, ZN => n5413);
   U17356 : OAI22_X1 port map( A1 => n4327, A2 => n21801, B1 => n21804, B2 => 
                           n22506, ZN => n5415);
   U17357 : OAI22_X1 port map( A1 => n4329, A2 => n21801, B1 => n21804, B2 => 
                           n22512, ZN => n5417);
   U17358 : OAI22_X1 port map( A1 => n4331, A2 => n16832, B1 => n21804, B2 => 
                           n22518, ZN => n5419);
   U17359 : OAI22_X1 port map( A1 => n4333, A2 => n16832, B1 => n21804, B2 => 
                           n22524, ZN => n5421);
   U17360 : OAI22_X1 port map( A1 => n4335, A2 => n16832, B1 => n21803, B2 => 
                           n22530, ZN => n5423);
   U17361 : OAI22_X1 port map( A1 => n4337, A2 => n16832, B1 => n21803, B2 => 
                           n22536, ZN => n5425);
   U17362 : OAI22_X1 port map( A1 => n4339, A2 => n16832, B1 => n21803, B2 => 
                           n22542, ZN => n5427);
   U17363 : OAI22_X1 port map( A1 => n4341, A2 => n16832, B1 => n21803, B2 => 
                           n22548, ZN => n5429);
   U17364 : OAI22_X1 port map( A1 => n4343, A2 => n16832, B1 => n21802, B2 => 
                           n22554, ZN => n5431);
   U17365 : OAI22_X1 port map( A1 => n4345, A2 => n21801, B1 => n21802, B2 => 
                           n22560, ZN => n5433);
   U17366 : OAI22_X1 port map( A1 => n4347, A2 => n21801, B1 => n21802, B2 => 
                           n22566, ZN => n5435);
   U17367 : OAI22_X1 port map( A1 => n4349, A2 => n21801, B1 => n21802, B2 => 
                           n22581, ZN => n5437);
   U17368 : OAI22_X1 port map( A1 => n19615, A2 => n19616, B1 => n4254, B2 => 
                           n18417, ZN => n5342);
   U17369 : NOR4_X1 port map( A1 => n19617, A2 => n19618, A3 => n19619, A4 => 
                           n19620, ZN => n19615);
   U17370 : OAI221_X1 port map( B1 => n16098, B2 => n21190, C1 => n16064, C2 =>
                           n21197, A => n19627, ZN => n19619);
   U17371 : NAND4_X1 port map( A1 => n19628, A2 => n19629, A3 => n19630, A4 => 
                           n19631, ZN => n19618);
   U17372 : OAI22_X1 port map( A1 => n18342, A2 => n18343, B1 => n4286, B2 => 
                           n16834, ZN => n5374);
   U17373 : NOR4_X1 port map( A1 => n18344, A2 => n18345, A3 => n18346, A4 => 
                           n18347, ZN => n18342);
   U17374 : OAI221_X1 port map( B1 => n16098, B2 => n21747, C1 => n16064, C2 =>
                           n21754, A => n18354, ZN => n18346);
   U17375 : NAND4_X1 port map( A1 => n18355, A2 => n18356, A3 => n18357, A4 => 
                           n18358, ZN => n18345);
   U17376 : OAI22_X1 port map( A1 => n21809, A2 => n22381, B1 => n4287, B2 => 
                           n21801, ZN => n5375);
   U17377 : OAI22_X1 port map( A1 => n21817, A2 => n22530, B1 => n4374, B2 => 
                           n16831, ZN => n5462);
   U17378 : OAI22_X1 port map( A1 => n21818, A2 => n22536, B1 => n4375, B2 => 
                           n16831, ZN => n5463);
   U17379 : OAI22_X1 port map( A1 => n21818, A2 => n22542, B1 => n4376, B2 => 
                           n16831, ZN => n5464);
   U17380 : OAI22_X1 port map( A1 => n21818, A2 => n22548, B1 => n4377, B2 => 
                           n21812, ZN => n5465);
   U17381 : OAI22_X1 port map( A1 => n21818, A2 => n22554, B1 => n4378, B2 => 
                           n21812, ZN => n5466);
   U17382 : OAI22_X1 port map( A1 => n21818, A2 => n22560, B1 => n4379, B2 => 
                           n21812, ZN => n5467);
   U17383 : OAI22_X1 port map( A1 => n21819, A2 => n22566, B1 => n4380, B2 => 
                           n21812, ZN => n5468);
   U17384 : OAI22_X1 port map( A1 => n21819, A2 => n22581, B1 => n4381, B2 => 
                           n16831, ZN => n5469);
   U17385 : OAI22_X1 port map( A1 => n21844, A2 => n22529, B1 => n4406, B2 => 
                           n16758, ZN => n5558);
   U17386 : OAI22_X1 port map( A1 => n21845, A2 => n22535, B1 => n4407, B2 => 
                           n16758, ZN => n5559);
   U17387 : OAI22_X1 port map( A1 => n21845, A2 => n22541, B1 => n4408, B2 => 
                           n16758, ZN => n5560);
   U17388 : OAI22_X1 port map( A1 => n21845, A2 => n22547, B1 => n4409, B2 => 
                           n21839, ZN => n5561);
   U17389 : OAI22_X1 port map( A1 => n21845, A2 => n22553, B1 => n4410, B2 => 
                           n21839, ZN => n5562);
   U17390 : OAI22_X1 port map( A1 => n21845, A2 => n22559, B1 => n4411, B2 => 
                           n21839, ZN => n5563);
   U17391 : OAI22_X1 port map( A1 => n21846, A2 => n22565, B1 => n4412, B2 => 
                           n21839, ZN => n5564);
   U17392 : OAI22_X1 port map( A1 => n21846, A2 => n22580, B1 => n4413, B2 => 
                           n16758, ZN => n5565);
   U17393 : OAI22_X1 port map( A1 => n21889, A2 => n22529, B1 => n4502, B2 => 
                           n16618, ZN => n5718);
   U17394 : OAI22_X1 port map( A1 => n21890, A2 => n22535, B1 => n4503, B2 => 
                           n16618, ZN => n5719);
   U17395 : OAI22_X1 port map( A1 => n21890, A2 => n22541, B1 => n4504, B2 => 
                           n16618, ZN => n5720);
   U17396 : OAI22_X1 port map( A1 => n21890, A2 => n22547, B1 => n4505, B2 => 
                           n21884, ZN => n5721);
   U17397 : OAI22_X1 port map( A1 => n21890, A2 => n22553, B1 => n4506, B2 => 
                           n21884, ZN => n5722);
   U17398 : OAI22_X1 port map( A1 => n21890, A2 => n22559, B1 => n4507, B2 => 
                           n21884, ZN => n5723);
   U17399 : OAI22_X1 port map( A1 => n21891, A2 => n22565, B1 => n4508, B2 => 
                           n21884, ZN => n5724);
   U17400 : OAI22_X1 port map( A1 => n21891, A2 => n22580, B1 => n4509, B2 => 
                           n16618, ZN => n5725);
   U17401 : OAI22_X1 port map( A1 => n21898, A2 => n22529, B1 => n8224, B2 => 
                           n16616, ZN => n5750);
   U17402 : OAI22_X1 port map( A1 => n21899, A2 => n22535, B1 => n8256, B2 => 
                           n16616, ZN => n5751);
   U17403 : OAI22_X1 port map( A1 => n21899, A2 => n22541, B1 => n8288, B2 => 
                           n16616, ZN => n5752);
   U17404 : OAI22_X1 port map( A1 => n21899, A2 => n22547, B1 => n8320, B2 => 
                           n21893, ZN => n5753);
   U17405 : OAI22_X1 port map( A1 => n21899, A2 => n22553, B1 => n8352, B2 => 
                           n21893, ZN => n5754);
   U17406 : OAI22_X1 port map( A1 => n21899, A2 => n22559, B1 => n8384, B2 => 
                           n21893, ZN => n5755);
   U17407 : OAI22_X1 port map( A1 => n21900, A2 => n22565, B1 => n8416, B2 => 
                           n21893, ZN => n5756);
   U17408 : OAI22_X1 port map( A1 => n21900, A2 => n22580, B1 => n8448, B2 => 
                           n16616, ZN => n5757);
   U17409 : OAI22_X1 port map( A1 => n21907, A2 => n22529, B1 => n8225, B2 => 
                           n16613, ZN => n5782);
   U17410 : OAI22_X1 port map( A1 => n21908, A2 => n22535, B1 => n8257, B2 => 
                           n16613, ZN => n5783);
   U17411 : OAI22_X1 port map( A1 => n21908, A2 => n22541, B1 => n8289, B2 => 
                           n16613, ZN => n5784);
   U17412 : OAI22_X1 port map( A1 => n21908, A2 => n22547, B1 => n8321, B2 => 
                           n21902, ZN => n5785);
   U17413 : OAI22_X1 port map( A1 => n21908, A2 => n22553, B1 => n8353, B2 => 
                           n21902, ZN => n5786);
   U17414 : OAI22_X1 port map( A1 => n21908, A2 => n22559, B1 => n8385, B2 => 
                           n21902, ZN => n5787);
   U17415 : OAI22_X1 port map( A1 => n21909, A2 => n22565, B1 => n8417, B2 => 
                           n21902, ZN => n5788);
   U17416 : OAI22_X1 port map( A1 => n21909, A2 => n22580, B1 => n8449, B2 => 
                           n16613, ZN => n5789);
   U17417 : OAI22_X1 port map( A1 => n21916, A2 => n22529, B1 => n4534, B2 => 
                           n16610, ZN => n5814);
   U17418 : OAI22_X1 port map( A1 => n21917, A2 => n22535, B1 => n4535, B2 => 
                           n16610, ZN => n5815);
   U17419 : OAI22_X1 port map( A1 => n21917, A2 => n22541, B1 => n4536, B2 => 
                           n16610, ZN => n5816);
   U17420 : OAI22_X1 port map( A1 => n21917, A2 => n22547, B1 => n4537, B2 => 
                           n21911, ZN => n5817);
   U17421 : OAI22_X1 port map( A1 => n21917, A2 => n22553, B1 => n4538, B2 => 
                           n21911, ZN => n5818);
   U17422 : OAI22_X1 port map( A1 => n21917, A2 => n22559, B1 => n4539, B2 => 
                           n21911, ZN => n5819);
   U17423 : OAI22_X1 port map( A1 => n21918, A2 => n22565, B1 => n4540, B2 => 
                           n21911, ZN => n5820);
   U17424 : OAI22_X1 port map( A1 => n21918, A2 => n22580, B1 => n4541, B2 => 
                           n16610, ZN => n5821);
   U17425 : OAI22_X1 port map( A1 => n21997, A2 => n22528, B1 => n4694, B2 => 
                           n16348, ZN => n6102);
   U17426 : OAI22_X1 port map( A1 => n21998, A2 => n22534, B1 => n4695, B2 => 
                           n16348, ZN => n6103);
   U17427 : OAI22_X1 port map( A1 => n21998, A2 => n22540, B1 => n4696, B2 => 
                           n16348, ZN => n6104);
   U17428 : OAI22_X1 port map( A1 => n21998, A2 => n22546, B1 => n4697, B2 => 
                           n21992, ZN => n6105);
   U17429 : OAI22_X1 port map( A1 => n21998, A2 => n22552, B1 => n4698, B2 => 
                           n21992, ZN => n6106);
   U17430 : OAI22_X1 port map( A1 => n21998, A2 => n22558, B1 => n4699, B2 => 
                           n21992, ZN => n6107);
   U17431 : OAI22_X1 port map( A1 => n21999, A2 => n22564, B1 => n4700, B2 => 
                           n21992, ZN => n6108);
   U17432 : OAI22_X1 port map( A1 => n21999, A2 => n22579, B1 => n4701, B2 => 
                           n16348, ZN => n6109);
   U17433 : OAI22_X1 port map( A1 => n22006, A2 => n22528, B1 => n8234, B2 => 
                           n16346, ZN => n6134);
   U17434 : OAI22_X1 port map( A1 => n22007, A2 => n22534, B1 => n8266, B2 => 
                           n16346, ZN => n6135);
   U17435 : OAI22_X1 port map( A1 => n22007, A2 => n22540, B1 => n8298, B2 => 
                           n16346, ZN => n6136);
   U17436 : OAI22_X1 port map( A1 => n22007, A2 => n22546, B1 => n8330, B2 => 
                           n22001, ZN => n6137);
   U17437 : OAI22_X1 port map( A1 => n22007, A2 => n22552, B1 => n8362, B2 => 
                           n22001, ZN => n6138);
   U17438 : OAI22_X1 port map( A1 => n22007, A2 => n22558, B1 => n8394, B2 => 
                           n22001, ZN => n6139);
   U17439 : OAI22_X1 port map( A1 => n22008, A2 => n22564, B1 => n8426, B2 => 
                           n22001, ZN => n6140);
   U17440 : OAI22_X1 port map( A1 => n22008, A2 => n22579, B1 => n8458, B2 => 
                           n16346, ZN => n6141);
   U17441 : OAI22_X1 port map( A1 => n22015, A2 => n22528, B1 => n8235, B2 => 
                           n16343, ZN => n6166);
   U17442 : OAI22_X1 port map( A1 => n22016, A2 => n22534, B1 => n8267, B2 => 
                           n16343, ZN => n6167);
   U17443 : OAI22_X1 port map( A1 => n22016, A2 => n22540, B1 => n8299, B2 => 
                           n16343, ZN => n6168);
   U17444 : OAI22_X1 port map( A1 => n22016, A2 => n22546, B1 => n8331, B2 => 
                           n22010, ZN => n6169);
   U17445 : OAI22_X1 port map( A1 => n22016, A2 => n22552, B1 => n8363, B2 => 
                           n22010, ZN => n6170);
   U17446 : OAI22_X1 port map( A1 => n22016, A2 => n22558, B1 => n8395, B2 => 
                           n22010, ZN => n6171);
   U17447 : OAI22_X1 port map( A1 => n22017, A2 => n22564, B1 => n8427, B2 => 
                           n22010, ZN => n6172);
   U17448 : OAI22_X1 port map( A1 => n22017, A2 => n22579, B1 => n8459, B2 => 
                           n16343, ZN => n6173);
   U17449 : OAI22_X1 port map( A1 => n22069, A2 => n22527, B1 => n4822, B2 => 
                           n16169, ZN => n6358);
   U17450 : OAI22_X1 port map( A1 => n22070, A2 => n22533, B1 => n4823, B2 => 
                           n16169, ZN => n6359);
   U17451 : OAI22_X1 port map( A1 => n22070, A2 => n22539, B1 => n4824, B2 => 
                           n16169, ZN => n6360);
   U17452 : OAI22_X1 port map( A1 => n22070, A2 => n22545, B1 => n4825, B2 => 
                           n22064, ZN => n6361);
   U17453 : OAI22_X1 port map( A1 => n22070, A2 => n22551, B1 => n4826, B2 => 
                           n22064, ZN => n6362);
   U17454 : OAI22_X1 port map( A1 => n22070, A2 => n22557, B1 => n4827, B2 => 
                           n22064, ZN => n6363);
   U17455 : OAI22_X1 port map( A1 => n22071, A2 => n22563, B1 => n4828, B2 => 
                           n22064, ZN => n6364);
   U17456 : OAI22_X1 port map( A1 => n22071, A2 => n22578, B1 => n4829, B2 => 
                           n16169, ZN => n6365);
   U17457 : OAI22_X1 port map( A1 => n22150, A2 => n22527, B1 => n8242, B2 => 
                           n15893, ZN => n6646);
   U17458 : OAI22_X1 port map( A1 => n22151, A2 => n22533, B1 => n8274, B2 => 
                           n15893, ZN => n6647);
   U17459 : OAI22_X1 port map( A1 => n22151, A2 => n22539, B1 => n8306, B2 => 
                           n15893, ZN => n6648);
   U17460 : OAI22_X1 port map( A1 => n22151, A2 => n22545, B1 => n8338, B2 => 
                           n22145, ZN => n6649);
   U17461 : OAI22_X1 port map( A1 => n22151, A2 => n22551, B1 => n8370, B2 => 
                           n22145, ZN => n6650);
   U17462 : OAI22_X1 port map( A1 => n22151, A2 => n22557, B1 => n8402, B2 => 
                           n22145, ZN => n6651);
   U17463 : OAI22_X1 port map( A1 => n22152, A2 => n22563, B1 => n8434, B2 => 
                           n22145, ZN => n6652);
   U17464 : OAI22_X1 port map( A1 => n22152, A2 => n22578, B1 => n8466, B2 => 
                           n15893, ZN => n6653);
   U17465 : OAI22_X1 port map( A1 => n22159, A2 => n22527, B1 => n8243, B2 => 
                           n15890, ZN => n6678);
   U17466 : OAI22_X1 port map( A1 => n22160, A2 => n22533, B1 => n8275, B2 => 
                           n15890, ZN => n6679);
   U17467 : OAI22_X1 port map( A1 => n22160, A2 => n22539, B1 => n8307, B2 => 
                           n15890, ZN => n6680);
   U17468 : OAI22_X1 port map( A1 => n22160, A2 => n22545, B1 => n8339, B2 => 
                           n22154, ZN => n6681);
   U17469 : OAI22_X1 port map( A1 => n22160, A2 => n22551, B1 => n8371, B2 => 
                           n22154, ZN => n6682);
   U17470 : OAI22_X1 port map( A1 => n22160, A2 => n22557, B1 => n8403, B2 => 
                           n22154, ZN => n6683);
   U17471 : OAI22_X1 port map( A1 => n22161, A2 => n22563, B1 => n8435, B2 => 
                           n22154, ZN => n6684);
   U17472 : OAI22_X1 port map( A1 => n22161, A2 => n22578, B1 => n8467, B2 => 
                           n15890, ZN => n6685);
   U17473 : OAI22_X1 port map( A1 => n22204, A2 => n22526, B1 => n5046, B2 => 
                           n15750, ZN => n6838);
   U17474 : OAI22_X1 port map( A1 => n22205, A2 => n22532, B1 => n5047, B2 => 
                           n15750, ZN => n6839);
   U17475 : OAI22_X1 port map( A1 => n22205, A2 => n22538, B1 => n5048, B2 => 
                           n15750, ZN => n6840);
   U17476 : OAI22_X1 port map( A1 => n22205, A2 => n22544, B1 => n5049, B2 => 
                           n22199, ZN => n6841);
   U17477 : OAI22_X1 port map( A1 => n22205, A2 => n22550, B1 => n5050, B2 => 
                           n22199, ZN => n6842);
   U17478 : OAI22_X1 port map( A1 => n22205, A2 => n22556, B1 => n5051, B2 => 
                           n22199, ZN => n6843);
   U17479 : OAI22_X1 port map( A1 => n22206, A2 => n22562, B1 => n5052, B2 => 
                           n22199, ZN => n6844);
   U17480 : OAI22_X1 port map( A1 => n22206, A2 => n22577, B1 => n5053, B2 => 
                           n15750, ZN => n6845);
   U17481 : OAI22_X1 port map( A1 => n22366, A2 => n22525, B1 => n8246, B2 => 
                           n15155, ZN => n7414);
   U17482 : OAI22_X1 port map( A1 => n22367, A2 => n22531, B1 => n8278, B2 => 
                           n15155, ZN => n7415);
   U17483 : OAI22_X1 port map( A1 => n22367, A2 => n22537, B1 => n8310, B2 => 
                           n15155, ZN => n7416);
   U17484 : OAI22_X1 port map( A1 => n22367, A2 => n22543, B1 => n8342, B2 => 
                           n22361, ZN => n7417);
   U17485 : OAI22_X1 port map( A1 => n22367, A2 => n22549, B1 => n8374, B2 => 
                           n22361, ZN => n7418);
   U17486 : OAI22_X1 port map( A1 => n22367, A2 => n22555, B1 => n8406, B2 => 
                           n22361, ZN => n7419);
   U17487 : OAI22_X1 port map( A1 => n22368, A2 => n22561, B1 => n8438, B2 => 
                           n22361, ZN => n7420);
   U17488 : OAI22_X1 port map( A1 => n22368, A2 => n22576, B1 => n8470, B2 => 
                           n15155, ZN => n7421);
   U17489 : OAI22_X1 port map( A1 => n22572, A2 => n22525, B1 => n8247, B2 => 
                           n15119, ZN => n7446);
   U17490 : OAI22_X1 port map( A1 => n22573, A2 => n22531, B1 => n8279, B2 => 
                           n15119, ZN => n7447);
   U17491 : OAI22_X1 port map( A1 => n22573, A2 => n22537, B1 => n8311, B2 => 
                           n15119, ZN => n7448);
   U17492 : OAI22_X1 port map( A1 => n22573, A2 => n22543, B1 => n8343, B2 => 
                           n22567, ZN => n7449);
   U17493 : OAI22_X1 port map( A1 => n22573, A2 => n22549, B1 => n8375, B2 => 
                           n22567, ZN => n7450);
   U17494 : OAI22_X1 port map( A1 => n22573, A2 => n22555, B1 => n8407, B2 => 
                           n22567, ZN => n7451);
   U17495 : OAI22_X1 port map( A1 => n22574, A2 => n22561, B1 => n8439, B2 => 
                           n22567, ZN => n7452);
   U17496 : OAI22_X1 port map( A1 => n22574, A2 => n22576, B1 => n8471, B2 => 
                           n15119, ZN => n7453);
   U17497 : AOI22_X1 port map( A1 => n21070, A2 => n9803, B1 => n21101, B2 => 
                           n19998, ZN => n18971);
   U17498 : AOI22_X1 port map( A1 => n20783, A2 => n9169, B1 => n20837, B2 => 
                           n8721, ZN => n18973);
   U17499 : AOI22_X1 port map( A1 => n20976, A2 => n19935, B1 => n20934, B2 => 
                           n9899, ZN => n18974);
   U17500 : AOI22_X1 port map( A1 => n21070, A2 => n9802, B1 => n21102, B2 => 
                           n19690, ZN => n18934);
   U17501 : AOI22_X1 port map( A1 => n20783, A2 => n9158, B1 => n20838, B2 => 
                           n8710, ZN => n18936);
   U17502 : AOI22_X1 port map( A1 => n20976, A2 => n19687, B1 => n20935, B2 => 
                           n9898, ZN => n18937);
   U17503 : AOI22_X1 port map( A1 => n21025, A2 => n19688, B1 => n20719, B2 => 
                           n8701, ZN => n18898);
   U17504 : AOI22_X1 port map( A1 => n20781, A2 => n9147, B1 => n20838, B2 => 
                           n8699, ZN => n18899);
   U17505 : AOI22_X1 port map( A1 => n20977, A2 => n19689, B1 => n20935, B2 => 
                           n9897, ZN => n18900);
   U17506 : AOI22_X1 port map( A1 => n21065, A2 => n9800, B1 => n21103, B2 => 
                           n19691, ZN => n18860);
   U17507 : AOI22_X1 port map( A1 => n20778, A2 => n9136, B1 => n20837, B2 => 
                           n8688, ZN => n18862);
   U17508 : AOI22_X1 port map( A1 => n20970, A2 => n19936, B1 => n20934, B2 => 
                           n9896, ZN => n18863);
   U17509 : AOI22_X1 port map( A1 => n21627, A2 => n9803, B1 => n21658, B2 => 
                           n19998, ZN => n17520);
   U17510 : AOI22_X1 port map( A1 => n21340, A2 => n9169, B1 => n21394, B2 => 
                           n8721, ZN => n17524);
   U17511 : AOI22_X1 port map( A1 => n21533, A2 => n19935, B1 => n21491, B2 => 
                           n9899, ZN => n17525);
   U17512 : AOI22_X1 port map( A1 => n21627, A2 => n9802, B1 => n21659, B2 => 
                           n19690, ZN => n17473);
   U17513 : AOI22_X1 port map( A1 => n21340, A2 => n9158, B1 => n21395, B2 => 
                           n8710, ZN => n17477);
   U17514 : AOI22_X1 port map( A1 => n21533, A2 => n19687, B1 => n21492, B2 => 
                           n9898, ZN => n17478);
   U17515 : AOI22_X1 port map( A1 => n21582, A2 => n19688, B1 => n21276, B2 => 
                           n8701, ZN => n17428);
   U17516 : AOI22_X1 port map( A1 => n21338, A2 => n9147, B1 => n21395, B2 => 
                           n8699, ZN => n17430);
   U17517 : AOI22_X1 port map( A1 => n21534, A2 => n19689, B1 => n21492, B2 => 
                           n9897, ZN => n17431);
   U17518 : AOI22_X1 port map( A1 => n21622, A2 => n9800, B1 => n21660, B2 => 
                           n19691, ZN => n17379);
   U17519 : AOI22_X1 port map( A1 => n21335, A2 => n9136, B1 => n21394, B2 => 
                           n8688, ZN => n17383);
   U17520 : AOI22_X1 port map( A1 => n21527, A2 => n19936, B1 => n21491, B2 => 
                           n9896, ZN => n17384);
   U17521 : AOI22_X1 port map( A1 => n21206, A2 => n8572, B1 => n21210, B2 => 
                           n9020, ZN => n19627);
   U17522 : AOI22_X1 port map( A1 => n21763, A2 => n8572, B1 => n21767, B2 => 
                           n9020, ZN => n18354);
   U17523 : OAI22_X1 port map( A1 => n21822, A2 => n22381, B1 => n21821, B2 => 
                           n20046, ZN => n5470);
   U17524 : OAI22_X1 port map( A1 => n21822, A2 => n22392, B1 => n21821, B2 => 
                           n16828, ZN => n5471);
   U17525 : OAI22_X1 port map( A1 => n21822, A2 => n22398, B1 => n21821, B2 => 
                           n16827, ZN => n5472);
   U17526 : OAI22_X1 port map( A1 => n21822, A2 => n22404, B1 => n21821, B2 => 
                           n16826, ZN => n5473);
   U17527 : OAI22_X1 port map( A1 => n21822, A2 => n22410, B1 => n21821, B2 => 
                           n16825, ZN => n5474);
   U17528 : OAI22_X1 port map( A1 => n21823, A2 => n22416, B1 => n21821, B2 => 
                           n16824, ZN => n5475);
   U17529 : OAI22_X1 port map( A1 => n21823, A2 => n22422, B1 => n21821, B2 => 
                           n16823, ZN => n5476);
   U17530 : OAI22_X1 port map( A1 => n21823, A2 => n22428, B1 => n21821, B2 => 
                           n16822, ZN => n5477);
   U17531 : OAI22_X1 port map( A1 => n21823, A2 => n22434, B1 => n21821, B2 => 
                           n16821, ZN => n5478);
   U17532 : OAI22_X1 port map( A1 => n21823, A2 => n22440, B1 => n21821, B2 => 
                           n16820, ZN => n5479);
   U17533 : OAI22_X1 port map( A1 => n21824, A2 => n22446, B1 => n21821, B2 => 
                           n16819, ZN => n5480);
   U17534 : OAI22_X1 port map( A1 => n21824, A2 => n22452, B1 => n21821, B2 => 
                           n16818, ZN => n5481);
   U17535 : OAI22_X1 port map( A1 => n21824, A2 => n22458, B1 => n21821, B2 => 
                           n16817, ZN => n5482);
   U17536 : OAI22_X1 port map( A1 => n21824, A2 => n22464, B1 => n21821, B2 => 
                           n16816, ZN => n5483);
   U17537 : OAI22_X1 port map( A1 => n21824, A2 => n22470, B1 => n16797, B2 => 
                           n16815, ZN => n5484);
   U17538 : OAI22_X1 port map( A1 => n21825, A2 => n22476, B1 => n16797, B2 => 
                           n16814, ZN => n5485);
   U17539 : OAI22_X1 port map( A1 => n21825, A2 => n22482, B1 => n16797, B2 => 
                           n16813, ZN => n5486);
   U17540 : OAI22_X1 port map( A1 => n21825, A2 => n22488, B1 => n16797, B2 => 
                           n16812, ZN => n5487);
   U17541 : OAI22_X1 port map( A1 => n21825, A2 => n22494, B1 => n16797, B2 => 
                           n16811, ZN => n5488);
   U17542 : OAI22_X1 port map( A1 => n21825, A2 => n22500, B1 => n16797, B2 => 
                           n16810, ZN => n5489);
   U17543 : OAI22_X1 port map( A1 => n21826, A2 => n22506, B1 => n16797, B2 => 
                           n16809, ZN => n5490);
   U17544 : OAI22_X1 port map( A1 => n21826, A2 => n22512, B1 => n21821, B2 => 
                           n16808, ZN => n5491);
   U17545 : OAI22_X1 port map( A1 => n21826, A2 => n22518, B1 => n21821, B2 => 
                           n16807, ZN => n5492);
   U17546 : OAI22_X1 port map( A1 => n21826, A2 => n22524, B1 => n21821, B2 => 
                           n16806, ZN => n5493);
   U17547 : OAI22_X1 port map( A1 => n21831, A2 => n22381, B1 => n21830, B2 => 
                           n20047, ZN => n5502);
   U17548 : OAI22_X1 port map( A1 => n21831, A2 => n22392, B1 => n21830, B2 => 
                           n16791, ZN => n5503);
   U17549 : OAI22_X1 port map( A1 => n21831, A2 => n22398, B1 => n21830, B2 => 
                           n16790, ZN => n5504);
   U17550 : OAI22_X1 port map( A1 => n21831, A2 => n22404, B1 => n21830, B2 => 
                           n16789, ZN => n5505);
   U17551 : OAI22_X1 port map( A1 => n21831, A2 => n22410, B1 => n21830, B2 => 
                           n16788, ZN => n5506);
   U17552 : OAI22_X1 port map( A1 => n21832, A2 => n22416, B1 => n21830, B2 => 
                           n16787, ZN => n5507);
   U17553 : OAI22_X1 port map( A1 => n21832, A2 => n22422, B1 => n21830, B2 => 
                           n16786, ZN => n5508);
   U17554 : OAI22_X1 port map( A1 => n21832, A2 => n22428, B1 => n21830, B2 => 
                           n16785, ZN => n5509);
   U17555 : OAI22_X1 port map( A1 => n21832, A2 => n22434, B1 => n21830, B2 => 
                           n16784, ZN => n5510);
   U17556 : OAI22_X1 port map( A1 => n21832, A2 => n22440, B1 => n21830, B2 => 
                           n16783, ZN => n5511);
   U17557 : OAI22_X1 port map( A1 => n21833, A2 => n22446, B1 => n21830, B2 => 
                           n16782, ZN => n5512);
   U17558 : OAI22_X1 port map( A1 => n21833, A2 => n22452, B1 => n21830, B2 => 
                           n16781, ZN => n5513);
   U17559 : OAI22_X1 port map( A1 => n21833, A2 => n22458, B1 => n21830, B2 => 
                           n16780, ZN => n5514);
   U17560 : OAI22_X1 port map( A1 => n21833, A2 => n22464, B1 => n21830, B2 => 
                           n16779, ZN => n5515);
   U17561 : OAI22_X1 port map( A1 => n21833, A2 => n22470, B1 => n16760, B2 => 
                           n16778, ZN => n5516);
   U17562 : OAI22_X1 port map( A1 => n21834, A2 => n22476, B1 => n16760, B2 => 
                           n16777, ZN => n5517);
   U17563 : OAI22_X1 port map( A1 => n21834, A2 => n22482, B1 => n16760, B2 => 
                           n16776, ZN => n5518);
   U17564 : OAI22_X1 port map( A1 => n21834, A2 => n22488, B1 => n16760, B2 => 
                           n16775, ZN => n5519);
   U17565 : OAI22_X1 port map( A1 => n21834, A2 => n22494, B1 => n16760, B2 => 
                           n16774, ZN => n5520);
   U17566 : OAI22_X1 port map( A1 => n21834, A2 => n22500, B1 => n16760, B2 => 
                           n16773, ZN => n5521);
   U17567 : OAI22_X1 port map( A1 => n21835, A2 => n22506, B1 => n16760, B2 => 
                           n16772, ZN => n5522);
   U17568 : OAI22_X1 port map( A1 => n21835, A2 => n22512, B1 => n21830, B2 => 
                           n16771, ZN => n5523);
   U17569 : OAI22_X1 port map( A1 => n21835, A2 => n22518, B1 => n21830, B2 => 
                           n16770, ZN => n5524);
   U17570 : OAI22_X1 port map( A1 => n21835, A2 => n22524, B1 => n21830, B2 => 
                           n16769, ZN => n5525);
   U17571 : OAI22_X1 port map( A1 => n21858, A2 => n22381, B1 => n21857, B2 => 
                           n20212, ZN => n5598);
   U17572 : OAI22_X1 port map( A1 => n21858, A2 => n22391, B1 => n21857, B2 => 
                           n20213, ZN => n5599);
   U17573 : OAI22_X1 port map( A1 => n21858, A2 => n22397, B1 => n21857, B2 => 
                           n20214, ZN => n5600);
   U17574 : OAI22_X1 port map( A1 => n21858, A2 => n22403, B1 => n21857, B2 => 
                           n20215, ZN => n5601);
   U17575 : OAI22_X1 port map( A1 => n21858, A2 => n22409, B1 => n21857, B2 => 
                           n20216, ZN => n5602);
   U17576 : OAI22_X1 port map( A1 => n21859, A2 => n22415, B1 => n21857, B2 => 
                           n20217, ZN => n5603);
   U17577 : OAI22_X1 port map( A1 => n21859, A2 => n22421, B1 => n21857, B2 => 
                           n20218, ZN => n5604);
   U17578 : OAI22_X1 port map( A1 => n21859, A2 => n22427, B1 => n21857, B2 => 
                           n20219, ZN => n5605);
   U17579 : OAI22_X1 port map( A1 => n21859, A2 => n22433, B1 => n21857, B2 => 
                           n20220, ZN => n5606);
   U17580 : OAI22_X1 port map( A1 => n21859, A2 => n22439, B1 => n21857, B2 => 
                           n20221, ZN => n5607);
   U17581 : OAI22_X1 port map( A1 => n21860, A2 => n22445, B1 => n21857, B2 => 
                           n20222, ZN => n5608);
   U17582 : OAI22_X1 port map( A1 => n21860, A2 => n22451, B1 => n21857, B2 => 
                           n20223, ZN => n5609);
   U17583 : OAI22_X1 port map( A1 => n21860, A2 => n22457, B1 => n21857, B2 => 
                           n20224, ZN => n5610);
   U17584 : OAI22_X1 port map( A1 => n21860, A2 => n22463, B1 => n21857, B2 => 
                           n20225, ZN => n5611);
   U17585 : OAI22_X1 port map( A1 => n21860, A2 => n22469, B1 => n16690, B2 => 
                           n20226, ZN => n5612);
   U17586 : OAI22_X1 port map( A1 => n21861, A2 => n22475, B1 => n16690, B2 => 
                           n20227, ZN => n5613);
   U17587 : OAI22_X1 port map( A1 => n21861, A2 => n22481, B1 => n16690, B2 => 
                           n20228, ZN => n5614);
   U17588 : OAI22_X1 port map( A1 => n21861, A2 => n22487, B1 => n16690, B2 => 
                           n20229, ZN => n5615);
   U17589 : OAI22_X1 port map( A1 => n21861, A2 => n22493, B1 => n16690, B2 => 
                           n20230, ZN => n5616);
   U17590 : OAI22_X1 port map( A1 => n21861, A2 => n22499, B1 => n16690, B2 => 
                           n20231, ZN => n5617);
   U17591 : OAI22_X1 port map( A1 => n21862, A2 => n22505, B1 => n16690, B2 => 
                           n20232, ZN => n5618);
   U17592 : OAI22_X1 port map( A1 => n21862, A2 => n22511, B1 => n21857, B2 => 
                           n20233, ZN => n5619);
   U17593 : OAI22_X1 port map( A1 => n21862, A2 => n22517, B1 => n21857, B2 => 
                           n20234, ZN => n5620);
   U17594 : OAI22_X1 port map( A1 => n21862, A2 => n22523, B1 => n21857, B2 => 
                           n20235, ZN => n5621);
   U17595 : OAI22_X1 port map( A1 => n21867, A2 => n22381, B1 => n21866, B2 => 
                           n20236, ZN => n5630);
   U17596 : OAI22_X1 port map( A1 => n21867, A2 => n22391, B1 => n21866, B2 => 
                           n20237, ZN => n5631);
   U17597 : OAI22_X1 port map( A1 => n21867, A2 => n22397, B1 => n21866, B2 => 
                           n20238, ZN => n5632);
   U17598 : OAI22_X1 port map( A1 => n21867, A2 => n22403, B1 => n21866, B2 => 
                           n20239, ZN => n5633);
   U17599 : OAI22_X1 port map( A1 => n21867, A2 => n22409, B1 => n21866, B2 => 
                           n20240, ZN => n5634);
   U17600 : OAI22_X1 port map( A1 => n21868, A2 => n22415, B1 => n21866, B2 => 
                           n20241, ZN => n5635);
   U17601 : OAI22_X1 port map( A1 => n21868, A2 => n22421, B1 => n21866, B2 => 
                           n20242, ZN => n5636);
   U17602 : OAI22_X1 port map( A1 => n21868, A2 => n22427, B1 => n21866, B2 => 
                           n20243, ZN => n5637);
   U17603 : OAI22_X1 port map( A1 => n21868, A2 => n22433, B1 => n21866, B2 => 
                           n20244, ZN => n5638);
   U17604 : OAI22_X1 port map( A1 => n21868, A2 => n22439, B1 => n21866, B2 => 
                           n20245, ZN => n5639);
   U17605 : OAI22_X1 port map( A1 => n21869, A2 => n22445, B1 => n21866, B2 => 
                           n20246, ZN => n5640);
   U17606 : OAI22_X1 port map( A1 => n21869, A2 => n22451, B1 => n21866, B2 => 
                           n20247, ZN => n5641);
   U17607 : OAI22_X1 port map( A1 => n21869, A2 => n22457, B1 => n21866, B2 => 
                           n20248, ZN => n5642);
   U17608 : OAI22_X1 port map( A1 => n21869, A2 => n22463, B1 => n21866, B2 => 
                           n20249, ZN => n5643);
   U17609 : OAI22_X1 port map( A1 => n21869, A2 => n22469, B1 => n16655, B2 => 
                           n20250, ZN => n5644);
   U17610 : OAI22_X1 port map( A1 => n21870, A2 => n22475, B1 => n16655, B2 => 
                           n20251, ZN => n5645);
   U17611 : OAI22_X1 port map( A1 => n21870, A2 => n22481, B1 => n16655, B2 => 
                           n20252, ZN => n5646);
   U17612 : OAI22_X1 port map( A1 => n21870, A2 => n22487, B1 => n16655, B2 => 
                           n20253, ZN => n5647);
   U17613 : OAI22_X1 port map( A1 => n21870, A2 => n22493, B1 => n16655, B2 => 
                           n20254, ZN => n5648);
   U17614 : OAI22_X1 port map( A1 => n21870, A2 => n22499, B1 => n16655, B2 => 
                           n20255, ZN => n5649);
   U17615 : OAI22_X1 port map( A1 => n21871, A2 => n22505, B1 => n16655, B2 => 
                           n20256, ZN => n5650);
   U17616 : OAI22_X1 port map( A1 => n21871, A2 => n22511, B1 => n21866, B2 => 
                           n20257, ZN => n5651);
   U17617 : OAI22_X1 port map( A1 => n21871, A2 => n22517, B1 => n21866, B2 => 
                           n20258, ZN => n5652);
   U17618 : OAI22_X1 port map( A1 => n21871, A2 => n22523, B1 => n21866, B2 => 
                           n20259, ZN => n5653);
   U17619 : OAI22_X1 port map( A1 => n21876, A2 => n22381, B1 => n21875, B2 => 
                           n16652, ZN => n5662);
   U17620 : OAI22_X1 port map( A1 => n21876, A2 => n22391, B1 => n21875, B2 => 
                           n20097, ZN => n5663);
   U17621 : OAI22_X1 port map( A1 => n21876, A2 => n22397, B1 => n21875, B2 => 
                           n20098, ZN => n5664);
   U17622 : OAI22_X1 port map( A1 => n21876, A2 => n22403, B1 => n21875, B2 => 
                           n20099, ZN => n5665);
   U17623 : OAI22_X1 port map( A1 => n21876, A2 => n22409, B1 => n21875, B2 => 
                           n20100, ZN => n5666);
   U17624 : OAI22_X1 port map( A1 => n21877, A2 => n22415, B1 => n21875, B2 => 
                           n20101, ZN => n5667);
   U17625 : OAI22_X1 port map( A1 => n21877, A2 => n22421, B1 => n21875, B2 => 
                           n20102, ZN => n5668);
   U17626 : OAI22_X1 port map( A1 => n21877, A2 => n22427, B1 => n21875, B2 => 
                           n20103, ZN => n5669);
   U17627 : OAI22_X1 port map( A1 => n21877, A2 => n22433, B1 => n21875, B2 => 
                           n20104, ZN => n5670);
   U17628 : OAI22_X1 port map( A1 => n21877, A2 => n22439, B1 => n21875, B2 => 
                           n20105, ZN => n5671);
   U17629 : OAI22_X1 port map( A1 => n21878, A2 => n22445, B1 => n21875, B2 => 
                           n20106, ZN => n5672);
   U17630 : OAI22_X1 port map( A1 => n21878, A2 => n22451, B1 => n21875, B2 => 
                           n20107, ZN => n5673);
   U17631 : OAI22_X1 port map( A1 => n21878, A2 => n22457, B1 => n21875, B2 => 
                           n20108, ZN => n5674);
   U17632 : OAI22_X1 port map( A1 => n21878, A2 => n22463, B1 => n21875, B2 => 
                           n20109, ZN => n5675);
   U17633 : OAI22_X1 port map( A1 => n21878, A2 => n22469, B1 => n16620, B2 => 
                           n20110, ZN => n5676);
   U17634 : OAI22_X1 port map( A1 => n21879, A2 => n22475, B1 => n16620, B2 => 
                           n20111, ZN => n5677);
   U17635 : OAI22_X1 port map( A1 => n21879, A2 => n22481, B1 => n16620, B2 => 
                           n20112, ZN => n5678);
   U17636 : OAI22_X1 port map( A1 => n21879, A2 => n22487, B1 => n16620, B2 => 
                           n20113, ZN => n5679);
   U17637 : OAI22_X1 port map( A1 => n21879, A2 => n22493, B1 => n16620, B2 => 
                           n20114, ZN => n5680);
   U17638 : OAI22_X1 port map( A1 => n21879, A2 => n22499, B1 => n16620, B2 => 
                           n20115, ZN => n5681);
   U17639 : OAI22_X1 port map( A1 => n21880, A2 => n22505, B1 => n16620, B2 => 
                           n20116, ZN => n5682);
   U17640 : OAI22_X1 port map( A1 => n21880, A2 => n22511, B1 => n21875, B2 => 
                           n20117, ZN => n5683);
   U17641 : OAI22_X1 port map( A1 => n21880, A2 => n22517, B1 => n21875, B2 => 
                           n20118, ZN => n5684);
   U17642 : OAI22_X1 port map( A1 => n21880, A2 => n22523, B1 => n21875, B2 => 
                           n20119, ZN => n5685);
   U17643 : OAI22_X1 port map( A1 => n21921, A2 => n22382, B1 => n21920, B2 => 
                           n16608, ZN => n5822);
   U17644 : OAI22_X1 port map( A1 => n21921, A2 => n22391, B1 => n21920, B2 => 
                           n20000, ZN => n5823);
   U17645 : OAI22_X1 port map( A1 => n21921, A2 => n22397, B1 => n21920, B2 => 
                           n20001, ZN => n5824);
   U17646 : OAI22_X1 port map( A1 => n21921, A2 => n22403, B1 => n21920, B2 => 
                           n20002, ZN => n5825);
   U17647 : OAI22_X1 port map( A1 => n21921, A2 => n22409, B1 => n21920, B2 => 
                           n20003, ZN => n5826);
   U17648 : OAI22_X1 port map( A1 => n21922, A2 => n22415, B1 => n21920, B2 => 
                           n20004, ZN => n5827);
   U17649 : OAI22_X1 port map( A1 => n21922, A2 => n22421, B1 => n21920, B2 => 
                           n20005, ZN => n5828);
   U17650 : OAI22_X1 port map( A1 => n21922, A2 => n22427, B1 => n21920, B2 => 
                           n20006, ZN => n5829);
   U17651 : OAI22_X1 port map( A1 => n21922, A2 => n22433, B1 => n21920, B2 => 
                           n20007, ZN => n5830);
   U17652 : OAI22_X1 port map( A1 => n21922, A2 => n22439, B1 => n21920, B2 => 
                           n20008, ZN => n5831);
   U17653 : OAI22_X1 port map( A1 => n21923, A2 => n22445, B1 => n21920, B2 => 
                           n20009, ZN => n5832);
   U17654 : OAI22_X1 port map( A1 => n21923, A2 => n22451, B1 => n21920, B2 => 
                           n20010, ZN => n5833);
   U17655 : OAI22_X1 port map( A1 => n21923, A2 => n22457, B1 => n21920, B2 => 
                           n20011, ZN => n5834);
   U17656 : OAI22_X1 port map( A1 => n21923, A2 => n22463, B1 => n21920, B2 => 
                           n20012, ZN => n5835);
   U17657 : OAI22_X1 port map( A1 => n21923, A2 => n22469, B1 => n16576, B2 => 
                           n20013, ZN => n5836);
   U17658 : OAI22_X1 port map( A1 => n21924, A2 => n22475, B1 => n16576, B2 => 
                           n20014, ZN => n5837);
   U17659 : OAI22_X1 port map( A1 => n21924, A2 => n22481, B1 => n16576, B2 => 
                           n20015, ZN => n5838);
   U17660 : OAI22_X1 port map( A1 => n21924, A2 => n22487, B1 => n16576, B2 => 
                           n20016, ZN => n5839);
   U17661 : OAI22_X1 port map( A1 => n21924, A2 => n22493, B1 => n16576, B2 => 
                           n20017, ZN => n5840);
   U17662 : OAI22_X1 port map( A1 => n21924, A2 => n22499, B1 => n16576, B2 => 
                           n20018, ZN => n5841);
   U17663 : OAI22_X1 port map( A1 => n21925, A2 => n22505, B1 => n16576, B2 => 
                           n20019, ZN => n5842);
   U17664 : OAI22_X1 port map( A1 => n21925, A2 => n22511, B1 => n21920, B2 => 
                           n20020, ZN => n5843);
   U17665 : OAI22_X1 port map( A1 => n21925, A2 => n22517, B1 => n21920, B2 => 
                           n20021, ZN => n5844);
   U17666 : OAI22_X1 port map( A1 => n21925, A2 => n22523, B1 => n21920, B2 => 
                           n20022, ZN => n5845);
   U17667 : OAI22_X1 port map( A1 => n21957, A2 => n22382, B1 => n21956, B2 => 
                           n16485, ZN => n5950);
   U17668 : OAI22_X1 port map( A1 => n21957, A2 => n22390, B1 => n21956, B2 => 
                           n16484, ZN => n5951);
   U17669 : OAI22_X1 port map( A1 => n21957, A2 => n22396, B1 => n21956, B2 => 
                           n16483, ZN => n5952);
   U17670 : OAI22_X1 port map( A1 => n21957, A2 => n22402, B1 => n21956, B2 => 
                           n16482, ZN => n5953);
   U17671 : OAI22_X1 port map( A1 => n21957, A2 => n22408, B1 => n21956, B2 => 
                           n16481, ZN => n5954);
   U17672 : OAI22_X1 port map( A1 => n21958, A2 => n22414, B1 => n21956, B2 => 
                           n16480, ZN => n5955);
   U17673 : OAI22_X1 port map( A1 => n21958, A2 => n22420, B1 => n21956, B2 => 
                           n16479, ZN => n5956);
   U17674 : OAI22_X1 port map( A1 => n21958, A2 => n22426, B1 => n21956, B2 => 
                           n16478, ZN => n5957);
   U17675 : OAI22_X1 port map( A1 => n21958, A2 => n22432, B1 => n21956, B2 => 
                           n16477, ZN => n5958);
   U17676 : OAI22_X1 port map( A1 => n21958, A2 => n22438, B1 => n21956, B2 => 
                           n16476, ZN => n5959);
   U17677 : OAI22_X1 port map( A1 => n21959, A2 => n22444, B1 => n21956, B2 => 
                           n16475, ZN => n5960);
   U17678 : OAI22_X1 port map( A1 => n21959, A2 => n22450, B1 => n21956, B2 => 
                           n16474, ZN => n5961);
   U17679 : OAI22_X1 port map( A1 => n21959, A2 => n22456, B1 => n21956, B2 => 
                           n16473, ZN => n5962);
   U17680 : OAI22_X1 port map( A1 => n21959, A2 => n22462, B1 => n21956, B2 => 
                           n16472, ZN => n5963);
   U17681 : OAI22_X1 port map( A1 => n21959, A2 => n22468, B1 => n16453, B2 => 
                           n16471, ZN => n5964);
   U17682 : OAI22_X1 port map( A1 => n21960, A2 => n22474, B1 => n16453, B2 => 
                           n16470, ZN => n5965);
   U17683 : OAI22_X1 port map( A1 => n21960, A2 => n22480, B1 => n16453, B2 => 
                           n16469, ZN => n5966);
   U17684 : OAI22_X1 port map( A1 => n21960, A2 => n22486, B1 => n16453, B2 => 
                           n16468, ZN => n5967);
   U17685 : OAI22_X1 port map( A1 => n21960, A2 => n22492, B1 => n16453, B2 => 
                           n16467, ZN => n5968);
   U17686 : OAI22_X1 port map( A1 => n21960, A2 => n22498, B1 => n16453, B2 => 
                           n16466, ZN => n5969);
   U17687 : OAI22_X1 port map( A1 => n21961, A2 => n22504, B1 => n16453, B2 => 
                           n16465, ZN => n5970);
   U17688 : OAI22_X1 port map( A1 => n21961, A2 => n22510, B1 => n21956, B2 => 
                           n16464, ZN => n5971);
   U17689 : OAI22_X1 port map( A1 => n21961, A2 => n22516, B1 => n21956, B2 => 
                           n16463, ZN => n5972);
   U17690 : OAI22_X1 port map( A1 => n21961, A2 => n22522, B1 => n21956, B2 => 
                           n16462, ZN => n5973);
   U17691 : OAI22_X1 port map( A1 => n21966, A2 => n22382, B1 => n21965, B2 => 
                           n16451, ZN => n5982);
   U17692 : OAI22_X1 port map( A1 => n21966, A2 => n22390, B1 => n21965, B2 => 
                           n16450, ZN => n5983);
   U17693 : OAI22_X1 port map( A1 => n21966, A2 => n22396, B1 => n21965, B2 => 
                           n16449, ZN => n5984);
   U17694 : OAI22_X1 port map( A1 => n21966, A2 => n22402, B1 => n21965, B2 => 
                           n16448, ZN => n5985);
   U17695 : OAI22_X1 port map( A1 => n21966, A2 => n22408, B1 => n21965, B2 => 
                           n16447, ZN => n5986);
   U17696 : OAI22_X1 port map( A1 => n21967, A2 => n22414, B1 => n21965, B2 => 
                           n16446, ZN => n5987);
   U17697 : OAI22_X1 port map( A1 => n21967, A2 => n22420, B1 => n21965, B2 => 
                           n16445, ZN => n5988);
   U17698 : OAI22_X1 port map( A1 => n21967, A2 => n22426, B1 => n21965, B2 => 
                           n16444, ZN => n5989);
   U17699 : OAI22_X1 port map( A1 => n21967, A2 => n22432, B1 => n21965, B2 => 
                           n16443, ZN => n5990);
   U17700 : OAI22_X1 port map( A1 => n21967, A2 => n22438, B1 => n21965, B2 => 
                           n16442, ZN => n5991);
   U17701 : OAI22_X1 port map( A1 => n21968, A2 => n22444, B1 => n21965, B2 => 
                           n16441, ZN => n5992);
   U17702 : OAI22_X1 port map( A1 => n21968, A2 => n22450, B1 => n21965, B2 => 
                           n16440, ZN => n5993);
   U17703 : OAI22_X1 port map( A1 => n21968, A2 => n22456, B1 => n21965, B2 => 
                           n16439, ZN => n5994);
   U17704 : OAI22_X1 port map( A1 => n21968, A2 => n22462, B1 => n21965, B2 => 
                           n16438, ZN => n5995);
   U17705 : OAI22_X1 port map( A1 => n21968, A2 => n22468, B1 => n16419, B2 => 
                           n16437, ZN => n5996);
   U17706 : OAI22_X1 port map( A1 => n21969, A2 => n22474, B1 => n16419, B2 => 
                           n16436, ZN => n5997);
   U17707 : OAI22_X1 port map( A1 => n21969, A2 => n22480, B1 => n16419, B2 => 
                           n16435, ZN => n5998);
   U17708 : OAI22_X1 port map( A1 => n21969, A2 => n22486, B1 => n16419, B2 => 
                           n16434, ZN => n5999);
   U17709 : OAI22_X1 port map( A1 => n21969, A2 => n22492, B1 => n16419, B2 => 
                           n16433, ZN => n6000);
   U17710 : OAI22_X1 port map( A1 => n21969, A2 => n22498, B1 => n16419, B2 => 
                           n16432, ZN => n6001);
   U17711 : OAI22_X1 port map( A1 => n21970, A2 => n22504, B1 => n16419, B2 => 
                           n16431, ZN => n6002);
   U17712 : OAI22_X1 port map( A1 => n21970, A2 => n22510, B1 => n21965, B2 => 
                           n16430, ZN => n6003);
   U17713 : OAI22_X1 port map( A1 => n21970, A2 => n22516, B1 => n21965, B2 => 
                           n16429, ZN => n6004);
   U17714 : OAI22_X1 port map( A1 => n21970, A2 => n22522, B1 => n21965, B2 => 
                           n16428, ZN => n6005);
   U17715 : OAI22_X1 port map( A1 => n21975, A2 => n22382, B1 => n21974, B2 => 
                           n16416, ZN => n6014);
   U17716 : OAI22_X1 port map( A1 => n21975, A2 => n22390, B1 => n21974, B2 => 
                           n16415, ZN => n6015);
   U17717 : OAI22_X1 port map( A1 => n21975, A2 => n22396, B1 => n21974, B2 => 
                           n16414, ZN => n6016);
   U17718 : OAI22_X1 port map( A1 => n21975, A2 => n22402, B1 => n21974, B2 => 
                           n16413, ZN => n6017);
   U17719 : OAI22_X1 port map( A1 => n21975, A2 => n22408, B1 => n21974, B2 => 
                           n16412, ZN => n6018);
   U17720 : OAI22_X1 port map( A1 => n21976, A2 => n22414, B1 => n21974, B2 => 
                           n16411, ZN => n6019);
   U17721 : OAI22_X1 port map( A1 => n21976, A2 => n22420, B1 => n21974, B2 => 
                           n16410, ZN => n6020);
   U17722 : OAI22_X1 port map( A1 => n21976, A2 => n22426, B1 => n21974, B2 => 
                           n16409, ZN => n6021);
   U17723 : OAI22_X1 port map( A1 => n21976, A2 => n22432, B1 => n21974, B2 => 
                           n16408, ZN => n6022);
   U17724 : OAI22_X1 port map( A1 => n21976, A2 => n22438, B1 => n21974, B2 => 
                           n16407, ZN => n6023);
   U17725 : OAI22_X1 port map( A1 => n21977, A2 => n22444, B1 => n21974, B2 => 
                           n16406, ZN => n6024);
   U17726 : OAI22_X1 port map( A1 => n21977, A2 => n22450, B1 => n21974, B2 => 
                           n16405, ZN => n6025);
   U17727 : OAI22_X1 port map( A1 => n21977, A2 => n22456, B1 => n21974, B2 => 
                           n16404, ZN => n6026);
   U17728 : OAI22_X1 port map( A1 => n21977, A2 => n22462, B1 => n21974, B2 => 
                           n16403, ZN => n6027);
   U17729 : OAI22_X1 port map( A1 => n21977, A2 => n22468, B1 => n16384, B2 => 
                           n16402, ZN => n6028);
   U17730 : OAI22_X1 port map( A1 => n21978, A2 => n22474, B1 => n16384, B2 => 
                           n16401, ZN => n6029);
   U17731 : OAI22_X1 port map( A1 => n21978, A2 => n22480, B1 => n16384, B2 => 
                           n16400, ZN => n6030);
   U17732 : OAI22_X1 port map( A1 => n21978, A2 => n22486, B1 => n16384, B2 => 
                           n16399, ZN => n6031);
   U17733 : OAI22_X1 port map( A1 => n21978, A2 => n22492, B1 => n16384, B2 => 
                           n16398, ZN => n6032);
   U17734 : OAI22_X1 port map( A1 => n21978, A2 => n22498, B1 => n16384, B2 => 
                           n16397, ZN => n6033);
   U17735 : OAI22_X1 port map( A1 => n21979, A2 => n22504, B1 => n16384, B2 => 
                           n16396, ZN => n6034);
   U17736 : OAI22_X1 port map( A1 => n21979, A2 => n22510, B1 => n21974, B2 => 
                           n16395, ZN => n6035);
   U17737 : OAI22_X1 port map( A1 => n21979, A2 => n22516, B1 => n21974, B2 => 
                           n16394, ZN => n6036);
   U17738 : OAI22_X1 port map( A1 => n21979, A2 => n22522, B1 => n21974, B2 => 
                           n16393, ZN => n6037);
   U17739 : OAI22_X1 port map( A1 => n22029, A2 => n22383, B1 => n22028, B2 => 
                           n16307, ZN => n6206);
   U17740 : OAI22_X1 port map( A1 => n22029, A2 => n22390, B1 => n22028, B2 => 
                           n16306, ZN => n6207);
   U17741 : OAI22_X1 port map( A1 => n22029, A2 => n22396, B1 => n22028, B2 => 
                           n16305, ZN => n6208);
   U17742 : OAI22_X1 port map( A1 => n22029, A2 => n22402, B1 => n22028, B2 => 
                           n16304, ZN => n6209);
   U17743 : OAI22_X1 port map( A1 => n22029, A2 => n22408, B1 => n22028, B2 => 
                           n16303, ZN => n6210);
   U17744 : OAI22_X1 port map( A1 => n22030, A2 => n22414, B1 => n22028, B2 => 
                           n16302, ZN => n6211);
   U17745 : OAI22_X1 port map( A1 => n22030, A2 => n22420, B1 => n22028, B2 => 
                           n16301, ZN => n6212);
   U17746 : OAI22_X1 port map( A1 => n22030, A2 => n22426, B1 => n22028, B2 => 
                           n16300, ZN => n6213);
   U17747 : OAI22_X1 port map( A1 => n22030, A2 => n22432, B1 => n22028, B2 => 
                           n16299, ZN => n6214);
   U17748 : OAI22_X1 port map( A1 => n22030, A2 => n22438, B1 => n22028, B2 => 
                           n16298, ZN => n6215);
   U17749 : OAI22_X1 port map( A1 => n22031, A2 => n22444, B1 => n22028, B2 => 
                           n16297, ZN => n6216);
   U17750 : OAI22_X1 port map( A1 => n22031, A2 => n22450, B1 => n22028, B2 => 
                           n16296, ZN => n6217);
   U17751 : OAI22_X1 port map( A1 => n22031, A2 => n22456, B1 => n22028, B2 => 
                           n16295, ZN => n6218);
   U17752 : OAI22_X1 port map( A1 => n22031, A2 => n22462, B1 => n22028, B2 => 
                           n16294, ZN => n6219);
   U17753 : OAI22_X1 port map( A1 => n22031, A2 => n22468, B1 => n16275, B2 => 
                           n16293, ZN => n6220);
   U17754 : OAI22_X1 port map( A1 => n22032, A2 => n22474, B1 => n16275, B2 => 
                           n16292, ZN => n6221);
   U17755 : OAI22_X1 port map( A1 => n22032, A2 => n22480, B1 => n16275, B2 => 
                           n16291, ZN => n6222);
   U17756 : OAI22_X1 port map( A1 => n22032, A2 => n22486, B1 => n16275, B2 => 
                           n16290, ZN => n6223);
   U17757 : OAI22_X1 port map( A1 => n22032, A2 => n22492, B1 => n16275, B2 => 
                           n16289, ZN => n6224);
   U17758 : OAI22_X1 port map( A1 => n22032, A2 => n22498, B1 => n16275, B2 => 
                           n16288, ZN => n6225);
   U17759 : OAI22_X1 port map( A1 => n22033, A2 => n22504, B1 => n16275, B2 => 
                           n16287, ZN => n6226);
   U17760 : OAI22_X1 port map( A1 => n22033, A2 => n22510, B1 => n22028, B2 => 
                           n16286, ZN => n6227);
   U17761 : OAI22_X1 port map( A1 => n22033, A2 => n22516, B1 => n22028, B2 => 
                           n16285, ZN => n6228);
   U17762 : OAI22_X1 port map( A1 => n22033, A2 => n22522, B1 => n22028, B2 => 
                           n16284, ZN => n6229);
   U17763 : OAI22_X1 port map( A1 => n22110, A2 => n22383, B1 => n22109, B2 => 
                           n20048, ZN => n6494);
   U17764 : OAI22_X1 port map( A1 => n22110, A2 => n22389, B1 => n22109, B2 => 
                           n20049, ZN => n6495);
   U17765 : OAI22_X1 port map( A1 => n22110, A2 => n22395, B1 => n22109, B2 => 
                           n20050, ZN => n6496);
   U17766 : OAI22_X1 port map( A1 => n22110, A2 => n22401, B1 => n22109, B2 => 
                           n20051, ZN => n6497);
   U17767 : OAI22_X1 port map( A1 => n22110, A2 => n22407, B1 => n22109, B2 => 
                           n20052, ZN => n6498);
   U17768 : OAI22_X1 port map( A1 => n22111, A2 => n22413, B1 => n22109, B2 => 
                           n20053, ZN => n6499);
   U17769 : OAI22_X1 port map( A1 => n22111, A2 => n22419, B1 => n22109, B2 => 
                           n20054, ZN => n6500);
   U17770 : OAI22_X1 port map( A1 => n22111, A2 => n22425, B1 => n22109, B2 => 
                           n20055, ZN => n6501);
   U17771 : OAI22_X1 port map( A1 => n22111, A2 => n22431, B1 => n22109, B2 => 
                           n20056, ZN => n6502);
   U17772 : OAI22_X1 port map( A1 => n22111, A2 => n22437, B1 => n22109, B2 => 
                           n20057, ZN => n6503);
   U17773 : OAI22_X1 port map( A1 => n22112, A2 => n22443, B1 => n22109, B2 => 
                           n20058, ZN => n6504);
   U17774 : OAI22_X1 port map( A1 => n22112, A2 => n22449, B1 => n22109, B2 => 
                           n20059, ZN => n6505);
   U17775 : OAI22_X1 port map( A1 => n22112, A2 => n22455, B1 => n22109, B2 => 
                           n20060, ZN => n6506);
   U17776 : OAI22_X1 port map( A1 => n22112, A2 => n22461, B1 => n22109, B2 => 
                           n20061, ZN => n6507);
   U17777 : OAI22_X1 port map( A1 => n22112, A2 => n22467, B1 => n15998, B2 => 
                           n20062, ZN => n6508);
   U17778 : OAI22_X1 port map( A1 => n22113, A2 => n22473, B1 => n15998, B2 => 
                           n20063, ZN => n6509);
   U17779 : OAI22_X1 port map( A1 => n22113, A2 => n22479, B1 => n15998, B2 => 
                           n20064, ZN => n6510);
   U17780 : OAI22_X1 port map( A1 => n22113, A2 => n22485, B1 => n15998, B2 => 
                           n20065, ZN => n6511);
   U17781 : OAI22_X1 port map( A1 => n22113, A2 => n22491, B1 => n15998, B2 => 
                           n20066, ZN => n6512);
   U17782 : OAI22_X1 port map( A1 => n22113, A2 => n22497, B1 => n15998, B2 => 
                           n20067, ZN => n6513);
   U17783 : OAI22_X1 port map( A1 => n22114, A2 => n22503, B1 => n15998, B2 => 
                           n20068, ZN => n6514);
   U17784 : OAI22_X1 port map( A1 => n22114, A2 => n22509, B1 => n22109, B2 => 
                           n20069, ZN => n6515);
   U17785 : OAI22_X1 port map( A1 => n22114, A2 => n22515, B1 => n22109, B2 => 
                           n20070, ZN => n6516);
   U17786 : OAI22_X1 port map( A1 => n22114, A2 => n22521, B1 => n22109, B2 => 
                           n20071, ZN => n6517);
   U17787 : OAI22_X1 port map( A1 => n22119, A2 => n22383, B1 => n22118, B2 => 
                           n20072, ZN => n6526);
   U17788 : OAI22_X1 port map( A1 => n22119, A2 => n22389, B1 => n22118, B2 => 
                           n20073, ZN => n6527);
   U17789 : OAI22_X1 port map( A1 => n22119, A2 => n22395, B1 => n22118, B2 => 
                           n20074, ZN => n6528);
   U17790 : OAI22_X1 port map( A1 => n22119, A2 => n22401, B1 => n22118, B2 => 
                           n20075, ZN => n6529);
   U17791 : OAI22_X1 port map( A1 => n22119, A2 => n22407, B1 => n22118, B2 => 
                           n20076, ZN => n6530);
   U17792 : OAI22_X1 port map( A1 => n22120, A2 => n22413, B1 => n22118, B2 => 
                           n20077, ZN => n6531);
   U17793 : OAI22_X1 port map( A1 => n22120, A2 => n22419, B1 => n22118, B2 => 
                           n20078, ZN => n6532);
   U17794 : OAI22_X1 port map( A1 => n22120, A2 => n22425, B1 => n22118, B2 => 
                           n20079, ZN => n6533);
   U17795 : OAI22_X1 port map( A1 => n22120, A2 => n22431, B1 => n22118, B2 => 
                           n20080, ZN => n6534);
   U17796 : OAI22_X1 port map( A1 => n22120, A2 => n22437, B1 => n22118, B2 => 
                           n20081, ZN => n6535);
   U17797 : OAI22_X1 port map( A1 => n22121, A2 => n22443, B1 => n22118, B2 => 
                           n20082, ZN => n6536);
   U17798 : OAI22_X1 port map( A1 => n22121, A2 => n22449, B1 => n22118, B2 => 
                           n20083, ZN => n6537);
   U17799 : OAI22_X1 port map( A1 => n22121, A2 => n22455, B1 => n22118, B2 => 
                           n20084, ZN => n6538);
   U17800 : OAI22_X1 port map( A1 => n22121, A2 => n22461, B1 => n22118, B2 => 
                           n20085, ZN => n6539);
   U17801 : OAI22_X1 port map( A1 => n22121, A2 => n22467, B1 => n15963, B2 => 
                           n20086, ZN => n6540);
   U17802 : OAI22_X1 port map( A1 => n22122, A2 => n22473, B1 => n15963, B2 => 
                           n20087, ZN => n6541);
   U17803 : OAI22_X1 port map( A1 => n22122, A2 => n22479, B1 => n15963, B2 => 
                           n20088, ZN => n6542);
   U17804 : OAI22_X1 port map( A1 => n22122, A2 => n22485, B1 => n15963, B2 => 
                           n20089, ZN => n6543);
   U17805 : OAI22_X1 port map( A1 => n22122, A2 => n22491, B1 => n15963, B2 => 
                           n20090, ZN => n6544);
   U17806 : OAI22_X1 port map( A1 => n22122, A2 => n22497, B1 => n15963, B2 => 
                           n20091, ZN => n6545);
   U17807 : OAI22_X1 port map( A1 => n22123, A2 => n22503, B1 => n15963, B2 => 
                           n20092, ZN => n6546);
   U17808 : OAI22_X1 port map( A1 => n22123, A2 => n22509, B1 => n22118, B2 => 
                           n20093, ZN => n6547);
   U17809 : OAI22_X1 port map( A1 => n22123, A2 => n22515, B1 => n22118, B2 => 
                           n20094, ZN => n6548);
   U17810 : OAI22_X1 port map( A1 => n22123, A2 => n22521, B1 => n22118, B2 => 
                           n20095, ZN => n6549);
   U17811 : OAI22_X1 port map( A1 => n22128, A2 => n22384, B1 => n22127, B2 => 
                           n15961, ZN => n6558);
   U17812 : OAI22_X1 port map( A1 => n22128, A2 => n22389, B1 => n22127, B2 => 
                           n15960, ZN => n6559);
   U17813 : OAI22_X1 port map( A1 => n22128, A2 => n22395, B1 => n22127, B2 => 
                           n15959, ZN => n6560);
   U17814 : OAI22_X1 port map( A1 => n22128, A2 => n22401, B1 => n22127, B2 => 
                           n15958, ZN => n6561);
   U17815 : OAI22_X1 port map( A1 => n22128, A2 => n22407, B1 => n22127, B2 => 
                           n15957, ZN => n6562);
   U17816 : OAI22_X1 port map( A1 => n22129, A2 => n22413, B1 => n22127, B2 => 
                           n15956, ZN => n6563);
   U17817 : OAI22_X1 port map( A1 => n22129, A2 => n22419, B1 => n22127, B2 => 
                           n15955, ZN => n6564);
   U17818 : OAI22_X1 port map( A1 => n22129, A2 => n22425, B1 => n22127, B2 => 
                           n15954, ZN => n6565);
   U17819 : OAI22_X1 port map( A1 => n22129, A2 => n22431, B1 => n22127, B2 => 
                           n15953, ZN => n6566);
   U17820 : OAI22_X1 port map( A1 => n22129, A2 => n22437, B1 => n22127, B2 => 
                           n15952, ZN => n6567);
   U17821 : OAI22_X1 port map( A1 => n22130, A2 => n22443, B1 => n22127, B2 => 
                           n15951, ZN => n6568);
   U17822 : OAI22_X1 port map( A1 => n22130, A2 => n22449, B1 => n22127, B2 => 
                           n15950, ZN => n6569);
   U17823 : OAI22_X1 port map( A1 => n22130, A2 => n22455, B1 => n22127, B2 => 
                           n15949, ZN => n6570);
   U17824 : OAI22_X1 port map( A1 => n22130, A2 => n22461, B1 => n22127, B2 => 
                           n15948, ZN => n6571);
   U17825 : OAI22_X1 port map( A1 => n22130, A2 => n22467, B1 => n15929, B2 => 
                           n15947, ZN => n6572);
   U17826 : OAI22_X1 port map( A1 => n22131, A2 => n22473, B1 => n15929, B2 => 
                           n15946, ZN => n6573);
   U17827 : OAI22_X1 port map( A1 => n22131, A2 => n22479, B1 => n15929, B2 => 
                           n15945, ZN => n6574);
   U17828 : OAI22_X1 port map( A1 => n22131, A2 => n22485, B1 => n15929, B2 => 
                           n15944, ZN => n6575);
   U17829 : OAI22_X1 port map( A1 => n22131, A2 => n22491, B1 => n15929, B2 => 
                           n15943, ZN => n6576);
   U17830 : OAI22_X1 port map( A1 => n22131, A2 => n22497, B1 => n15929, B2 => 
                           n15942, ZN => n6577);
   U17831 : OAI22_X1 port map( A1 => n22132, A2 => n22503, B1 => n15929, B2 => 
                           n15941, ZN => n6578);
   U17832 : OAI22_X1 port map( A1 => n22132, A2 => n22509, B1 => n22127, B2 => 
                           n15940, ZN => n6579);
   U17833 : OAI22_X1 port map( A1 => n22132, A2 => n22515, B1 => n22127, B2 => 
                           n15939, ZN => n6580);
   U17834 : OAI22_X1 port map( A1 => n22132, A2 => n22521, B1 => n22127, B2 => 
                           n15938, ZN => n6581);
   U17835 : OAI22_X1 port map( A1 => n22164, A2 => n22384, B1 => n22163, B2 => 
                           n15888, ZN => n6686);
   U17836 : OAI22_X1 port map( A1 => n22164, A2 => n22388, B1 => n22163, B2 => 
                           n15887, ZN => n6687);
   U17837 : OAI22_X1 port map( A1 => n22164, A2 => n22394, B1 => n22163, B2 => 
                           n15886, ZN => n6688);
   U17838 : OAI22_X1 port map( A1 => n22164, A2 => n22400, B1 => n22163, B2 => 
                           n15885, ZN => n6689);
   U17839 : OAI22_X1 port map( A1 => n22164, A2 => n22406, B1 => n22163, B2 => 
                           n15884, ZN => n6690);
   U17840 : OAI22_X1 port map( A1 => n22165, A2 => n22412, B1 => n22163, B2 => 
                           n15883, ZN => n6691);
   U17841 : OAI22_X1 port map( A1 => n22165, A2 => n22418, B1 => n22163, B2 => 
                           n15882, ZN => n6692);
   U17842 : OAI22_X1 port map( A1 => n22165, A2 => n22424, B1 => n22163, B2 => 
                           n15881, ZN => n6693);
   U17843 : OAI22_X1 port map( A1 => n22165, A2 => n22430, B1 => n22163, B2 => 
                           n15880, ZN => n6694);
   U17844 : OAI22_X1 port map( A1 => n22165, A2 => n22436, B1 => n22163, B2 => 
                           n15879, ZN => n6695);
   U17845 : OAI22_X1 port map( A1 => n22166, A2 => n22442, B1 => n22163, B2 => 
                           n15878, ZN => n6696);
   U17846 : OAI22_X1 port map( A1 => n22166, A2 => n22448, B1 => n22163, B2 => 
                           n15877, ZN => n6697);
   U17847 : OAI22_X1 port map( A1 => n22166, A2 => n22454, B1 => n22163, B2 => 
                           n15876, ZN => n6698);
   U17848 : OAI22_X1 port map( A1 => n22166, A2 => n22460, B1 => n22163, B2 => 
                           n15875, ZN => n6699);
   U17849 : OAI22_X1 port map( A1 => n22166, A2 => n22466, B1 => n15856, B2 => 
                           n15874, ZN => n6700);
   U17850 : OAI22_X1 port map( A1 => n22167, A2 => n22472, B1 => n15856, B2 => 
                           n15873, ZN => n6701);
   U17851 : OAI22_X1 port map( A1 => n22167, A2 => n22478, B1 => n15856, B2 => 
                           n15872, ZN => n6702);
   U17852 : OAI22_X1 port map( A1 => n22167, A2 => n22484, B1 => n15856, B2 => 
                           n15871, ZN => n6703);
   U17853 : OAI22_X1 port map( A1 => n22167, A2 => n22490, B1 => n15856, B2 => 
                           n15870, ZN => n6704);
   U17854 : OAI22_X1 port map( A1 => n22167, A2 => n22496, B1 => n15856, B2 => 
                           n15869, ZN => n6705);
   U17855 : OAI22_X1 port map( A1 => n22168, A2 => n22502, B1 => n15856, B2 => 
                           n15868, ZN => n6706);
   U17856 : OAI22_X1 port map( A1 => n22168, A2 => n22508, B1 => n22163, B2 => 
                           n15867, ZN => n6707);
   U17857 : OAI22_X1 port map( A1 => n22168, A2 => n22514, B1 => n22163, B2 => 
                           n15866, ZN => n6708);
   U17858 : OAI22_X1 port map( A1 => n22168, A2 => n22520, B1 => n22163, B2 => 
                           n15865, ZN => n6709);
   U17859 : OAI22_X1 port map( A1 => n22209, A2 => n22384, B1 => n22208, B2 => 
                           n15748, ZN => n6846);
   U17860 : OAI22_X1 port map( A1 => n22209, A2 => n22388, B1 => n22208, B2 => 
                           n20120, ZN => n6847);
   U17861 : OAI22_X1 port map( A1 => n22209, A2 => n22394, B1 => n22208, B2 => 
                           n20121, ZN => n6848);
   U17862 : OAI22_X1 port map( A1 => n22209, A2 => n22400, B1 => n22208, B2 => 
                           n20122, ZN => n6849);
   U17863 : OAI22_X1 port map( A1 => n22209, A2 => n22406, B1 => n22208, B2 => 
                           n20123, ZN => n6850);
   U17864 : OAI22_X1 port map( A1 => n22210, A2 => n22412, B1 => n22208, B2 => 
                           n20124, ZN => n6851);
   U17865 : OAI22_X1 port map( A1 => n22210, A2 => n22418, B1 => n22208, B2 => 
                           n20125, ZN => n6852);
   U17866 : OAI22_X1 port map( A1 => n22210, A2 => n22424, B1 => n22208, B2 => 
                           n20126, ZN => n6853);
   U17867 : OAI22_X1 port map( A1 => n22210, A2 => n22430, B1 => n22208, B2 => 
                           n20127, ZN => n6854);
   U17868 : OAI22_X1 port map( A1 => n22210, A2 => n22436, B1 => n22208, B2 => 
                           n20128, ZN => n6855);
   U17869 : OAI22_X1 port map( A1 => n22211, A2 => n22442, B1 => n22208, B2 => 
                           n20129, ZN => n6856);
   U17870 : OAI22_X1 port map( A1 => n22211, A2 => n22448, B1 => n22208, B2 => 
                           n20130, ZN => n6857);
   U17871 : OAI22_X1 port map( A1 => n22211, A2 => n22454, B1 => n22208, B2 => 
                           n20131, ZN => n6858);
   U17872 : OAI22_X1 port map( A1 => n22211, A2 => n22460, B1 => n22208, B2 => 
                           n20132, ZN => n6859);
   U17873 : OAI22_X1 port map( A1 => n22211, A2 => n22466, B1 => n15716, B2 => 
                           n20133, ZN => n6860);
   U17874 : OAI22_X1 port map( A1 => n22212, A2 => n22472, B1 => n15716, B2 => 
                           n20134, ZN => n6861);
   U17875 : OAI22_X1 port map( A1 => n22212, A2 => n22478, B1 => n15716, B2 => 
                           n20135, ZN => n6862);
   U17876 : OAI22_X1 port map( A1 => n22212, A2 => n22484, B1 => n15716, B2 => 
                           n20136, ZN => n6863);
   U17877 : OAI22_X1 port map( A1 => n22212, A2 => n22490, B1 => n15716, B2 => 
                           n20137, ZN => n6864);
   U17878 : OAI22_X1 port map( A1 => n22212, A2 => n22496, B1 => n15716, B2 => 
                           n20138, ZN => n6865);
   U17879 : OAI22_X1 port map( A1 => n22213, A2 => n22502, B1 => n15716, B2 => 
                           n20139, ZN => n6866);
   U17880 : OAI22_X1 port map( A1 => n22213, A2 => n22508, B1 => n22208, B2 => 
                           n20140, ZN => n6867);
   U17881 : OAI22_X1 port map( A1 => n22213, A2 => n22514, B1 => n22208, B2 => 
                           n20141, ZN => n6868);
   U17882 : OAI22_X1 port map( A1 => n22213, A2 => n22520, B1 => n22208, B2 => 
                           n20142, ZN => n6869);
   U17883 : OAI22_X1 port map( A1 => n22236, A2 => n22385, B1 => n22235, B2 => 
                           n15641, ZN => n6942);
   U17884 : OAI22_X1 port map( A1 => n22236, A2 => n22388, B1 => n22235, B2 => 
                           n20143, ZN => n6943);
   U17885 : OAI22_X1 port map( A1 => n22236, A2 => n22394, B1 => n22235, B2 => 
                           n20144, ZN => n6944);
   U17886 : OAI22_X1 port map( A1 => n22236, A2 => n22400, B1 => n22235, B2 => 
                           n20145, ZN => n6945);
   U17887 : OAI22_X1 port map( A1 => n22236, A2 => n22406, B1 => n22235, B2 => 
                           n20146, ZN => n6946);
   U17888 : OAI22_X1 port map( A1 => n22237, A2 => n22412, B1 => n22235, B2 => 
                           n20147, ZN => n6947);
   U17889 : OAI22_X1 port map( A1 => n22237, A2 => n22418, B1 => n22235, B2 => 
                           n20148, ZN => n6948);
   U17890 : OAI22_X1 port map( A1 => n22237, A2 => n22424, B1 => n22235, B2 => 
                           n20149, ZN => n6949);
   U17891 : OAI22_X1 port map( A1 => n22237, A2 => n22430, B1 => n22235, B2 => 
                           n20150, ZN => n6950);
   U17892 : OAI22_X1 port map( A1 => n22237, A2 => n22436, B1 => n22235, B2 => 
                           n20151, ZN => n6951);
   U17893 : OAI22_X1 port map( A1 => n22238, A2 => n22442, B1 => n22235, B2 => 
                           n20152, ZN => n6952);
   U17894 : OAI22_X1 port map( A1 => n22238, A2 => n22448, B1 => n22235, B2 => 
                           n20153, ZN => n6953);
   U17895 : OAI22_X1 port map( A1 => n22238, A2 => n22454, B1 => n22235, B2 => 
                           n20154, ZN => n6954);
   U17896 : OAI22_X1 port map( A1 => n22238, A2 => n22460, B1 => n22235, B2 => 
                           n20155, ZN => n6955);
   U17897 : OAI22_X1 port map( A1 => n22238, A2 => n22466, B1 => n15609, B2 => 
                           n20156, ZN => n6956);
   U17898 : OAI22_X1 port map( A1 => n22239, A2 => n22472, B1 => n15609, B2 => 
                           n20157, ZN => n6957);
   U17899 : OAI22_X1 port map( A1 => n22239, A2 => n22478, B1 => n15609, B2 => 
                           n20158, ZN => n6958);
   U17900 : OAI22_X1 port map( A1 => n22239, A2 => n22484, B1 => n15609, B2 => 
                           n20159, ZN => n6959);
   U17901 : OAI22_X1 port map( A1 => n22239, A2 => n22490, B1 => n15609, B2 => 
                           n20160, ZN => n6960);
   U17902 : OAI22_X1 port map( A1 => n22239, A2 => n22496, B1 => n15609, B2 => 
                           n20161, ZN => n6961);
   U17903 : OAI22_X1 port map( A1 => n22240, A2 => n22502, B1 => n15609, B2 => 
                           n20162, ZN => n6962);
   U17904 : OAI22_X1 port map( A1 => n22240, A2 => n22508, B1 => n22235, B2 => 
                           n20163, ZN => n6963);
   U17905 : OAI22_X1 port map( A1 => n22240, A2 => n22514, B1 => n22235, B2 => 
                           n20164, ZN => n6964);
   U17906 : OAI22_X1 port map( A1 => n22240, A2 => n22520, B1 => n22235, B2 => 
                           n20165, ZN => n6965);
   U17907 : OAI22_X1 port map( A1 => n22254, A2 => n22385, B1 => n22253, B2 => 
                           n20260, ZN => n7006);
   U17908 : OAI22_X1 port map( A1 => n22254, A2 => n22388, B1 => n22253, B2 => 
                           n20261, ZN => n7007);
   U17909 : OAI22_X1 port map( A1 => n22254, A2 => n22394, B1 => n22253, B2 => 
                           n20262, ZN => n7008);
   U17910 : OAI22_X1 port map( A1 => n22254, A2 => n22400, B1 => n22253, B2 => 
                           n20263, ZN => n7009);
   U17911 : OAI22_X1 port map( A1 => n22254, A2 => n22406, B1 => n22253, B2 => 
                           n20264, ZN => n7010);
   U17912 : OAI22_X1 port map( A1 => n22255, A2 => n22412, B1 => n22253, B2 => 
                           n20265, ZN => n7011);
   U17913 : OAI22_X1 port map( A1 => n22255, A2 => n22418, B1 => n22253, B2 => 
                           n20266, ZN => n7012);
   U17914 : OAI22_X1 port map( A1 => n22255, A2 => n22424, B1 => n22253, B2 => 
                           n20267, ZN => n7013);
   U17915 : OAI22_X1 port map( A1 => n22255, A2 => n22430, B1 => n22253, B2 => 
                           n20268, ZN => n7014);
   U17916 : OAI22_X1 port map( A1 => n22255, A2 => n22436, B1 => n22253, B2 => 
                           n20269, ZN => n7015);
   U17917 : OAI22_X1 port map( A1 => n22256, A2 => n22442, B1 => n22253, B2 => 
                           n20270, ZN => n7016);
   U17918 : OAI22_X1 port map( A1 => n22256, A2 => n22448, B1 => n22253, B2 => 
                           n20271, ZN => n7017);
   U17919 : OAI22_X1 port map( A1 => n22256, A2 => n22454, B1 => n22253, B2 => 
                           n20272, ZN => n7018);
   U17920 : OAI22_X1 port map( A1 => n22256, A2 => n22460, B1 => n22253, B2 => 
                           n20273, ZN => n7019);
   U17921 : OAI22_X1 port map( A1 => n22256, A2 => n22466, B1 => n15541, B2 => 
                           n20274, ZN => n7020);
   U17922 : OAI22_X1 port map( A1 => n22257, A2 => n22472, B1 => n15541, B2 => 
                           n20275, ZN => n7021);
   U17923 : OAI22_X1 port map( A1 => n22257, A2 => n22478, B1 => n15541, B2 => 
                           n20276, ZN => n7022);
   U17924 : OAI22_X1 port map( A1 => n22257, A2 => n22484, B1 => n15541, B2 => 
                           n20277, ZN => n7023);
   U17925 : OAI22_X1 port map( A1 => n22257, A2 => n22490, B1 => n15541, B2 => 
                           n20278, ZN => n7024);
   U17926 : OAI22_X1 port map( A1 => n22257, A2 => n22496, B1 => n15541, B2 => 
                           n20279, ZN => n7025);
   U17927 : OAI22_X1 port map( A1 => n22258, A2 => n22502, B1 => n15541, B2 => 
                           n20280, ZN => n7026);
   U17928 : OAI22_X1 port map( A1 => n22258, A2 => n22508, B1 => n22253, B2 => 
                           n20281, ZN => n7027);
   U17929 : OAI22_X1 port map( A1 => n22258, A2 => n22514, B1 => n22253, B2 => 
                           n20282, ZN => n7028);
   U17930 : OAI22_X1 port map( A1 => n22258, A2 => n22520, B1 => n22253, B2 => 
                           n20283, ZN => n7029);
   U17931 : OAI22_X1 port map( A1 => n22263, A2 => n22385, B1 => n22262, B2 => 
                           n20284, ZN => n7038);
   U17932 : OAI22_X1 port map( A1 => n22263, A2 => n22388, B1 => n22262, B2 => 
                           n20285, ZN => n7039);
   U17933 : OAI22_X1 port map( A1 => n22263, A2 => n22394, B1 => n22262, B2 => 
                           n20286, ZN => n7040);
   U17934 : OAI22_X1 port map( A1 => n22263, A2 => n22400, B1 => n22262, B2 => 
                           n20287, ZN => n7041);
   U17935 : OAI22_X1 port map( A1 => n22263, A2 => n22406, B1 => n22262, B2 => 
                           n20288, ZN => n7042);
   U17936 : OAI22_X1 port map( A1 => n22264, A2 => n22412, B1 => n22262, B2 => 
                           n20289, ZN => n7043);
   U17937 : OAI22_X1 port map( A1 => n22264, A2 => n22418, B1 => n22262, B2 => 
                           n20290, ZN => n7044);
   U17938 : OAI22_X1 port map( A1 => n22264, A2 => n22424, B1 => n22262, B2 => 
                           n20291, ZN => n7045);
   U17939 : OAI22_X1 port map( A1 => n22264, A2 => n22430, B1 => n22262, B2 => 
                           n20292, ZN => n7046);
   U17940 : OAI22_X1 port map( A1 => n22264, A2 => n22436, B1 => n22262, B2 => 
                           n20293, ZN => n7047);
   U17941 : OAI22_X1 port map( A1 => n22265, A2 => n22442, B1 => n22262, B2 => 
                           n20294, ZN => n7048);
   U17942 : OAI22_X1 port map( A1 => n22265, A2 => n22448, B1 => n22262, B2 => 
                           n20295, ZN => n7049);
   U17943 : OAI22_X1 port map( A1 => n22265, A2 => n22454, B1 => n22262, B2 => 
                           n20296, ZN => n7050);
   U17944 : OAI22_X1 port map( A1 => n22265, A2 => n22460, B1 => n22262, B2 => 
                           n20297, ZN => n7051);
   U17945 : OAI22_X1 port map( A1 => n22265, A2 => n22466, B1 => n15506, B2 => 
                           n20298, ZN => n7052);
   U17946 : OAI22_X1 port map( A1 => n22266, A2 => n22472, B1 => n15506, B2 => 
                           n20299, ZN => n7053);
   U17947 : OAI22_X1 port map( A1 => n22266, A2 => n22478, B1 => n15506, B2 => 
                           n20300, ZN => n7054);
   U17948 : OAI22_X1 port map( A1 => n22266, A2 => n22484, B1 => n15506, B2 => 
                           n20301, ZN => n7055);
   U17949 : OAI22_X1 port map( A1 => n22266, A2 => n22490, B1 => n15506, B2 => 
                           n20302, ZN => n7056);
   U17950 : OAI22_X1 port map( A1 => n22266, A2 => n22496, B1 => n15506, B2 => 
                           n20303, ZN => n7057);
   U17951 : OAI22_X1 port map( A1 => n22267, A2 => n22502, B1 => n15506, B2 => 
                           n20304, ZN => n7058);
   U17952 : OAI22_X1 port map( A1 => n22267, A2 => n22508, B1 => n22262, B2 => 
                           n20305, ZN => n7059);
   U17953 : OAI22_X1 port map( A1 => n22267, A2 => n22514, B1 => n22262, B2 => 
                           n20306, ZN => n7060);
   U17954 : OAI22_X1 port map( A1 => n22267, A2 => n22520, B1 => n22262, B2 => 
                           n20307, ZN => n7061);
   U17955 : OAI22_X1 port map( A1 => n22308, A2 => n22385, B1 => n22307, B2 => 
                           n15365, ZN => n7198);
   U17956 : OAI22_X1 port map( A1 => n22308, A2 => n22387, B1 => n22307, B2 => 
                           n20023, ZN => n7199);
   U17957 : OAI22_X1 port map( A1 => n22308, A2 => n22393, B1 => n22307, B2 => 
                           n20024, ZN => n7200);
   U17958 : OAI22_X1 port map( A1 => n22308, A2 => n22399, B1 => n22307, B2 => 
                           n20025, ZN => n7201);
   U17959 : OAI22_X1 port map( A1 => n22308, A2 => n22405, B1 => n22307, B2 => 
                           n20026, ZN => n7202);
   U17960 : OAI22_X1 port map( A1 => n22309, A2 => n22411, B1 => n22307, B2 => 
                           n20027, ZN => n7203);
   U17961 : OAI22_X1 port map( A1 => n22309, A2 => n22417, B1 => n22307, B2 => 
                           n20028, ZN => n7204);
   U17962 : OAI22_X1 port map( A1 => n22309, A2 => n22423, B1 => n22307, B2 => 
                           n20029, ZN => n7205);
   U17963 : OAI22_X1 port map( A1 => n22309, A2 => n22429, B1 => n22307, B2 => 
                           n20030, ZN => n7206);
   U17964 : OAI22_X1 port map( A1 => n22309, A2 => n22435, B1 => n22307, B2 => 
                           n20031, ZN => n7207);
   U17965 : OAI22_X1 port map( A1 => n22310, A2 => n22441, B1 => n22307, B2 => 
                           n20032, ZN => n7208);
   U17966 : OAI22_X1 port map( A1 => n22310, A2 => n22447, B1 => n22307, B2 => 
                           n20033, ZN => n7209);
   U17967 : OAI22_X1 port map( A1 => n22310, A2 => n22453, B1 => n22307, B2 => 
                           n20034, ZN => n7210);
   U17968 : OAI22_X1 port map( A1 => n22310, A2 => n22459, B1 => n22307, B2 => 
                           n20035, ZN => n7211);
   U17969 : OAI22_X1 port map( A1 => n22310, A2 => n22465, B1 => n15333, B2 => 
                           n20036, ZN => n7212);
   U17970 : OAI22_X1 port map( A1 => n22311, A2 => n22471, B1 => n15333, B2 => 
                           n20037, ZN => n7213);
   U17971 : OAI22_X1 port map( A1 => n22311, A2 => n22477, B1 => n15333, B2 => 
                           n20038, ZN => n7214);
   U17972 : OAI22_X1 port map( A1 => n22311, A2 => n22483, B1 => n15333, B2 => 
                           n20039, ZN => n7215);
   U17973 : OAI22_X1 port map( A1 => n22311, A2 => n22489, B1 => n15333, B2 => 
                           n20040, ZN => n7216);
   U17974 : OAI22_X1 port map( A1 => n22311, A2 => n22495, B1 => n15333, B2 => 
                           n20041, ZN => n7217);
   U17975 : OAI22_X1 port map( A1 => n22312, A2 => n22501, B1 => n15333, B2 => 
                           n20042, ZN => n7218);
   U17976 : OAI22_X1 port map( A1 => n22312, A2 => n22507, B1 => n22307, B2 => 
                           n20043, ZN => n7219);
   U17977 : OAI22_X1 port map( A1 => n22312, A2 => n22513, B1 => n22307, B2 => 
                           n20044, ZN => n7220);
   U17978 : OAI22_X1 port map( A1 => n22312, A2 => n22519, B1 => n22307, B2 => 
                           n20045, ZN => n7221);
   U17979 : OAI22_X1 port map( A1 => n22317, A2 => n22385, B1 => n22316, B2 => 
                           n15331, ZN => n7230);
   U17980 : OAI22_X1 port map( A1 => n22317, A2 => n22387, B1 => n22316, B2 => 
                           n20166, ZN => n7231);
   U17981 : OAI22_X1 port map( A1 => n22317, A2 => n22393, B1 => n22316, B2 => 
                           n20167, ZN => n7232);
   U17982 : OAI22_X1 port map( A1 => n22317, A2 => n22399, B1 => n22316, B2 => 
                           n20168, ZN => n7233);
   U17983 : OAI22_X1 port map( A1 => n22317, A2 => n22405, B1 => n22316, B2 => 
                           n20169, ZN => n7234);
   U17984 : OAI22_X1 port map( A1 => n22318, A2 => n22411, B1 => n22316, B2 => 
                           n20170, ZN => n7235);
   U17985 : OAI22_X1 port map( A1 => n22318, A2 => n22417, B1 => n22316, B2 => 
                           n20171, ZN => n7236);
   U17986 : OAI22_X1 port map( A1 => n22318, A2 => n22423, B1 => n22316, B2 => 
                           n20172, ZN => n7237);
   U17987 : OAI22_X1 port map( A1 => n22318, A2 => n22429, B1 => n22316, B2 => 
                           n20173, ZN => n7238);
   U17988 : OAI22_X1 port map( A1 => n22318, A2 => n22435, B1 => n22316, B2 => 
                           n20174, ZN => n7239);
   U17989 : OAI22_X1 port map( A1 => n22319, A2 => n22441, B1 => n22316, B2 => 
                           n20175, ZN => n7240);
   U17990 : OAI22_X1 port map( A1 => n22319, A2 => n22447, B1 => n22316, B2 => 
                           n20176, ZN => n7241);
   U17991 : OAI22_X1 port map( A1 => n22319, A2 => n22453, B1 => n22316, B2 => 
                           n20177, ZN => n7242);
   U17992 : OAI22_X1 port map( A1 => n22319, A2 => n22459, B1 => n22316, B2 => 
                           n20178, ZN => n7243);
   U17993 : OAI22_X1 port map( A1 => n22319, A2 => n22465, B1 => n15299, B2 => 
                           n20179, ZN => n7244);
   U17994 : OAI22_X1 port map( A1 => n22320, A2 => n22471, B1 => n15299, B2 => 
                           n20180, ZN => n7245);
   U17995 : OAI22_X1 port map( A1 => n22320, A2 => n22477, B1 => n15299, B2 => 
                           n20181, ZN => n7246);
   U17996 : OAI22_X1 port map( A1 => n22320, A2 => n22483, B1 => n15299, B2 => 
                           n20182, ZN => n7247);
   U17997 : OAI22_X1 port map( A1 => n22320, A2 => n22489, B1 => n15299, B2 => 
                           n20183, ZN => n7248);
   U17998 : OAI22_X1 port map( A1 => n22320, A2 => n22495, B1 => n15299, B2 => 
                           n20184, ZN => n7249);
   U17999 : OAI22_X1 port map( A1 => n22321, A2 => n22501, B1 => n15299, B2 => 
                           n20185, ZN => n7250);
   U18000 : OAI22_X1 port map( A1 => n22321, A2 => n22507, B1 => n22316, B2 => 
                           n20186, ZN => n7251);
   U18001 : OAI22_X1 port map( A1 => n22321, A2 => n22513, B1 => n22316, B2 => 
                           n20187, ZN => n7252);
   U18002 : OAI22_X1 port map( A1 => n22321, A2 => n22519, B1 => n22316, B2 => 
                           n20188, ZN => n7253);
   U18003 : OAI22_X1 port map( A1 => n22344, A2 => n22386, B1 => n22343, B2 => 
                           n20096, ZN => n7326);
   U18004 : OAI22_X1 port map( A1 => n22344, A2 => n22387, B1 => n22343, B2 => 
                           n20189, ZN => n7327);
   U18005 : OAI22_X1 port map( A1 => n22344, A2 => n22393, B1 => n22343, B2 => 
                           n20190, ZN => n7328);
   U18006 : OAI22_X1 port map( A1 => n22344, A2 => n22399, B1 => n22343, B2 => 
                           n20191, ZN => n7329);
   U18007 : OAI22_X1 port map( A1 => n22344, A2 => n22405, B1 => n22343, B2 => 
                           n20192, ZN => n7330);
   U18008 : OAI22_X1 port map( A1 => n22345, A2 => n22411, B1 => n22343, B2 => 
                           n20193, ZN => n7331);
   U18009 : OAI22_X1 port map( A1 => n22345, A2 => n22417, B1 => n22343, B2 => 
                           n20194, ZN => n7332);
   U18010 : OAI22_X1 port map( A1 => n22345, A2 => n22423, B1 => n22343, B2 => 
                           n20195, ZN => n7333);
   U18011 : OAI22_X1 port map( A1 => n22345, A2 => n22429, B1 => n22343, B2 => 
                           n20196, ZN => n7334);
   U18012 : OAI22_X1 port map( A1 => n22345, A2 => n22435, B1 => n22343, B2 => 
                           n20197, ZN => n7335);
   U18013 : OAI22_X1 port map( A1 => n22346, A2 => n22441, B1 => n22343, B2 => 
                           n20198, ZN => n7336);
   U18014 : OAI22_X1 port map( A1 => n22346, A2 => n22447, B1 => n22343, B2 => 
                           n20199, ZN => n7337);
   U18015 : OAI22_X1 port map( A1 => n22346, A2 => n22453, B1 => n22343, B2 => 
                           n20200, ZN => n7338);
   U18016 : OAI22_X1 port map( A1 => n22346, A2 => n22459, B1 => n22343, B2 => 
                           n20201, ZN => n7339);
   U18017 : OAI22_X1 port map( A1 => n22346, A2 => n22465, B1 => n15193, B2 => 
                           n20202, ZN => n7340);
   U18018 : OAI22_X1 port map( A1 => n22347, A2 => n22471, B1 => n15193, B2 => 
                           n20203, ZN => n7341);
   U18019 : OAI22_X1 port map( A1 => n22347, A2 => n22477, B1 => n15193, B2 => 
                           n20204, ZN => n7342);
   U18020 : OAI22_X1 port map( A1 => n22347, A2 => n22483, B1 => n15193, B2 => 
                           n20205, ZN => n7343);
   U18021 : OAI22_X1 port map( A1 => n22347, A2 => n22489, B1 => n15193, B2 => 
                           n20206, ZN => n7344);
   U18022 : OAI22_X1 port map( A1 => n22347, A2 => n22495, B1 => n15193, B2 => 
                           n20207, ZN => n7345);
   U18023 : OAI22_X1 port map( A1 => n22348, A2 => n22501, B1 => n15193, B2 => 
                           n20208, ZN => n7346);
   U18024 : OAI22_X1 port map( A1 => n22348, A2 => n22507, B1 => n22343, B2 => 
                           n20209, ZN => n7347);
   U18025 : OAI22_X1 port map( A1 => n22348, A2 => n22513, B1 => n22343, B2 => 
                           n20210, ZN => n7348);
   U18026 : OAI22_X1 port map( A1 => n22348, A2 => n22519, B1 => n22343, B2 => 
                           n20211, ZN => n7349);
   U18027 : OAI22_X1 port map( A1 => n22353, A2 => n22386, B1 => n22352, B2 => 
                           n15190, ZN => n7358);
   U18028 : OAI22_X1 port map( A1 => n22353, A2 => n22387, B1 => n22352, B2 => 
                           n15189, ZN => n7359);
   U18029 : OAI22_X1 port map( A1 => n22353, A2 => n22393, B1 => n22352, B2 => 
                           n15188, ZN => n7360);
   U18030 : OAI22_X1 port map( A1 => n22353, A2 => n22399, B1 => n22352, B2 => 
                           n15187, ZN => n7361);
   U18031 : OAI22_X1 port map( A1 => n22353, A2 => n22405, B1 => n22352, B2 => 
                           n15186, ZN => n7362);
   U18032 : OAI22_X1 port map( A1 => n22354, A2 => n22411, B1 => n22352, B2 => 
                           n15185, ZN => n7363);
   U18033 : OAI22_X1 port map( A1 => n22354, A2 => n22417, B1 => n22352, B2 => 
                           n15184, ZN => n7364);
   U18034 : OAI22_X1 port map( A1 => n22354, A2 => n22423, B1 => n22352, B2 => 
                           n15183, ZN => n7365);
   U18035 : OAI22_X1 port map( A1 => n22354, A2 => n22429, B1 => n22352, B2 => 
                           n15182, ZN => n7366);
   U18036 : OAI22_X1 port map( A1 => n22354, A2 => n22435, B1 => n22352, B2 => 
                           n15181, ZN => n7367);
   U18037 : OAI22_X1 port map( A1 => n22355, A2 => n22441, B1 => n22352, B2 => 
                           n15180, ZN => n7368);
   U18038 : OAI22_X1 port map( A1 => n22355, A2 => n22447, B1 => n22352, B2 => 
                           n15179, ZN => n7369);
   U18039 : OAI22_X1 port map( A1 => n22355, A2 => n22453, B1 => n22352, B2 => 
                           n15178, ZN => n7370);
   U18040 : OAI22_X1 port map( A1 => n22355, A2 => n22459, B1 => n22352, B2 => 
                           n15177, ZN => n7371);
   U18041 : OAI22_X1 port map( A1 => n22355, A2 => n22465, B1 => n15158, B2 => 
                           n15176, ZN => n7372);
   U18042 : OAI22_X1 port map( A1 => n22356, A2 => n22471, B1 => n15158, B2 => 
                           n15175, ZN => n7373);
   U18043 : OAI22_X1 port map( A1 => n22356, A2 => n22477, B1 => n15158, B2 => 
                           n15174, ZN => n7374);
   U18044 : OAI22_X1 port map( A1 => n22356, A2 => n22483, B1 => n15158, B2 => 
                           n15173, ZN => n7375);
   U18045 : OAI22_X1 port map( A1 => n22356, A2 => n22489, B1 => n15158, B2 => 
                           n15172, ZN => n7376);
   U18046 : OAI22_X1 port map( A1 => n22356, A2 => n22495, B1 => n15158, B2 => 
                           n15171, ZN => n7377);
   U18047 : OAI22_X1 port map( A1 => n22357, A2 => n22501, B1 => n15158, B2 => 
                           n15170, ZN => n7378);
   U18048 : OAI22_X1 port map( A1 => n22357, A2 => n22507, B1 => n22352, B2 => 
                           n15169, ZN => n7379);
   U18049 : OAI22_X1 port map( A1 => n22357, A2 => n22513, B1 => n22352, B2 => 
                           n15168, ZN => n7380);
   U18050 : OAI22_X1 port map( A1 => n22357, A2 => n22519, B1 => n22352, B2 => 
                           n15167, ZN => n7381);
   U18051 : AOI22_X1 port map( A1 => n21147, A2 => n9533, B1 => n18426, B2 => 
                           n9629, ZN => n19630);
   U18052 : AOI22_X1 port map( A1 => n21704, A2 => n9533, B1 => n16843, B2 => 
                           n9629, ZN => n18357);
   U18053 : OAI22_X1 port map( A1 => n21894, A2 => n22381, B1 => n7456, B2 => 
                           n21893, ZN => n5726);
   U18054 : OAI22_X1 port map( A1 => n21894, A2 => n22391, B1 => n7488, B2 => 
                           n21893, ZN => n5727);
   U18055 : OAI22_X1 port map( A1 => n21894, A2 => n22397, B1 => n7520, B2 => 
                           n21893, ZN => n5728);
   U18056 : OAI22_X1 port map( A1 => n21894, A2 => n22403, B1 => n7552, B2 => 
                           n21893, ZN => n5729);
   U18057 : OAI22_X1 port map( A1 => n21894, A2 => n22409, B1 => n7584, B2 => 
                           n21893, ZN => n5730);
   U18058 : OAI22_X1 port map( A1 => n21895, A2 => n22415, B1 => n7616, B2 => 
                           n21893, ZN => n5731);
   U18059 : OAI22_X1 port map( A1 => n21895, A2 => n22421, B1 => n7648, B2 => 
                           n21893, ZN => n5732);
   U18060 : OAI22_X1 port map( A1 => n21895, A2 => n22427, B1 => n7680, B2 => 
                           n21893, ZN => n5733);
   U18061 : OAI22_X1 port map( A1 => n21895, A2 => n22433, B1 => n7712, B2 => 
                           n21893, ZN => n5734);
   U18062 : OAI22_X1 port map( A1 => n21895, A2 => n22439, B1 => n7744, B2 => 
                           n21893, ZN => n5735);
   U18063 : OAI22_X1 port map( A1 => n21896, A2 => n22445, B1 => n7776, B2 => 
                           n21893, ZN => n5736);
   U18064 : OAI22_X1 port map( A1 => n21896, A2 => n22451, B1 => n7808, B2 => 
                           n21893, ZN => n5737);
   U18065 : OAI22_X1 port map( A1 => n21896, A2 => n22457, B1 => n7840, B2 => 
                           n21893, ZN => n5738);
   U18066 : OAI22_X1 port map( A1 => n21896, A2 => n22463, B1 => n7872, B2 => 
                           n21893, ZN => n5739);
   U18067 : OAI22_X1 port map( A1 => n21896, A2 => n22469, B1 => n7904, B2 => 
                           n16616, ZN => n5740);
   U18068 : OAI22_X1 port map( A1 => n21897, A2 => n22475, B1 => n7936, B2 => 
                           n16616, ZN => n5741);
   U18069 : OAI22_X1 port map( A1 => n21897, A2 => n22481, B1 => n7968, B2 => 
                           n16616, ZN => n5742);
   U18070 : OAI22_X1 port map( A1 => n21897, A2 => n22487, B1 => n8000, B2 => 
                           n16616, ZN => n5743);
   U18071 : OAI22_X1 port map( A1 => n21897, A2 => n22493, B1 => n8032, B2 => 
                           n16616, ZN => n5744);
   U18072 : OAI22_X1 port map( A1 => n21897, A2 => n22499, B1 => n8064, B2 => 
                           n16616, ZN => n5745);
   U18073 : OAI22_X1 port map( A1 => n21898, A2 => n22505, B1 => n8096, B2 => 
                           n16616, ZN => n5746);
   U18074 : OAI22_X1 port map( A1 => n21898, A2 => n22511, B1 => n8128, B2 => 
                           n21893, ZN => n5747);
   U18075 : OAI22_X1 port map( A1 => n21898, A2 => n22517, B1 => n8160, B2 => 
                           n21893, ZN => n5748);
   U18076 : OAI22_X1 port map( A1 => n21898, A2 => n22523, B1 => n8192, B2 => 
                           n21893, ZN => n5749);
   U18077 : OAI22_X1 port map( A1 => n21903, A2 => n22381, B1 => n7457, B2 => 
                           n21902, ZN => n5758);
   U18078 : OAI22_X1 port map( A1 => n21903, A2 => n22391, B1 => n7489, B2 => 
                           n21902, ZN => n5759);
   U18079 : OAI22_X1 port map( A1 => n21903, A2 => n22397, B1 => n7521, B2 => 
                           n21902, ZN => n5760);
   U18080 : OAI22_X1 port map( A1 => n21903, A2 => n22403, B1 => n7553, B2 => 
                           n21902, ZN => n5761);
   U18081 : OAI22_X1 port map( A1 => n21903, A2 => n22409, B1 => n7585, B2 => 
                           n21902, ZN => n5762);
   U18082 : OAI22_X1 port map( A1 => n21904, A2 => n22415, B1 => n7617, B2 => 
                           n21902, ZN => n5763);
   U18083 : OAI22_X1 port map( A1 => n21904, A2 => n22421, B1 => n7649, B2 => 
                           n21902, ZN => n5764);
   U18084 : OAI22_X1 port map( A1 => n21904, A2 => n22427, B1 => n7681, B2 => 
                           n21902, ZN => n5765);
   U18085 : OAI22_X1 port map( A1 => n21904, A2 => n22433, B1 => n7713, B2 => 
                           n21902, ZN => n5766);
   U18086 : OAI22_X1 port map( A1 => n21904, A2 => n22439, B1 => n7745, B2 => 
                           n21902, ZN => n5767);
   U18087 : OAI22_X1 port map( A1 => n21905, A2 => n22445, B1 => n7777, B2 => 
                           n21902, ZN => n5768);
   U18088 : OAI22_X1 port map( A1 => n21905, A2 => n22451, B1 => n7809, B2 => 
                           n21902, ZN => n5769);
   U18089 : OAI22_X1 port map( A1 => n21905, A2 => n22457, B1 => n7841, B2 => 
                           n21902, ZN => n5770);
   U18090 : OAI22_X1 port map( A1 => n21905, A2 => n22463, B1 => n7873, B2 => 
                           n21902, ZN => n5771);
   U18091 : OAI22_X1 port map( A1 => n21905, A2 => n22469, B1 => n7905, B2 => 
                           n16613, ZN => n5772);
   U18092 : OAI22_X1 port map( A1 => n21906, A2 => n22475, B1 => n7937, B2 => 
                           n16613, ZN => n5773);
   U18093 : OAI22_X1 port map( A1 => n21906, A2 => n22481, B1 => n7969, B2 => 
                           n16613, ZN => n5774);
   U18094 : OAI22_X1 port map( A1 => n21906, A2 => n22487, B1 => n8001, B2 => 
                           n16613, ZN => n5775);
   U18095 : OAI22_X1 port map( A1 => n21906, A2 => n22493, B1 => n8033, B2 => 
                           n16613, ZN => n5776);
   U18096 : OAI22_X1 port map( A1 => n21906, A2 => n22499, B1 => n8065, B2 => 
                           n16613, ZN => n5777);
   U18097 : OAI22_X1 port map( A1 => n21907, A2 => n22505, B1 => n8097, B2 => 
                           n16613, ZN => n5778);
   U18098 : OAI22_X1 port map( A1 => n21907, A2 => n22511, B1 => n8129, B2 => 
                           n21902, ZN => n5779);
   U18099 : OAI22_X1 port map( A1 => n21907, A2 => n22517, B1 => n8161, B2 => 
                           n21902, ZN => n5780);
   U18100 : OAI22_X1 port map( A1 => n21907, A2 => n22523, B1 => n8193, B2 => 
                           n21902, ZN => n5781);
   U18101 : OAI22_X1 port map( A1 => n21813, A2 => n22381, B1 => n4350, B2 => 
                           n21812, ZN => n5438);
   U18102 : OAI22_X1 port map( A1 => n21813, A2 => n22392, B1 => n4351, B2 => 
                           n21812, ZN => n5439);
   U18103 : OAI22_X1 port map( A1 => n21813, A2 => n22398, B1 => n4352, B2 => 
                           n21812, ZN => n5440);
   U18104 : OAI22_X1 port map( A1 => n21813, A2 => n22404, B1 => n4353, B2 => 
                           n21812, ZN => n5441);
   U18105 : OAI22_X1 port map( A1 => n21813, A2 => n22410, B1 => n4354, B2 => 
                           n21812, ZN => n5442);
   U18106 : OAI22_X1 port map( A1 => n21814, A2 => n22416, B1 => n4355, B2 => 
                           n21812, ZN => n5443);
   U18107 : OAI22_X1 port map( A1 => n21814, A2 => n22422, B1 => n4356, B2 => 
                           n21812, ZN => n5444);
   U18108 : OAI22_X1 port map( A1 => n21814, A2 => n22428, B1 => n4357, B2 => 
                           n21812, ZN => n5445);
   U18109 : OAI22_X1 port map( A1 => n21814, A2 => n22434, B1 => n4358, B2 => 
                           n21812, ZN => n5446);
   U18110 : OAI22_X1 port map( A1 => n21814, A2 => n22440, B1 => n4359, B2 => 
                           n21812, ZN => n5447);
   U18111 : OAI22_X1 port map( A1 => n21815, A2 => n22446, B1 => n4360, B2 => 
                           n21812, ZN => n5448);
   U18112 : OAI22_X1 port map( A1 => n21815, A2 => n22452, B1 => n4361, B2 => 
                           n21812, ZN => n5449);
   U18113 : OAI22_X1 port map( A1 => n21815, A2 => n22458, B1 => n4362, B2 => 
                           n21812, ZN => n5450);
   U18114 : OAI22_X1 port map( A1 => n21815, A2 => n22464, B1 => n4363, B2 => 
                           n21812, ZN => n5451);
   U18115 : OAI22_X1 port map( A1 => n21815, A2 => n22470, B1 => n4364, B2 => 
                           n16831, ZN => n5452);
   U18116 : OAI22_X1 port map( A1 => n21816, A2 => n22476, B1 => n4365, B2 => 
                           n16831, ZN => n5453);
   U18117 : OAI22_X1 port map( A1 => n21816, A2 => n22482, B1 => n4366, B2 => 
                           n16831, ZN => n5454);
   U18118 : OAI22_X1 port map( A1 => n21816, A2 => n22488, B1 => n4367, B2 => 
                           n16831, ZN => n5455);
   U18119 : OAI22_X1 port map( A1 => n21816, A2 => n22494, B1 => n4368, B2 => 
                           n16831, ZN => n5456);
   U18120 : OAI22_X1 port map( A1 => n21816, A2 => n22500, B1 => n4369, B2 => 
                           n16831, ZN => n5457);
   U18121 : OAI22_X1 port map( A1 => n21817, A2 => n22506, B1 => n4370, B2 => 
                           n16831, ZN => n5458);
   U18122 : OAI22_X1 port map( A1 => n21817, A2 => n22512, B1 => n4371, B2 => 
                           n21812, ZN => n5459);
   U18123 : OAI22_X1 port map( A1 => n21817, A2 => n22518, B1 => n4372, B2 => 
                           n21812, ZN => n5460);
   U18124 : OAI22_X1 port map( A1 => n21817, A2 => n22524, B1 => n4373, B2 => 
                           n21812, ZN => n5461);
   U18125 : OAI22_X1 port map( A1 => n21840, A2 => n22381, B1 => n4382, B2 => 
                           n21839, ZN => n5534);
   U18126 : OAI22_X1 port map( A1 => n21840, A2 => n22391, B1 => n4383, B2 => 
                           n21839, ZN => n5535);
   U18127 : OAI22_X1 port map( A1 => n21840, A2 => n22397, B1 => n4384, B2 => 
                           n21839, ZN => n5536);
   U18128 : OAI22_X1 port map( A1 => n21840, A2 => n22403, B1 => n4385, B2 => 
                           n21839, ZN => n5537);
   U18129 : OAI22_X1 port map( A1 => n21840, A2 => n22409, B1 => n4386, B2 => 
                           n21839, ZN => n5538);
   U18130 : OAI22_X1 port map( A1 => n21841, A2 => n22415, B1 => n4387, B2 => 
                           n21839, ZN => n5539);
   U18131 : OAI22_X1 port map( A1 => n21841, A2 => n22421, B1 => n4388, B2 => 
                           n21839, ZN => n5540);
   U18132 : OAI22_X1 port map( A1 => n21841, A2 => n22427, B1 => n4389, B2 => 
                           n21839, ZN => n5541);
   U18133 : OAI22_X1 port map( A1 => n21841, A2 => n22433, B1 => n4390, B2 => 
                           n21839, ZN => n5542);
   U18134 : OAI22_X1 port map( A1 => n21841, A2 => n22439, B1 => n4391, B2 => 
                           n21839, ZN => n5543);
   U18135 : OAI22_X1 port map( A1 => n21842, A2 => n22445, B1 => n4392, B2 => 
                           n21839, ZN => n5544);
   U18136 : OAI22_X1 port map( A1 => n21842, A2 => n22451, B1 => n4393, B2 => 
                           n21839, ZN => n5545);
   U18137 : OAI22_X1 port map( A1 => n21842, A2 => n22457, B1 => n4394, B2 => 
                           n21839, ZN => n5546);
   U18138 : OAI22_X1 port map( A1 => n21842, A2 => n22463, B1 => n4395, B2 => 
                           n21839, ZN => n5547);
   U18139 : OAI22_X1 port map( A1 => n21842, A2 => n22469, B1 => n4396, B2 => 
                           n16758, ZN => n5548);
   U18140 : OAI22_X1 port map( A1 => n21843, A2 => n22475, B1 => n4397, B2 => 
                           n16758, ZN => n5549);
   U18141 : OAI22_X1 port map( A1 => n21843, A2 => n22481, B1 => n4398, B2 => 
                           n16758, ZN => n5550);
   U18142 : OAI22_X1 port map( A1 => n21843, A2 => n22487, B1 => n4399, B2 => 
                           n16758, ZN => n5551);
   U18143 : OAI22_X1 port map( A1 => n21843, A2 => n22493, B1 => n4400, B2 => 
                           n16758, ZN => n5552);
   U18144 : OAI22_X1 port map( A1 => n21843, A2 => n22499, B1 => n4401, B2 => 
                           n16758, ZN => n5553);
   U18145 : OAI22_X1 port map( A1 => n21844, A2 => n22505, B1 => n4402, B2 => 
                           n16758, ZN => n5554);
   U18146 : OAI22_X1 port map( A1 => n21844, A2 => n22511, B1 => n4403, B2 => 
                           n21839, ZN => n5555);
   U18147 : OAI22_X1 port map( A1 => n21844, A2 => n22517, B1 => n4404, B2 => 
                           n21839, ZN => n5556);
   U18148 : OAI22_X1 port map( A1 => n21844, A2 => n22523, B1 => n4405, B2 => 
                           n21839, ZN => n5557);
   U18149 : OAI22_X1 port map( A1 => n21885, A2 => n22381, B1 => n4478, B2 => 
                           n21884, ZN => n5694);
   U18150 : OAI22_X1 port map( A1 => n21885, A2 => n22391, B1 => n4479, B2 => 
                           n21884, ZN => n5695);
   U18151 : OAI22_X1 port map( A1 => n21885, A2 => n22397, B1 => n4480, B2 => 
                           n21884, ZN => n5696);
   U18152 : OAI22_X1 port map( A1 => n21885, A2 => n22403, B1 => n4481, B2 => 
                           n21884, ZN => n5697);
   U18153 : OAI22_X1 port map( A1 => n21885, A2 => n22409, B1 => n4482, B2 => 
                           n21884, ZN => n5698);
   U18154 : OAI22_X1 port map( A1 => n21886, A2 => n22415, B1 => n4483, B2 => 
                           n21884, ZN => n5699);
   U18155 : OAI22_X1 port map( A1 => n21886, A2 => n22421, B1 => n4484, B2 => 
                           n21884, ZN => n5700);
   U18156 : OAI22_X1 port map( A1 => n21886, A2 => n22427, B1 => n4485, B2 => 
                           n21884, ZN => n5701);
   U18157 : OAI22_X1 port map( A1 => n21886, A2 => n22433, B1 => n4486, B2 => 
                           n21884, ZN => n5702);
   U18158 : OAI22_X1 port map( A1 => n21886, A2 => n22439, B1 => n4487, B2 => 
                           n21884, ZN => n5703);
   U18159 : OAI22_X1 port map( A1 => n21887, A2 => n22445, B1 => n4488, B2 => 
                           n21884, ZN => n5704);
   U18160 : OAI22_X1 port map( A1 => n21887, A2 => n22451, B1 => n4489, B2 => 
                           n21884, ZN => n5705);
   U18161 : OAI22_X1 port map( A1 => n21887, A2 => n22457, B1 => n4490, B2 => 
                           n21884, ZN => n5706);
   U18162 : OAI22_X1 port map( A1 => n21887, A2 => n22463, B1 => n4491, B2 => 
                           n21884, ZN => n5707);
   U18163 : OAI22_X1 port map( A1 => n21887, A2 => n22469, B1 => n4492, B2 => 
                           n16618, ZN => n5708);
   U18164 : OAI22_X1 port map( A1 => n21888, A2 => n22475, B1 => n4493, B2 => 
                           n16618, ZN => n5709);
   U18165 : OAI22_X1 port map( A1 => n21888, A2 => n22481, B1 => n4494, B2 => 
                           n16618, ZN => n5710);
   U18166 : OAI22_X1 port map( A1 => n21888, A2 => n22487, B1 => n4495, B2 => 
                           n16618, ZN => n5711);
   U18167 : OAI22_X1 port map( A1 => n21888, A2 => n22493, B1 => n4496, B2 => 
                           n16618, ZN => n5712);
   U18168 : OAI22_X1 port map( A1 => n21888, A2 => n22499, B1 => n4497, B2 => 
                           n16618, ZN => n5713);
   U18169 : OAI22_X1 port map( A1 => n21889, A2 => n22505, B1 => n4498, B2 => 
                           n16618, ZN => n5714);
   U18170 : OAI22_X1 port map( A1 => n21889, A2 => n22511, B1 => n4499, B2 => 
                           n21884, ZN => n5715);
   U18171 : OAI22_X1 port map( A1 => n21889, A2 => n22517, B1 => n4500, B2 => 
                           n21884, ZN => n5716);
   U18172 : OAI22_X1 port map( A1 => n21889, A2 => n22523, B1 => n4501, B2 => 
                           n21884, ZN => n5717);
   U18173 : OAI22_X1 port map( A1 => n21912, A2 => n22382, B1 => n4510, B2 => 
                           n21911, ZN => n5790);
   U18174 : OAI22_X1 port map( A1 => n21912, A2 => n22391, B1 => n4511, B2 => 
                           n21911, ZN => n5791);
   U18175 : OAI22_X1 port map( A1 => n21912, A2 => n22397, B1 => n4512, B2 => 
                           n21911, ZN => n5792);
   U18176 : OAI22_X1 port map( A1 => n21912, A2 => n22403, B1 => n4513, B2 => 
                           n21911, ZN => n5793);
   U18177 : OAI22_X1 port map( A1 => n21912, A2 => n22409, B1 => n4514, B2 => 
                           n21911, ZN => n5794);
   U18178 : OAI22_X1 port map( A1 => n21913, A2 => n22415, B1 => n4515, B2 => 
                           n21911, ZN => n5795);
   U18179 : OAI22_X1 port map( A1 => n21913, A2 => n22421, B1 => n4516, B2 => 
                           n21911, ZN => n5796);
   U18180 : OAI22_X1 port map( A1 => n21913, A2 => n22427, B1 => n4517, B2 => 
                           n21911, ZN => n5797);
   U18181 : OAI22_X1 port map( A1 => n21913, A2 => n22433, B1 => n4518, B2 => 
                           n21911, ZN => n5798);
   U18182 : OAI22_X1 port map( A1 => n21913, A2 => n22439, B1 => n4519, B2 => 
                           n21911, ZN => n5799);
   U18183 : OAI22_X1 port map( A1 => n21914, A2 => n22445, B1 => n4520, B2 => 
                           n21911, ZN => n5800);
   U18184 : OAI22_X1 port map( A1 => n21914, A2 => n22451, B1 => n4521, B2 => 
                           n21911, ZN => n5801);
   U18185 : OAI22_X1 port map( A1 => n21914, A2 => n22457, B1 => n4522, B2 => 
                           n21911, ZN => n5802);
   U18186 : OAI22_X1 port map( A1 => n21914, A2 => n22463, B1 => n4523, B2 => 
                           n21911, ZN => n5803);
   U18187 : OAI22_X1 port map( A1 => n21914, A2 => n22469, B1 => n4524, B2 => 
                           n16610, ZN => n5804);
   U18188 : OAI22_X1 port map( A1 => n21915, A2 => n22475, B1 => n4525, B2 => 
                           n16610, ZN => n5805);
   U18189 : OAI22_X1 port map( A1 => n21915, A2 => n22481, B1 => n4526, B2 => 
                           n16610, ZN => n5806);
   U18190 : OAI22_X1 port map( A1 => n21915, A2 => n22487, B1 => n4527, B2 => 
                           n16610, ZN => n5807);
   U18191 : OAI22_X1 port map( A1 => n21915, A2 => n22493, B1 => n4528, B2 => 
                           n16610, ZN => n5808);
   U18192 : OAI22_X1 port map( A1 => n21915, A2 => n22499, B1 => n4529, B2 => 
                           n16610, ZN => n5809);
   U18193 : OAI22_X1 port map( A1 => n21916, A2 => n22505, B1 => n4530, B2 => 
                           n16610, ZN => n5810);
   U18194 : OAI22_X1 port map( A1 => n21916, A2 => n22511, B1 => n4531, B2 => 
                           n21911, ZN => n5811);
   U18195 : OAI22_X1 port map( A1 => n21916, A2 => n22517, B1 => n4532, B2 => 
                           n21911, ZN => n5812);
   U18196 : OAI22_X1 port map( A1 => n21916, A2 => n22523, B1 => n4533, B2 => 
                           n21911, ZN => n5813);
   U18197 : OAI22_X1 port map( A1 => n21930, A2 => n22382, B1 => n7454, B2 => 
                           n21929, ZN => n5854);
   U18198 : OAI22_X1 port map( A1 => n21930, A2 => n22391, B1 => n7486, B2 => 
                           n21929, ZN => n5855);
   U18199 : OAI22_X1 port map( A1 => n21930, A2 => n22397, B1 => n7518, B2 => 
                           n16556, ZN => n5856);
   U18200 : OAI22_X1 port map( A1 => n21930, A2 => n22403, B1 => n7550, B2 => 
                           n16556, ZN => n5857);
   U18201 : OAI22_X1 port map( A1 => n21930, A2 => n22409, B1 => n7582, B2 => 
                           n16556, ZN => n5858);
   U18202 : OAI22_X1 port map( A1 => n21931, A2 => n22415, B1 => n7614, B2 => 
                           n21929, ZN => n5859);
   U18203 : OAI22_X1 port map( A1 => n21931, A2 => n22421, B1 => n7646, B2 => 
                           n21929, ZN => n5860);
   U18204 : OAI22_X1 port map( A1 => n21931, A2 => n22427, B1 => n7678, B2 => 
                           n16556, ZN => n5861);
   U18205 : OAI22_X1 port map( A1 => n21931, A2 => n22433, B1 => n7710, B2 => 
                           n16556, ZN => n5862);
   U18206 : OAI22_X1 port map( A1 => n21931, A2 => n22439, B1 => n7742, B2 => 
                           n16556, ZN => n5863);
   U18207 : OAI22_X1 port map( A1 => n21932, A2 => n22445, B1 => n7774, B2 => 
                           n21929, ZN => n5864);
   U18208 : OAI22_X1 port map( A1 => n21932, A2 => n22451, B1 => n7806, B2 => 
                           n16556, ZN => n5865);
   U18209 : OAI22_X1 port map( A1 => n21993, A2 => n22382, B1 => n4670, B2 => 
                           n21992, ZN => n6078);
   U18210 : OAI22_X1 port map( A1 => n21993, A2 => n22390, B1 => n4671, B2 => 
                           n21992, ZN => n6079);
   U18211 : OAI22_X1 port map( A1 => n21993, A2 => n22396, B1 => n4672, B2 => 
                           n21992, ZN => n6080);
   U18212 : OAI22_X1 port map( A1 => n21993, A2 => n22402, B1 => n4673, B2 => 
                           n21992, ZN => n6081);
   U18213 : OAI22_X1 port map( A1 => n21993, A2 => n22408, B1 => n4674, B2 => 
                           n21992, ZN => n6082);
   U18214 : OAI22_X1 port map( A1 => n21994, A2 => n22414, B1 => n4675, B2 => 
                           n21992, ZN => n6083);
   U18215 : OAI22_X1 port map( A1 => n21994, A2 => n22420, B1 => n4676, B2 => 
                           n21992, ZN => n6084);
   U18216 : OAI22_X1 port map( A1 => n21994, A2 => n22426, B1 => n4677, B2 => 
                           n21992, ZN => n6085);
   U18217 : OAI22_X1 port map( A1 => n21994, A2 => n22432, B1 => n4678, B2 => 
                           n21992, ZN => n6086);
   U18218 : OAI22_X1 port map( A1 => n21994, A2 => n22438, B1 => n4679, B2 => 
                           n21992, ZN => n6087);
   U18219 : OAI22_X1 port map( A1 => n21995, A2 => n22444, B1 => n4680, B2 => 
                           n21992, ZN => n6088);
   U18220 : OAI22_X1 port map( A1 => n21995, A2 => n22450, B1 => n4681, B2 => 
                           n21992, ZN => n6089);
   U18221 : OAI22_X1 port map( A1 => n21995, A2 => n22456, B1 => n4682, B2 => 
                           n21992, ZN => n6090);
   U18222 : OAI22_X1 port map( A1 => n21995, A2 => n22462, B1 => n4683, B2 => 
                           n21992, ZN => n6091);
   U18223 : OAI22_X1 port map( A1 => n21995, A2 => n22468, B1 => n4684, B2 => 
                           n16348, ZN => n6092);
   U18224 : OAI22_X1 port map( A1 => n21996, A2 => n22474, B1 => n4685, B2 => 
                           n16348, ZN => n6093);
   U18225 : OAI22_X1 port map( A1 => n21996, A2 => n22480, B1 => n4686, B2 => 
                           n16348, ZN => n6094);
   U18226 : OAI22_X1 port map( A1 => n21996, A2 => n22486, B1 => n4687, B2 => 
                           n16348, ZN => n6095);
   U18227 : OAI22_X1 port map( A1 => n21996, A2 => n22492, B1 => n4688, B2 => 
                           n16348, ZN => n6096);
   U18228 : OAI22_X1 port map( A1 => n21996, A2 => n22498, B1 => n4689, B2 => 
                           n16348, ZN => n6097);
   U18229 : OAI22_X1 port map( A1 => n21997, A2 => n22504, B1 => n4690, B2 => 
                           n16348, ZN => n6098);
   U18230 : OAI22_X1 port map( A1 => n21997, A2 => n22510, B1 => n4691, B2 => 
                           n21992, ZN => n6099);
   U18231 : OAI22_X1 port map( A1 => n21997, A2 => n22516, B1 => n4692, B2 => 
                           n21992, ZN => n6100);
   U18232 : OAI22_X1 port map( A1 => n21997, A2 => n22522, B1 => n4693, B2 => 
                           n21992, ZN => n6101);
   U18233 : OAI22_X1 port map( A1 => n22002, A2 => n22382, B1 => n7466, B2 => 
                           n22001, ZN => n6110);
   U18234 : OAI22_X1 port map( A1 => n22002, A2 => n22390, B1 => n7498, B2 => 
                           n22001, ZN => n6111);
   U18235 : OAI22_X1 port map( A1 => n22002, A2 => n22396, B1 => n7530, B2 => 
                           n22001, ZN => n6112);
   U18236 : OAI22_X1 port map( A1 => n22002, A2 => n22402, B1 => n7562, B2 => 
                           n22001, ZN => n6113);
   U18237 : OAI22_X1 port map( A1 => n22002, A2 => n22408, B1 => n7594, B2 => 
                           n22001, ZN => n6114);
   U18238 : OAI22_X1 port map( A1 => n22003, A2 => n22414, B1 => n7626, B2 => 
                           n22001, ZN => n6115);
   U18239 : OAI22_X1 port map( A1 => n22003, A2 => n22420, B1 => n7658, B2 => 
                           n22001, ZN => n6116);
   U18240 : OAI22_X1 port map( A1 => n22003, A2 => n22426, B1 => n7690, B2 => 
                           n22001, ZN => n6117);
   U18241 : OAI22_X1 port map( A1 => n22003, A2 => n22432, B1 => n7722, B2 => 
                           n22001, ZN => n6118);
   U18242 : OAI22_X1 port map( A1 => n22003, A2 => n22438, B1 => n7754, B2 => 
                           n22001, ZN => n6119);
   U18243 : OAI22_X1 port map( A1 => n22004, A2 => n22444, B1 => n7786, B2 => 
                           n22001, ZN => n6120);
   U18244 : OAI22_X1 port map( A1 => n22004, A2 => n22450, B1 => n7818, B2 => 
                           n22001, ZN => n6121);
   U18245 : OAI22_X1 port map( A1 => n22004, A2 => n22456, B1 => n7850, B2 => 
                           n22001, ZN => n6122);
   U18246 : OAI22_X1 port map( A1 => n22004, A2 => n22462, B1 => n7882, B2 => 
                           n22001, ZN => n6123);
   U18247 : OAI22_X1 port map( A1 => n22004, A2 => n22468, B1 => n7914, B2 => 
                           n16346, ZN => n6124);
   U18248 : OAI22_X1 port map( A1 => n22005, A2 => n22474, B1 => n7946, B2 => 
                           n16346, ZN => n6125);
   U18249 : OAI22_X1 port map( A1 => n22005, A2 => n22480, B1 => n7978, B2 => 
                           n16346, ZN => n6126);
   U18250 : OAI22_X1 port map( A1 => n22005, A2 => n22486, B1 => n8010, B2 => 
                           n16346, ZN => n6127);
   U18251 : OAI22_X1 port map( A1 => n22005, A2 => n22492, B1 => n8042, B2 => 
                           n16346, ZN => n6128);
   U18252 : OAI22_X1 port map( A1 => n22005, A2 => n22498, B1 => n8074, B2 => 
                           n16346, ZN => n6129);
   U18253 : OAI22_X1 port map( A1 => n22006, A2 => n22504, B1 => n8106, B2 => 
                           n16346, ZN => n6130);
   U18254 : OAI22_X1 port map( A1 => n22006, A2 => n22510, B1 => n8138, B2 => 
                           n22001, ZN => n6131);
   U18255 : OAI22_X1 port map( A1 => n22006, A2 => n22516, B1 => n8170, B2 => 
                           n22001, ZN => n6132);
   U18256 : OAI22_X1 port map( A1 => n22006, A2 => n22522, B1 => n8202, B2 => 
                           n22001, ZN => n6133);
   U18257 : OAI22_X1 port map( A1 => n22011, A2 => n22382, B1 => n7467, B2 => 
                           n22010, ZN => n6142);
   U18258 : OAI22_X1 port map( A1 => n22011, A2 => n22390, B1 => n7499, B2 => 
                           n22010, ZN => n6143);
   U18259 : OAI22_X1 port map( A1 => n22011, A2 => n22396, B1 => n7531, B2 => 
                           n22010, ZN => n6144);
   U18260 : OAI22_X1 port map( A1 => n22011, A2 => n22402, B1 => n7563, B2 => 
                           n22010, ZN => n6145);
   U18261 : OAI22_X1 port map( A1 => n22011, A2 => n22408, B1 => n7595, B2 => 
                           n22010, ZN => n6146);
   U18262 : OAI22_X1 port map( A1 => n22012, A2 => n22414, B1 => n7627, B2 => 
                           n22010, ZN => n6147);
   U18263 : OAI22_X1 port map( A1 => n22012, A2 => n22420, B1 => n7659, B2 => 
                           n22010, ZN => n6148);
   U18264 : OAI22_X1 port map( A1 => n22012, A2 => n22426, B1 => n7691, B2 => 
                           n22010, ZN => n6149);
   U18265 : OAI22_X1 port map( A1 => n22012, A2 => n22432, B1 => n7723, B2 => 
                           n22010, ZN => n6150);
   U18266 : OAI22_X1 port map( A1 => n22012, A2 => n22438, B1 => n7755, B2 => 
                           n22010, ZN => n6151);
   U18267 : OAI22_X1 port map( A1 => n22013, A2 => n22444, B1 => n7787, B2 => 
                           n22010, ZN => n6152);
   U18268 : OAI22_X1 port map( A1 => n22013, A2 => n22450, B1 => n7819, B2 => 
                           n22010, ZN => n6153);
   U18269 : OAI22_X1 port map( A1 => n22013, A2 => n22456, B1 => n7851, B2 => 
                           n22010, ZN => n6154);
   U18270 : OAI22_X1 port map( A1 => n22013, A2 => n22462, B1 => n7883, B2 => 
                           n22010, ZN => n6155);
   U18271 : OAI22_X1 port map( A1 => n22013, A2 => n22468, B1 => n7915, B2 => 
                           n16343, ZN => n6156);
   U18272 : OAI22_X1 port map( A1 => n22014, A2 => n22474, B1 => n7947, B2 => 
                           n16343, ZN => n6157);
   U18273 : OAI22_X1 port map( A1 => n22014, A2 => n22480, B1 => n7979, B2 => 
                           n16343, ZN => n6158);
   U18274 : OAI22_X1 port map( A1 => n22014, A2 => n22486, B1 => n8011, B2 => 
                           n16343, ZN => n6159);
   U18275 : OAI22_X1 port map( A1 => n22014, A2 => n22492, B1 => n8043, B2 => 
                           n16343, ZN => n6160);
   U18276 : OAI22_X1 port map( A1 => n22014, A2 => n22498, B1 => n8075, B2 => 
                           n16343, ZN => n6161);
   U18277 : OAI22_X1 port map( A1 => n22015, A2 => n22504, B1 => n8107, B2 => 
                           n16343, ZN => n6162);
   U18278 : OAI22_X1 port map( A1 => n22015, A2 => n22510, B1 => n8139, B2 => 
                           n22010, ZN => n6163);
   U18279 : OAI22_X1 port map( A1 => n22015, A2 => n22516, B1 => n8171, B2 => 
                           n22010, ZN => n6164);
   U18280 : OAI22_X1 port map( A1 => n22015, A2 => n22522, B1 => n8203, B2 => 
                           n22010, ZN => n6165);
   U18281 : OAI22_X1 port map( A1 => n22065, A2 => n22383, B1 => n4798, B2 => 
                           n22064, ZN => n6334);
   U18282 : OAI22_X1 port map( A1 => n22065, A2 => n22389, B1 => n4799, B2 => 
                           n22064, ZN => n6335);
   U18283 : OAI22_X1 port map( A1 => n22065, A2 => n22395, B1 => n4800, B2 => 
                           n22064, ZN => n6336);
   U18284 : OAI22_X1 port map( A1 => n22065, A2 => n22401, B1 => n4801, B2 => 
                           n22064, ZN => n6337);
   U18285 : OAI22_X1 port map( A1 => n22065, A2 => n22407, B1 => n4802, B2 => 
                           n22064, ZN => n6338);
   U18286 : OAI22_X1 port map( A1 => n22066, A2 => n22413, B1 => n4803, B2 => 
                           n22064, ZN => n6339);
   U18287 : OAI22_X1 port map( A1 => n22066, A2 => n22419, B1 => n4804, B2 => 
                           n22064, ZN => n6340);
   U18288 : OAI22_X1 port map( A1 => n22066, A2 => n22425, B1 => n4805, B2 => 
                           n22064, ZN => n6341);
   U18289 : OAI22_X1 port map( A1 => n22066, A2 => n22431, B1 => n4806, B2 => 
                           n22064, ZN => n6342);
   U18290 : OAI22_X1 port map( A1 => n22066, A2 => n22437, B1 => n4807, B2 => 
                           n22064, ZN => n6343);
   U18291 : OAI22_X1 port map( A1 => n22067, A2 => n22443, B1 => n4808, B2 => 
                           n22064, ZN => n6344);
   U18292 : OAI22_X1 port map( A1 => n22067, A2 => n22449, B1 => n4809, B2 => 
                           n22064, ZN => n6345);
   U18293 : OAI22_X1 port map( A1 => n22067, A2 => n22455, B1 => n4810, B2 => 
                           n22064, ZN => n6346);
   U18294 : OAI22_X1 port map( A1 => n22067, A2 => n22461, B1 => n4811, B2 => 
                           n22064, ZN => n6347);
   U18295 : OAI22_X1 port map( A1 => n22067, A2 => n22467, B1 => n4812, B2 => 
                           n16169, ZN => n6348);
   U18296 : OAI22_X1 port map( A1 => n22068, A2 => n22473, B1 => n4813, B2 => 
                           n16169, ZN => n6349);
   U18297 : OAI22_X1 port map( A1 => n22068, A2 => n22479, B1 => n4814, B2 => 
                           n16169, ZN => n6350);
   U18298 : OAI22_X1 port map( A1 => n22068, A2 => n22485, B1 => n4815, B2 => 
                           n16169, ZN => n6351);
   U18299 : OAI22_X1 port map( A1 => n22068, A2 => n22491, B1 => n4816, B2 => 
                           n16169, ZN => n6352);
   U18300 : OAI22_X1 port map( A1 => n22068, A2 => n22497, B1 => n4817, B2 => 
                           n16169, ZN => n6353);
   U18301 : OAI22_X1 port map( A1 => n22069, A2 => n22503, B1 => n4818, B2 => 
                           n16169, ZN => n6354);
   U18302 : OAI22_X1 port map( A1 => n22069, A2 => n22509, B1 => n4819, B2 => 
                           n22064, ZN => n6355);
   U18303 : OAI22_X1 port map( A1 => n22069, A2 => n22515, B1 => n4820, B2 => 
                           n22064, ZN => n6356);
   U18304 : OAI22_X1 port map( A1 => n22069, A2 => n22521, B1 => n4821, B2 => 
                           n22064, ZN => n6357);
   U18305 : OAI22_X1 port map( A1 => n22146, A2 => n22384, B1 => n7474, B2 => 
                           n22145, ZN => n6622);
   U18306 : OAI22_X1 port map( A1 => n22146, A2 => n22389, B1 => n7506, B2 => 
                           n22145, ZN => n6623);
   U18307 : OAI22_X1 port map( A1 => n22146, A2 => n22395, B1 => n7538, B2 => 
                           n22145, ZN => n6624);
   U18308 : OAI22_X1 port map( A1 => n22146, A2 => n22401, B1 => n7570, B2 => 
                           n22145, ZN => n6625);
   U18309 : OAI22_X1 port map( A1 => n22146, A2 => n22407, B1 => n7602, B2 => 
                           n22145, ZN => n6626);
   U18310 : OAI22_X1 port map( A1 => n22147, A2 => n22413, B1 => n7634, B2 => 
                           n22145, ZN => n6627);
   U18311 : OAI22_X1 port map( A1 => n22147, A2 => n22419, B1 => n7666, B2 => 
                           n22145, ZN => n6628);
   U18312 : OAI22_X1 port map( A1 => n22147, A2 => n22425, B1 => n7698, B2 => 
                           n22145, ZN => n6629);
   U18313 : OAI22_X1 port map( A1 => n22147, A2 => n22431, B1 => n7730, B2 => 
                           n22145, ZN => n6630);
   U18314 : OAI22_X1 port map( A1 => n22147, A2 => n22437, B1 => n7762, B2 => 
                           n22145, ZN => n6631);
   U18315 : OAI22_X1 port map( A1 => n22148, A2 => n22443, B1 => n7794, B2 => 
                           n22145, ZN => n6632);
   U18316 : OAI22_X1 port map( A1 => n22148, A2 => n22449, B1 => n7826, B2 => 
                           n22145, ZN => n6633);
   U18317 : OAI22_X1 port map( A1 => n22148, A2 => n22455, B1 => n7858, B2 => 
                           n22145, ZN => n6634);
   U18318 : OAI22_X1 port map( A1 => n22148, A2 => n22461, B1 => n7890, B2 => 
                           n22145, ZN => n6635);
   U18319 : OAI22_X1 port map( A1 => n22148, A2 => n22467, B1 => n7922, B2 => 
                           n15893, ZN => n6636);
   U18320 : OAI22_X1 port map( A1 => n22149, A2 => n22473, B1 => n7954, B2 => 
                           n15893, ZN => n6637);
   U18321 : OAI22_X1 port map( A1 => n22149, A2 => n22479, B1 => n7986, B2 => 
                           n15893, ZN => n6638);
   U18322 : OAI22_X1 port map( A1 => n22149, A2 => n22485, B1 => n8018, B2 => 
                           n15893, ZN => n6639);
   U18323 : OAI22_X1 port map( A1 => n22149, A2 => n22491, B1 => n8050, B2 => 
                           n15893, ZN => n6640);
   U18324 : OAI22_X1 port map( A1 => n22149, A2 => n22497, B1 => n8082, B2 => 
                           n15893, ZN => n6641);
   U18325 : OAI22_X1 port map( A1 => n22150, A2 => n22503, B1 => n8114, B2 => 
                           n15893, ZN => n6642);
   U18326 : OAI22_X1 port map( A1 => n22150, A2 => n22509, B1 => n8146, B2 => 
                           n22145, ZN => n6643);
   U18327 : OAI22_X1 port map( A1 => n22150, A2 => n22515, B1 => n8178, B2 => 
                           n22145, ZN => n6644);
   U18328 : OAI22_X1 port map( A1 => n22150, A2 => n22521, B1 => n8210, B2 => 
                           n22145, ZN => n6645);
   U18329 : OAI22_X1 port map( A1 => n22155, A2 => n22384, B1 => n7475, B2 => 
                           n22154, ZN => n6654);
   U18330 : OAI22_X1 port map( A1 => n22155, A2 => n22389, B1 => n7507, B2 => 
                           n22154, ZN => n6655);
   U18331 : OAI22_X1 port map( A1 => n22155, A2 => n22395, B1 => n7539, B2 => 
                           n22154, ZN => n6656);
   U18332 : OAI22_X1 port map( A1 => n22155, A2 => n22401, B1 => n7571, B2 => 
                           n22154, ZN => n6657);
   U18333 : OAI22_X1 port map( A1 => n22155, A2 => n22407, B1 => n7603, B2 => 
                           n22154, ZN => n6658);
   U18334 : OAI22_X1 port map( A1 => n22156, A2 => n22413, B1 => n7635, B2 => 
                           n22154, ZN => n6659);
   U18335 : OAI22_X1 port map( A1 => n22156, A2 => n22419, B1 => n7667, B2 => 
                           n22154, ZN => n6660);
   U18336 : OAI22_X1 port map( A1 => n22156, A2 => n22425, B1 => n7699, B2 => 
                           n22154, ZN => n6661);
   U18337 : OAI22_X1 port map( A1 => n22156, A2 => n22431, B1 => n7731, B2 => 
                           n22154, ZN => n6662);
   U18338 : OAI22_X1 port map( A1 => n22156, A2 => n22437, B1 => n7763, B2 => 
                           n22154, ZN => n6663);
   U18339 : OAI22_X1 port map( A1 => n22157, A2 => n22443, B1 => n7795, B2 => 
                           n22154, ZN => n6664);
   U18340 : OAI22_X1 port map( A1 => n22157, A2 => n22449, B1 => n7827, B2 => 
                           n22154, ZN => n6665);
   U18341 : OAI22_X1 port map( A1 => n22157, A2 => n22455, B1 => n7859, B2 => 
                           n22154, ZN => n6666);
   U18342 : OAI22_X1 port map( A1 => n22157, A2 => n22461, B1 => n7891, B2 => 
                           n22154, ZN => n6667);
   U18343 : OAI22_X1 port map( A1 => n22157, A2 => n22467, B1 => n7923, B2 => 
                           n15890, ZN => n6668);
   U18344 : OAI22_X1 port map( A1 => n22158, A2 => n22473, B1 => n7955, B2 => 
                           n15890, ZN => n6669);
   U18345 : OAI22_X1 port map( A1 => n22158, A2 => n22479, B1 => n7987, B2 => 
                           n15890, ZN => n6670);
   U18346 : OAI22_X1 port map( A1 => n22158, A2 => n22485, B1 => n8019, B2 => 
                           n15890, ZN => n6671);
   U18347 : OAI22_X1 port map( A1 => n22158, A2 => n22491, B1 => n8051, B2 => 
                           n15890, ZN => n6672);
   U18348 : OAI22_X1 port map( A1 => n22158, A2 => n22497, B1 => n8083, B2 => 
                           n15890, ZN => n6673);
   U18349 : OAI22_X1 port map( A1 => n22159, A2 => n22503, B1 => n8115, B2 => 
                           n15890, ZN => n6674);
   U18350 : OAI22_X1 port map( A1 => n22159, A2 => n22509, B1 => n8147, B2 => 
                           n22154, ZN => n6675);
   U18351 : OAI22_X1 port map( A1 => n22159, A2 => n22515, B1 => n8179, B2 => 
                           n22154, ZN => n6676);
   U18352 : OAI22_X1 port map( A1 => n22159, A2 => n22521, B1 => n8211, B2 => 
                           n22154, ZN => n6677);
   U18353 : OAI22_X1 port map( A1 => n22200, A2 => n22384, B1 => n5022, B2 => 
                           n22199, ZN => n6814);
   U18354 : OAI22_X1 port map( A1 => n22200, A2 => n22388, B1 => n5023, B2 => 
                           n22199, ZN => n6815);
   U18355 : OAI22_X1 port map( A1 => n22200, A2 => n22394, B1 => n5024, B2 => 
                           n22199, ZN => n6816);
   U18356 : OAI22_X1 port map( A1 => n22200, A2 => n22400, B1 => n5025, B2 => 
                           n22199, ZN => n6817);
   U18357 : OAI22_X1 port map( A1 => n22200, A2 => n22406, B1 => n5026, B2 => 
                           n22199, ZN => n6818);
   U18358 : OAI22_X1 port map( A1 => n22201, A2 => n22412, B1 => n5027, B2 => 
                           n22199, ZN => n6819);
   U18359 : OAI22_X1 port map( A1 => n22201, A2 => n22418, B1 => n5028, B2 => 
                           n22199, ZN => n6820);
   U18360 : OAI22_X1 port map( A1 => n22201, A2 => n22424, B1 => n5029, B2 => 
                           n22199, ZN => n6821);
   U18361 : OAI22_X1 port map( A1 => n22201, A2 => n22430, B1 => n5030, B2 => 
                           n22199, ZN => n6822);
   U18362 : OAI22_X1 port map( A1 => n22201, A2 => n22436, B1 => n5031, B2 => 
                           n22199, ZN => n6823);
   U18363 : OAI22_X1 port map( A1 => n22202, A2 => n22442, B1 => n5032, B2 => 
                           n22199, ZN => n6824);
   U18364 : OAI22_X1 port map( A1 => n22202, A2 => n22448, B1 => n5033, B2 => 
                           n22199, ZN => n6825);
   U18365 : OAI22_X1 port map( A1 => n22202, A2 => n22454, B1 => n5034, B2 => 
                           n22199, ZN => n6826);
   U18366 : OAI22_X1 port map( A1 => n22202, A2 => n22460, B1 => n5035, B2 => 
                           n22199, ZN => n6827);
   U18367 : OAI22_X1 port map( A1 => n22202, A2 => n22466, B1 => n5036, B2 => 
                           n15750, ZN => n6828);
   U18368 : OAI22_X1 port map( A1 => n22203, A2 => n22472, B1 => n5037, B2 => 
                           n15750, ZN => n6829);
   U18369 : OAI22_X1 port map( A1 => n22203, A2 => n22478, B1 => n5038, B2 => 
                           n15750, ZN => n6830);
   U18370 : OAI22_X1 port map( A1 => n22203, A2 => n22484, B1 => n5039, B2 => 
                           n15750, ZN => n6831);
   U18371 : OAI22_X1 port map( A1 => n22203, A2 => n22490, B1 => n5040, B2 => 
                           n15750, ZN => n6832);
   U18372 : OAI22_X1 port map( A1 => n22203, A2 => n22496, B1 => n5041, B2 => 
                           n15750, ZN => n6833);
   U18373 : OAI22_X1 port map( A1 => n22204, A2 => n22502, B1 => n5042, B2 => 
                           n15750, ZN => n6834);
   U18374 : OAI22_X1 port map( A1 => n22204, A2 => n22508, B1 => n5043, B2 => 
                           n22199, ZN => n6835);
   U18375 : OAI22_X1 port map( A1 => n22204, A2 => n22514, B1 => n5044, B2 => 
                           n22199, ZN => n6836);
   U18376 : OAI22_X1 port map( A1 => n22204, A2 => n22520, B1 => n5045, B2 => 
                           n22199, ZN => n6837);
   U18377 : OAI22_X1 port map( A1 => n22362, A2 => n22386, B1 => n7478, B2 => 
                           n22361, ZN => n7390);
   U18378 : OAI22_X1 port map( A1 => n22362, A2 => n22387, B1 => n7510, B2 => 
                           n22361, ZN => n7391);
   U18379 : OAI22_X1 port map( A1 => n22362, A2 => n22393, B1 => n7542, B2 => 
                           n22361, ZN => n7392);
   U18380 : OAI22_X1 port map( A1 => n22362, A2 => n22399, B1 => n7574, B2 => 
                           n22361, ZN => n7393);
   U18381 : OAI22_X1 port map( A1 => n22362, A2 => n22405, B1 => n7606, B2 => 
                           n22361, ZN => n7394);
   U18382 : OAI22_X1 port map( A1 => n22363, A2 => n22411, B1 => n7638, B2 => 
                           n22361, ZN => n7395);
   U18383 : OAI22_X1 port map( A1 => n22363, A2 => n22417, B1 => n7670, B2 => 
                           n22361, ZN => n7396);
   U18384 : OAI22_X1 port map( A1 => n22363, A2 => n22423, B1 => n7702, B2 => 
                           n22361, ZN => n7397);
   U18385 : OAI22_X1 port map( A1 => n22363, A2 => n22429, B1 => n7734, B2 => 
                           n22361, ZN => n7398);
   U18386 : OAI22_X1 port map( A1 => n22363, A2 => n22435, B1 => n7766, B2 => 
                           n22361, ZN => n7399);
   U18387 : OAI22_X1 port map( A1 => n22364, A2 => n22441, B1 => n7798, B2 => 
                           n22361, ZN => n7400);
   U18388 : OAI22_X1 port map( A1 => n22364, A2 => n22447, B1 => n7830, B2 => 
                           n22361, ZN => n7401);
   U18389 : OAI22_X1 port map( A1 => n22364, A2 => n22453, B1 => n7862, B2 => 
                           n22361, ZN => n7402);
   U18390 : OAI22_X1 port map( A1 => n22364, A2 => n22459, B1 => n7894, B2 => 
                           n22361, ZN => n7403);
   U18391 : OAI22_X1 port map( A1 => n22364, A2 => n22465, B1 => n7926, B2 => 
                           n15155, ZN => n7404);
   U18392 : OAI22_X1 port map( A1 => n22365, A2 => n22471, B1 => n7958, B2 => 
                           n15155, ZN => n7405);
   U18393 : OAI22_X1 port map( A1 => n22365, A2 => n22477, B1 => n7990, B2 => 
                           n15155, ZN => n7406);
   U18394 : OAI22_X1 port map( A1 => n22365, A2 => n22483, B1 => n8022, B2 => 
                           n15155, ZN => n7407);
   U18395 : OAI22_X1 port map( A1 => n22365, A2 => n22489, B1 => n8054, B2 => 
                           n15155, ZN => n7408);
   U18396 : OAI22_X1 port map( A1 => n22365, A2 => n22495, B1 => n8086, B2 => 
                           n15155, ZN => n7409);
   U18397 : OAI22_X1 port map( A1 => n22366, A2 => n22501, B1 => n8118, B2 => 
                           n15155, ZN => n7410);
   U18398 : OAI22_X1 port map( A1 => n22366, A2 => n22507, B1 => n8150, B2 => 
                           n22361, ZN => n7411);
   U18399 : OAI22_X1 port map( A1 => n22366, A2 => n22513, B1 => n8182, B2 => 
                           n22361, ZN => n7412);
   U18400 : OAI22_X1 port map( A1 => n22366, A2 => n22519, B1 => n8214, B2 => 
                           n22361, ZN => n7413);
   U18401 : OAI22_X1 port map( A1 => n22568, A2 => n22386, B1 => n7479, B2 => 
                           n22567, ZN => n7422);
   U18402 : OAI22_X1 port map( A1 => n22568, A2 => n22387, B1 => n7511, B2 => 
                           n22567, ZN => n7423);
   U18403 : OAI22_X1 port map( A1 => n22568, A2 => n22393, B1 => n7543, B2 => 
                           n22567, ZN => n7424);
   U18404 : OAI22_X1 port map( A1 => n22568, A2 => n22399, B1 => n7575, B2 => 
                           n22567, ZN => n7425);
   U18405 : OAI22_X1 port map( A1 => n22568, A2 => n22405, B1 => n7607, B2 => 
                           n22567, ZN => n7426);
   U18406 : OAI22_X1 port map( A1 => n22569, A2 => n22411, B1 => n7639, B2 => 
                           n22567, ZN => n7427);
   U18407 : OAI22_X1 port map( A1 => n22569, A2 => n22417, B1 => n7671, B2 => 
                           n22567, ZN => n7428);
   U18408 : OAI22_X1 port map( A1 => n22569, A2 => n22423, B1 => n7703, B2 => 
                           n22567, ZN => n7429);
   U18409 : OAI22_X1 port map( A1 => n22569, A2 => n22429, B1 => n7735, B2 => 
                           n22567, ZN => n7430);
   U18410 : OAI22_X1 port map( A1 => n22569, A2 => n22435, B1 => n7767, B2 => 
                           n22567, ZN => n7431);
   U18411 : OAI22_X1 port map( A1 => n22570, A2 => n22441, B1 => n7799, B2 => 
                           n22567, ZN => n7432);
   U18412 : OAI22_X1 port map( A1 => n22570, A2 => n22447, B1 => n7831, B2 => 
                           n22567, ZN => n7433);
   U18413 : OAI22_X1 port map( A1 => n22570, A2 => n22453, B1 => n7863, B2 => 
                           n22567, ZN => n7434);
   U18414 : OAI22_X1 port map( A1 => n22570, A2 => n22459, B1 => n7895, B2 => 
                           n22567, ZN => n7435);
   U18415 : OAI22_X1 port map( A1 => n22570, A2 => n22465, B1 => n7927, B2 => 
                           n15119, ZN => n7436);
   U18416 : OAI22_X1 port map( A1 => n22571, A2 => n22471, B1 => n7959, B2 => 
                           n15119, ZN => n7437);
   U18417 : OAI22_X1 port map( A1 => n22571, A2 => n22477, B1 => n7991, B2 => 
                           n15119, ZN => n7438);
   U18418 : OAI22_X1 port map( A1 => n22571, A2 => n22483, B1 => n8023, B2 => 
                           n15119, ZN => n7439);
   U18419 : OAI22_X1 port map( A1 => n22571, A2 => n22489, B1 => n8055, B2 => 
                           n15119, ZN => n7440);
   U18420 : OAI22_X1 port map( A1 => n22571, A2 => n22495, B1 => n8087, B2 => 
                           n15119, ZN => n7441);
   U18421 : OAI22_X1 port map( A1 => n22572, A2 => n22501, B1 => n8119, B2 => 
                           n15119, ZN => n7442);
   U18422 : OAI22_X1 port map( A1 => n22572, A2 => n22507, B1 => n8151, B2 => 
                           n22567, ZN => n7443);
   U18423 : OAI22_X1 port map( A1 => n22572, A2 => n22513, B1 => n8183, B2 => 
                           n22567, ZN => n7444);
   U18424 : OAI22_X1 port map( A1 => n22572, A2 => n22519, B1 => n8215, B2 => 
                           n22567, ZN => n7445);
   U18425 : OAI22_X1 port map( A1 => n21932, A2 => n22457, B1 => n7838, B2 => 
                           n21929, ZN => n5866);
   U18426 : OAI22_X1 port map( A1 => n21932, A2 => n22463, B1 => n7870, B2 => 
                           n21929, ZN => n5867);
   U18427 : AOI22_X1 port map( A1 => n21114, A2 => n9469, B1 => n18432, B2 => 
                           n19999, ZN => n19628);
   U18428 : AOI22_X1 port map( A1 => n21671, A2 => n9469, B1 => n16849, B2 => 
                           n19999, ZN => n18355);
   U18429 : NAND4_X1 port map( A1 => n19638, A2 => n19639, A3 => n19640, A4 => 
                           n19641, ZN => n19617);
   U18430 : AOI221_X1 port map( B1 => n18500, B2 => n8957, C1 => n18501, C2 => 
                           n8509, A => n19679, ZN => n19638);
   U18431 : AOI221_X1 port map( B1 => n18495, B2 => n8917, C1 => n20840, C2 => 
                           n19811, A => n19676, ZN => n19639);
   U18432 : AOI221_X1 port map( B1 => n18490, B2 => n8916, C1 => n18491, C2 => 
                           n19812, A => n19672, ZN => n19640);
   U18433 : NAND4_X1 port map( A1 => n18366, A2 => n18367, A3 => n18368, A4 => 
                           n18369, ZN => n18344);
   U18434 : AOI221_X1 port map( B1 => n16927, B2 => n8957, C1 => n16928, C2 => 
                           n8509, A => n18416, ZN => n18366);
   U18435 : AOI221_X1 port map( B1 => n16921, B2 => n8917, C1 => n21397, C2 => 
                           n19811, A => n18413, ZN => n18367);
   U18436 : AOI221_X1 port map( B1 => n16915, B2 => n8916, C1 => n16916, C2 => 
                           n19812, A => n18408, ZN => n18368);
   U18437 : AND3_X1 port map( A1 => n15645, A2 => n15643, A3 => ADD_WR(5), ZN 
                           => n16204);
   U18438 : AND3_X1 port map( A1 => n15645, A2 => n15644, A3 => ADD_WR(4), ZN 
                           => n15751);
   U18439 : AND3_X1 port map( A1 => ADD_WR(4), A2 => n15645, A3 => ADD_WR(5), 
                           ZN => n16611);
   U18440 : AND2_X1 port map( A1 => ADD_WR(3), A2 => n16653, ZN => n15504);
   U18441 : AND2_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(2), ZN => n15642);
   U18442 : INV_X1 port map( A => ADD_RD1(4), ZN => n19666);
   U18443 : INV_X1 port map( A => ADD_RD2(4), ZN => n18400);
   U18444 : INV_X1 port map( A => ADD_RD1(0), ZN => n19646);
   U18445 : INV_X1 port map( A => ADD_RD2(0), ZN => n18375);
   U18446 : INV_X1 port map( A => ADD_RD1(3), ZN => n19665);
   U18447 : INV_X1 port map( A => ADD_RD2(3), ZN => n18399);
   U18448 : INV_X1 port map( A => ADD_RD1(5), ZN => n19671);
   U18449 : INV_X1 port map( A => ADD_RD2(5), ZN => n18406);
   U18450 : OAI21_X1 port map( B1 => n4255, B2 => n18417, A => n19578, ZN => 
                           n5343);
   U18451 : OAI21_X1 port map( B1 => n19579, B2 => n19580, A => n18417, ZN => 
                           n19578);
   U18452 : NAND4_X1 port map( A1 => n19581, A2 => n19582, A3 => n19583, A4 => 
                           n19584, ZN => n19580);
   U18453 : NAND4_X1 port map( A1 => n19589, A2 => n19590, A3 => n19591, A4 => 
                           n19592, ZN => n19579);
   U18454 : OAI21_X1 port map( B1 => n4256, B2 => n18417, A => n19541, ZN => 
                           n5344);
   U18455 : OAI21_X1 port map( B1 => n19542, B2 => n19543, A => n18417, ZN => 
                           n19541);
   U18456 : NAND4_X1 port map( A1 => n19544, A2 => n19545, A3 => n19546, A4 => 
                           n19547, ZN => n19543);
   U18457 : NAND4_X1 port map( A1 => n19552, A2 => n19553, A3 => n19554, A4 => 
                           n19555, ZN => n19542);
   U18458 : OAI21_X1 port map( B1 => n4257, B2 => n18417, A => n19504, ZN => 
                           n5345);
   U18459 : OAI21_X1 port map( B1 => n19505, B2 => n19506, A => n18417, ZN => 
                           n19504);
   U18460 : NAND4_X1 port map( A1 => n19507, A2 => n19508, A3 => n19509, A4 => 
                           n19510, ZN => n19506);
   U18461 : NAND4_X1 port map( A1 => n19515, A2 => n19516, A3 => n19517, A4 => 
                           n19518, ZN => n19505);
   U18462 : OAI21_X1 port map( B1 => n4258, B2 => n18417, A => n19467, ZN => 
                           n5346);
   U18463 : OAI21_X1 port map( B1 => n19468, B2 => n19469, A => n18417, ZN => 
                           n19467);
   U18464 : NAND4_X1 port map( A1 => n19470, A2 => n19471, A3 => n19472, A4 => 
                           n19473, ZN => n19469);
   U18465 : NAND4_X1 port map( A1 => n19478, A2 => n19479, A3 => n19480, A4 => 
                           n19481, ZN => n19468);
   U18466 : OAI21_X1 port map( B1 => n4259, B2 => n18417, A => n19430, ZN => 
                           n5347);
   U18467 : OAI21_X1 port map( B1 => n19431, B2 => n19432, A => n18417, ZN => 
                           n19430);
   U18468 : NAND4_X1 port map( A1 => n19433, A2 => n19434, A3 => n19435, A4 => 
                           n19436, ZN => n19432);
   U18469 : NAND4_X1 port map( A1 => n19441, A2 => n19442, A3 => n19443, A4 => 
                           n19444, ZN => n19431);
   U18470 : OAI21_X1 port map( B1 => n4260, B2 => n18417, A => n19393, ZN => 
                           n5348);
   U18471 : OAI21_X1 port map( B1 => n19394, B2 => n19395, A => n18417, ZN => 
                           n19393);
   U18472 : NAND4_X1 port map( A1 => n19396, A2 => n19397, A3 => n19398, A4 => 
                           n19399, ZN => n19395);
   U18473 : NAND4_X1 port map( A1 => n19404, A2 => n19405, A3 => n19406, A4 => 
                           n19407, ZN => n19394);
   U18474 : OAI21_X1 port map( B1 => n4261, B2 => n18417, A => n19356, ZN => 
                           n5349);
   U18475 : OAI21_X1 port map( B1 => n19357, B2 => n19358, A => n18417, ZN => 
                           n19356);
   U18476 : NAND4_X1 port map( A1 => n19359, A2 => n19360, A3 => n19361, A4 => 
                           n19362, ZN => n19358);
   U18477 : NAND4_X1 port map( A1 => n19367, A2 => n19368, A3 => n19369, A4 => 
                           n19370, ZN => n19357);
   U18478 : OAI21_X1 port map( B1 => n4262, B2 => n18417, A => n19319, ZN => 
                           n5350);
   U18479 : OAI21_X1 port map( B1 => n19320, B2 => n19321, A => n18417, ZN => 
                           n19319);
   U18480 : NAND4_X1 port map( A1 => n19322, A2 => n19323, A3 => n19324, A4 => 
                           n19325, ZN => n19321);
   U18481 : NAND4_X1 port map( A1 => n19330, A2 => n19331, A3 => n19332, A4 => 
                           n19333, ZN => n19320);
   U18482 : OAI21_X1 port map( B1 => n4263, B2 => n18417, A => n19282, ZN => 
                           n5351);
   U18483 : OAI21_X1 port map( B1 => n19283, B2 => n19284, A => n18417, ZN => 
                           n19282);
   U18484 : NAND4_X1 port map( A1 => n19285, A2 => n19286, A3 => n19287, A4 => 
                           n19288, ZN => n19284);
   U18485 : NAND4_X1 port map( A1 => n19293, A2 => n19294, A3 => n19295, A4 => 
                           n19296, ZN => n19283);
   U18486 : OAI21_X1 port map( B1 => n4264, B2 => n18417, A => n19245, ZN => 
                           n5352);
   U18487 : OAI21_X1 port map( B1 => n19246, B2 => n19247, A => n18417, ZN => 
                           n19245);
   U18488 : NAND4_X1 port map( A1 => n19248, A2 => n19249, A3 => n19250, A4 => 
                           n19251, ZN => n19247);
   U18489 : NAND4_X1 port map( A1 => n19256, A2 => n19257, A3 => n19258, A4 => 
                           n19259, ZN => n19246);
   U18490 : OAI21_X1 port map( B1 => n4265, B2 => n18417, A => n19208, ZN => 
                           n5353);
   U18491 : OAI21_X1 port map( B1 => n19209, B2 => n19210, A => n18417, ZN => 
                           n19208);
   U18492 : NAND4_X1 port map( A1 => n19211, A2 => n19212, A3 => n19213, A4 => 
                           n19214, ZN => n19210);
   U18493 : NAND4_X1 port map( A1 => n19219, A2 => n19220, A3 => n19221, A4 => 
                           n19222, ZN => n19209);
   U18494 : OAI21_X1 port map( B1 => n4266, B2 => n18417, A => n19171, ZN => 
                           n5354);
   U18495 : OAI21_X1 port map( B1 => n19172, B2 => n19173, A => n18417, ZN => 
                           n19171);
   U18496 : NAND4_X1 port map( A1 => n19174, A2 => n19175, A3 => n19176, A4 => 
                           n19177, ZN => n19173);
   U18497 : NAND4_X1 port map( A1 => n19182, A2 => n19183, A3 => n19184, A4 => 
                           n19185, ZN => n19172);
   U18498 : OAI21_X1 port map( B1 => n4267, B2 => n18417, A => n19134, ZN => 
                           n5355);
   U18499 : OAI21_X1 port map( B1 => n19135, B2 => n19136, A => n18417, ZN => 
                           n19134);
   U18500 : NAND4_X1 port map( A1 => n19137, A2 => n19138, A3 => n19139, A4 => 
                           n19140, ZN => n19136);
   U18501 : NAND4_X1 port map( A1 => n19145, A2 => n19146, A3 => n19147, A4 => 
                           n19148, ZN => n19135);
   U18502 : OAI21_X1 port map( B1 => n4268, B2 => n18417, A => n19097, ZN => 
                           n5356);
   U18503 : OAI21_X1 port map( B1 => n19098, B2 => n19099, A => n18417, ZN => 
                           n19097);
   U18504 : NAND4_X1 port map( A1 => n19100, A2 => n19101, A3 => n19102, A4 => 
                           n19103, ZN => n19099);
   U18505 : NAND4_X1 port map( A1 => n19108, A2 => n19109, A3 => n19110, A4 => 
                           n19111, ZN => n19098);
   U18506 : OAI21_X1 port map( B1 => n4269, B2 => n18417, A => n19060, ZN => 
                           n5357);
   U18507 : OAI21_X1 port map( B1 => n19061, B2 => n19062, A => n18417, ZN => 
                           n19060);
   U18508 : NAND4_X1 port map( A1 => n19063, A2 => n19064, A3 => n19065, A4 => 
                           n19066, ZN => n19062);
   U18509 : NAND4_X1 port map( A1 => n19071, A2 => n19072, A3 => n19073, A4 => 
                           n19074, ZN => n19061);
   U18510 : OAI21_X1 port map( B1 => n4270, B2 => n18417, A => n19023, ZN => 
                           n5358);
   U18511 : OAI21_X1 port map( B1 => n19024, B2 => n19025, A => n18417, ZN => 
                           n19023);
   U18512 : NAND4_X1 port map( A1 => n19026, A2 => n19027, A3 => n19028, A4 => 
                           n19029, ZN => n19025);
   U18513 : NAND4_X1 port map( A1 => n19034, A2 => n19035, A3 => n19036, A4 => 
                           n19037, ZN => n19024);
   U18514 : OAI21_X1 port map( B1 => n4271, B2 => n18417, A => n18986, ZN => 
                           n5359);
   U18515 : OAI21_X1 port map( B1 => n18987, B2 => n18988, A => n18417, ZN => 
                           n18986);
   U18516 : NAND4_X1 port map( A1 => n18989, A2 => n18990, A3 => n18991, A4 => 
                           n18992, ZN => n18988);
   U18517 : NAND4_X1 port map( A1 => n18997, A2 => n18998, A3 => n18999, A4 => 
                           n19000, ZN => n18987);
   U18518 : OAI21_X1 port map( B1 => n4272, B2 => n18417, A => n18949, ZN => 
                           n5360);
   U18519 : OAI21_X1 port map( B1 => n18950, B2 => n18951, A => n18417, ZN => 
                           n18949);
   U18520 : NAND4_X1 port map( A1 => n18952, A2 => n18953, A3 => n18954, A4 => 
                           n18955, ZN => n18951);
   U18521 : NAND4_X1 port map( A1 => n18960, A2 => n18961, A3 => n18962, A4 => 
                           n18963, ZN => n18950);
   U18522 : OAI21_X1 port map( B1 => n4273, B2 => n18417, A => n18912, ZN => 
                           n5361);
   U18523 : OAI21_X1 port map( B1 => n18913, B2 => n18914, A => n18417, ZN => 
                           n18912);
   U18524 : NAND4_X1 port map( A1 => n18915, A2 => n18916, A3 => n18917, A4 => 
                           n18918, ZN => n18914);
   U18525 : NAND4_X1 port map( A1 => n18923, A2 => n18924, A3 => n18925, A4 => 
                           n18926, ZN => n18913);
   U18526 : OAI21_X1 port map( B1 => n4274, B2 => n18417, A => n18875, ZN => 
                           n5362);
   U18527 : OAI21_X1 port map( B1 => n18876, B2 => n18877, A => n18417, ZN => 
                           n18875);
   U18528 : NAND4_X1 port map( A1 => n18878, A2 => n18879, A3 => n18880, A4 => 
                           n18881, ZN => n18877);
   U18529 : NAND4_X1 port map( A1 => n18886, A2 => n18887, A3 => n18888, A4 => 
                           n18889, ZN => n18876);
   U18530 : OAI21_X1 port map( B1 => n4275, B2 => n18417, A => n18838, ZN => 
                           n5363);
   U18531 : OAI21_X1 port map( B1 => n18839, B2 => n18840, A => n18417, ZN => 
                           n18838);
   U18532 : NAND4_X1 port map( A1 => n18841, A2 => n18842, A3 => n18843, A4 => 
                           n18844, ZN => n18840);
   U18533 : NAND4_X1 port map( A1 => n18849, A2 => n18850, A3 => n18851, A4 => 
                           n18852, ZN => n18839);
   U18534 : OAI21_X1 port map( B1 => n4276, B2 => n18417, A => n18801, ZN => 
                           n5364);
   U18535 : OAI21_X1 port map( B1 => n18802, B2 => n18803, A => n18417, ZN => 
                           n18801);
   U18536 : NAND4_X1 port map( A1 => n18804, A2 => n18805, A3 => n18806, A4 => 
                           n18807, ZN => n18803);
   U18537 : NAND4_X1 port map( A1 => n18812, A2 => n18813, A3 => n18814, A4 => 
                           n18815, ZN => n18802);
   U18538 : OAI21_X1 port map( B1 => n4277, B2 => n18417, A => n18764, ZN => 
                           n5365);
   U18539 : OAI21_X1 port map( B1 => n18765, B2 => n18766, A => n18417, ZN => 
                           n18764);
   U18540 : NAND4_X1 port map( A1 => n18767, A2 => n18768, A3 => n18769, A4 => 
                           n18770, ZN => n18766);
   U18541 : NAND4_X1 port map( A1 => n18775, A2 => n18776, A3 => n18777, A4 => 
                           n18778, ZN => n18765);
   U18542 : OAI21_X1 port map( B1 => n4278, B2 => n18417, A => n18727, ZN => 
                           n5366);
   U18543 : OAI21_X1 port map( B1 => n18728, B2 => n18729, A => n18417, ZN => 
                           n18727);
   U18544 : NAND4_X1 port map( A1 => n18730, A2 => n18731, A3 => n18732, A4 => 
                           n18733, ZN => n18729);
   U18545 : NAND4_X1 port map( A1 => n18738, A2 => n18739, A3 => n18740, A4 => 
                           n18741, ZN => n18728);
   U18546 : OAI21_X1 port map( B1 => n4279, B2 => n18417, A => n18690, ZN => 
                           n5367);
   U18547 : OAI21_X1 port map( B1 => n18691, B2 => n18692, A => n18417, ZN => 
                           n18690);
   U18548 : NAND4_X1 port map( A1 => n18693, A2 => n18694, A3 => n18695, A4 => 
                           n18696, ZN => n18692);
   U18549 : NAND4_X1 port map( A1 => n18701, A2 => n18702, A3 => n18703, A4 => 
                           n18704, ZN => n18691);
   U18550 : OAI21_X1 port map( B1 => n4280, B2 => n18417, A => n18653, ZN => 
                           n5368);
   U18551 : OAI21_X1 port map( B1 => n18654, B2 => n18655, A => n18417, ZN => 
                           n18653);
   U18552 : NAND4_X1 port map( A1 => n18656, A2 => n18657, A3 => n18658, A4 => 
                           n18659, ZN => n18655);
   U18553 : NAND4_X1 port map( A1 => n18664, A2 => n18665, A3 => n18666, A4 => 
                           n18667, ZN => n18654);
   U18554 : OAI21_X1 port map( B1 => n4281, B2 => n18417, A => n18616, ZN => 
                           n5369);
   U18555 : OAI21_X1 port map( B1 => n18617, B2 => n18618, A => n18417, ZN => 
                           n18616);
   U18556 : NAND4_X1 port map( A1 => n18619, A2 => n18620, A3 => n18621, A4 => 
                           n18622, ZN => n18618);
   U18557 : NAND4_X1 port map( A1 => n18627, A2 => n18628, A3 => n18629, A4 => 
                           n18630, ZN => n18617);
   U18558 : OAI21_X1 port map( B1 => n4282, B2 => n18417, A => n18579, ZN => 
                           n5370);
   U18559 : OAI21_X1 port map( B1 => n18580, B2 => n18581, A => n18417, ZN => 
                           n18579);
   U18560 : NAND4_X1 port map( A1 => n18582, A2 => n18583, A3 => n18584, A4 => 
                           n18585, ZN => n18581);
   U18561 : NAND4_X1 port map( A1 => n18590, A2 => n18591, A3 => n18592, A4 => 
                           n18593, ZN => n18580);
   U18562 : OAI21_X1 port map( B1 => n4283, B2 => n18417, A => n18542, ZN => 
                           n5371);
   U18563 : OAI21_X1 port map( B1 => n18543, B2 => n18544, A => n18417, ZN => 
                           n18542);
   U18564 : NAND4_X1 port map( A1 => n18545, A2 => n18546, A3 => n18547, A4 => 
                           n18548, ZN => n18544);
   U18565 : NAND4_X1 port map( A1 => n18553, A2 => n18554, A3 => n18555, A4 => 
                           n18556, ZN => n18543);
   U18566 : OAI21_X1 port map( B1 => n4284, B2 => n18417, A => n18505, ZN => 
                           n5372);
   U18567 : OAI21_X1 port map( B1 => n18506, B2 => n18507, A => n18417, ZN => 
                           n18505);
   U18568 : NAND4_X1 port map( A1 => n18508, A2 => n18509, A3 => n18510, A4 => 
                           n18511, ZN => n18507);
   U18569 : NAND4_X1 port map( A1 => n18516, A2 => n18517, A3 => n18518, A4 => 
                           n18519, ZN => n18506);
   U18570 : OAI21_X1 port map( B1 => n4285, B2 => n18417, A => n18418, ZN => 
                           n5373);
   U18571 : OAI21_X1 port map( B1 => n18419, B2 => n18420, A => n18417, ZN => 
                           n18418);
   U18572 : NAND4_X1 port map( A1 => n18421, A2 => n18422, A3 => n18423, A4 => 
                           n18424, ZN => n18420);
   U18573 : NAND4_X1 port map( A1 => n18446, A2 => n18447, A3 => n18448, A4 => 
                           n18449, ZN => n18419);
   U18574 : OAI21_X1 port map( B1 => n4288, B2 => n16834, A => n18295, ZN => 
                           n5376);
   U18575 : OAI21_X1 port map( B1 => n18296, B2 => n18297, A => n16834, ZN => 
                           n18295);
   U18576 : NAND4_X1 port map( A1 => n18298, A2 => n18299, A3 => n18300, A4 => 
                           n18301, ZN => n18297);
   U18577 : NAND4_X1 port map( A1 => n18307, A2 => n18308, A3 => n18309, A4 => 
                           n18310, ZN => n18296);
   U18578 : OAI21_X1 port map( B1 => n4290, B2 => n16834, A => n18248, ZN => 
                           n5378);
   U18579 : OAI21_X1 port map( B1 => n18249, B2 => n18250, A => n16834, ZN => 
                           n18248);
   U18580 : NAND4_X1 port map( A1 => n18251, A2 => n18252, A3 => n18253, A4 => 
                           n18254, ZN => n18250);
   U18581 : NAND4_X1 port map( A1 => n18260, A2 => n18261, A3 => n18262, A4 => 
                           n18263, ZN => n18249);
   U18582 : OAI21_X1 port map( B1 => n4292, B2 => n16834, A => n18201, ZN => 
                           n5380);
   U18583 : OAI21_X1 port map( B1 => n18202, B2 => n18203, A => n16834, ZN => 
                           n18201);
   U18584 : NAND4_X1 port map( A1 => n18204, A2 => n18205, A3 => n18206, A4 => 
                           n18207, ZN => n18203);
   U18585 : NAND4_X1 port map( A1 => n18213, A2 => n18214, A3 => n18215, A4 => 
                           n18216, ZN => n18202);
   U18586 : OAI21_X1 port map( B1 => n4294, B2 => n16834, A => n18154, ZN => 
                           n5382);
   U18587 : OAI21_X1 port map( B1 => n18155, B2 => n18156, A => n16834, ZN => 
                           n18154);
   U18588 : NAND4_X1 port map( A1 => n18157, A2 => n18158, A3 => n18159, A4 => 
                           n18160, ZN => n18156);
   U18589 : NAND4_X1 port map( A1 => n18166, A2 => n18167, A3 => n18168, A4 => 
                           n18169, ZN => n18155);
   U18590 : OAI21_X1 port map( B1 => n4296, B2 => n16834, A => n18107, ZN => 
                           n5384);
   U18591 : OAI21_X1 port map( B1 => n18108, B2 => n18109, A => n16834, ZN => 
                           n18107);
   U18592 : NAND4_X1 port map( A1 => n18110, A2 => n18111, A3 => n18112, A4 => 
                           n18113, ZN => n18109);
   U18593 : NAND4_X1 port map( A1 => n18119, A2 => n18120, A3 => n18121, A4 => 
                           n18122, ZN => n18108);
   U18594 : OAI21_X1 port map( B1 => n4298, B2 => n16834, A => n18060, ZN => 
                           n5386);
   U18595 : OAI21_X1 port map( B1 => n18061, B2 => n18062, A => n16834, ZN => 
                           n18060);
   U18596 : NAND4_X1 port map( A1 => n18063, A2 => n18064, A3 => n18065, A4 => 
                           n18066, ZN => n18062);
   U18597 : NAND4_X1 port map( A1 => n18072, A2 => n18073, A3 => n18074, A4 => 
                           n18075, ZN => n18061);
   U18598 : OAI21_X1 port map( B1 => n4300, B2 => n16834, A => n18013, ZN => 
                           n5388);
   U18599 : OAI21_X1 port map( B1 => n18014, B2 => n18015, A => n16834, ZN => 
                           n18013);
   U18600 : NAND4_X1 port map( A1 => n18016, A2 => n18017, A3 => n18018, A4 => 
                           n18019, ZN => n18015);
   U18601 : NAND4_X1 port map( A1 => n18025, A2 => n18026, A3 => n18027, A4 => 
                           n18028, ZN => n18014);
   U18602 : OAI21_X1 port map( B1 => n4302, B2 => n16834, A => n17966, ZN => 
                           n5390);
   U18603 : OAI21_X1 port map( B1 => n17967, B2 => n17968, A => n16834, ZN => 
                           n17966);
   U18604 : NAND4_X1 port map( A1 => n17969, A2 => n17970, A3 => n17971, A4 => 
                           n17972, ZN => n17968);
   U18605 : NAND4_X1 port map( A1 => n17978, A2 => n17979, A3 => n17980, A4 => 
                           n17981, ZN => n17967);
   U18606 : OAI21_X1 port map( B1 => n4304, B2 => n16834, A => n17919, ZN => 
                           n5392);
   U18607 : OAI21_X1 port map( B1 => n17920, B2 => n17921, A => n16834, ZN => 
                           n17919);
   U18608 : NAND4_X1 port map( A1 => n17922, A2 => n17923, A3 => n17924, A4 => 
                           n17925, ZN => n17921);
   U18609 : NAND4_X1 port map( A1 => n17931, A2 => n17932, A3 => n17933, A4 => 
                           n17934, ZN => n17920);
   U18610 : OAI21_X1 port map( B1 => n4306, B2 => n16834, A => n17872, ZN => 
                           n5394);
   U18611 : OAI21_X1 port map( B1 => n17873, B2 => n17874, A => n16834, ZN => 
                           n17872);
   U18612 : NAND4_X1 port map( A1 => n17875, A2 => n17876, A3 => n17877, A4 => 
                           n17878, ZN => n17874);
   U18613 : NAND4_X1 port map( A1 => n17884, A2 => n17885, A3 => n17886, A4 => 
                           n17887, ZN => n17873);
   U18614 : OAI21_X1 port map( B1 => n4308, B2 => n16834, A => n17825, ZN => 
                           n5396);
   U18615 : OAI21_X1 port map( B1 => n17826, B2 => n17827, A => n16834, ZN => 
                           n17825);
   U18616 : NAND4_X1 port map( A1 => n17828, A2 => n17829, A3 => n17830, A4 => 
                           n17831, ZN => n17827);
   U18617 : NAND4_X1 port map( A1 => n17837, A2 => n17838, A3 => n17839, A4 => 
                           n17840, ZN => n17826);
   U18618 : OAI21_X1 port map( B1 => n4310, B2 => n16834, A => n17778, ZN => 
                           n5398);
   U18619 : OAI21_X1 port map( B1 => n17779, B2 => n17780, A => n16834, ZN => 
                           n17778);
   U18620 : NAND4_X1 port map( A1 => n17781, A2 => n17782, A3 => n17783, A4 => 
                           n17784, ZN => n17780);
   U18621 : NAND4_X1 port map( A1 => n17790, A2 => n17791, A3 => n17792, A4 => 
                           n17793, ZN => n17779);
   U18622 : OAI21_X1 port map( B1 => n4312, B2 => n16834, A => n17731, ZN => 
                           n5400);
   U18623 : OAI21_X1 port map( B1 => n17732, B2 => n17733, A => n16834, ZN => 
                           n17731);
   U18624 : NAND4_X1 port map( A1 => n17734, A2 => n17735, A3 => n17736, A4 => 
                           n17737, ZN => n17733);
   U18625 : NAND4_X1 port map( A1 => n17743, A2 => n17744, A3 => n17745, A4 => 
                           n17746, ZN => n17732);
   U18626 : OAI21_X1 port map( B1 => n4314, B2 => n16834, A => n17684, ZN => 
                           n5402);
   U18627 : OAI21_X1 port map( B1 => n17685, B2 => n17686, A => n16834, ZN => 
                           n17684);
   U18628 : NAND4_X1 port map( A1 => n17687, A2 => n17688, A3 => n17689, A4 => 
                           n17690, ZN => n17686);
   U18629 : NAND4_X1 port map( A1 => n17696, A2 => n17697, A3 => n17698, A4 => 
                           n17699, ZN => n17685);
   U18630 : OAI21_X1 port map( B1 => n4316, B2 => n16834, A => n17637, ZN => 
                           n5404);
   U18631 : OAI21_X1 port map( B1 => n17638, B2 => n17639, A => n16834, ZN => 
                           n17637);
   U18632 : NAND4_X1 port map( A1 => n17640, A2 => n17641, A3 => n17642, A4 => 
                           n17643, ZN => n17639);
   U18633 : NAND4_X1 port map( A1 => n17649, A2 => n17650, A3 => n17651, A4 => 
                           n17652, ZN => n17638);
   U18634 : OAI21_X1 port map( B1 => n4318, B2 => n16834, A => n17590, ZN => 
                           n5406);
   U18635 : OAI21_X1 port map( B1 => n17591, B2 => n17592, A => n16834, ZN => 
                           n17590);
   U18636 : NAND4_X1 port map( A1 => n17593, A2 => n17594, A3 => n17595, A4 => 
                           n17596, ZN => n17592);
   U18637 : NAND4_X1 port map( A1 => n17602, A2 => n17603, A3 => n17604, A4 => 
                           n17605, ZN => n17591);
   U18638 : OAI21_X1 port map( B1 => n4320, B2 => n16834, A => n17543, ZN => 
                           n5408);
   U18639 : OAI21_X1 port map( B1 => n17544, B2 => n17545, A => n16834, ZN => 
                           n17543);
   U18640 : NAND4_X1 port map( A1 => n17546, A2 => n17547, A3 => n17548, A4 => 
                           n17549, ZN => n17545);
   U18641 : NAND4_X1 port map( A1 => n17555, A2 => n17556, A3 => n17557, A4 => 
                           n17558, ZN => n17544);
   U18642 : OAI21_X1 port map( B1 => n4322, B2 => n16834, A => n17496, ZN => 
                           n5410);
   U18643 : OAI21_X1 port map( B1 => n17497, B2 => n17498, A => n16834, ZN => 
                           n17496);
   U18644 : NAND4_X1 port map( A1 => n17499, A2 => n17500, A3 => n17501, A4 => 
                           n17502, ZN => n17498);
   U18645 : NAND4_X1 port map( A1 => n17508, A2 => n17509, A3 => n17510, A4 => 
                           n17511, ZN => n17497);
   U18646 : OAI21_X1 port map( B1 => n4324, B2 => n16834, A => n17449, ZN => 
                           n5412);
   U18647 : OAI21_X1 port map( B1 => n17450, B2 => n17451, A => n16834, ZN => 
                           n17449);
   U18648 : NAND4_X1 port map( A1 => n17452, A2 => n17453, A3 => n17454, A4 => 
                           n17455, ZN => n17451);
   U18649 : NAND4_X1 port map( A1 => n17461, A2 => n17462, A3 => n17463, A4 => 
                           n17464, ZN => n17450);
   U18650 : OAI21_X1 port map( B1 => n4326, B2 => n16834, A => n17402, ZN => 
                           n5414);
   U18651 : OAI21_X1 port map( B1 => n17403, B2 => n17404, A => n16834, ZN => 
                           n17402);
   U18652 : NAND4_X1 port map( A1 => n17405, A2 => n17406, A3 => n17407, A4 => 
                           n17408, ZN => n17404);
   U18653 : NAND4_X1 port map( A1 => n17414, A2 => n17415, A3 => n17416, A4 => 
                           n17417, ZN => n17403);
   U18654 : OAI21_X1 port map( B1 => n4328, B2 => n16834, A => n17355, ZN => 
                           n5416);
   U18655 : OAI21_X1 port map( B1 => n17356, B2 => n17357, A => n16834, ZN => 
                           n17355);
   U18656 : NAND4_X1 port map( A1 => n17358, A2 => n17359, A3 => n17360, A4 => 
                           n17361, ZN => n17357);
   U18657 : NAND4_X1 port map( A1 => n17367, A2 => n17368, A3 => n17369, A4 => 
                           n17370, ZN => n17356);
   U18658 : OAI21_X1 port map( B1 => n4330, B2 => n16834, A => n17308, ZN => 
                           n5418);
   U18659 : OAI21_X1 port map( B1 => n17309, B2 => n17310, A => n16834, ZN => 
                           n17308);
   U18660 : NAND4_X1 port map( A1 => n17311, A2 => n17312, A3 => n17313, A4 => 
                           n17314, ZN => n17310);
   U18661 : NAND4_X1 port map( A1 => n17320, A2 => n17321, A3 => n17322, A4 => 
                           n17323, ZN => n17309);
   U18662 : OAI21_X1 port map( B1 => n4332, B2 => n16834, A => n17261, ZN => 
                           n5420);
   U18663 : OAI21_X1 port map( B1 => n17262, B2 => n17263, A => n16834, ZN => 
                           n17261);
   U18664 : NAND4_X1 port map( A1 => n17264, A2 => n17265, A3 => n17266, A4 => 
                           n17267, ZN => n17263);
   U18665 : NAND4_X1 port map( A1 => n17273, A2 => n17274, A3 => n17275, A4 => 
                           n17276, ZN => n17262);
   U18666 : OAI21_X1 port map( B1 => n4334, B2 => n16834, A => n17214, ZN => 
                           n5422);
   U18667 : OAI21_X1 port map( B1 => n17215, B2 => n17216, A => n16834, ZN => 
                           n17214);
   U18668 : NAND4_X1 port map( A1 => n17217, A2 => n17218, A3 => n17219, A4 => 
                           n17220, ZN => n17216);
   U18669 : NAND4_X1 port map( A1 => n17226, A2 => n17227, A3 => n17228, A4 => 
                           n17229, ZN => n17215);
   U18670 : OAI21_X1 port map( B1 => n4336, B2 => n16834, A => n17167, ZN => 
                           n5424);
   U18671 : OAI21_X1 port map( B1 => n17168, B2 => n17169, A => n16834, ZN => 
                           n17167);
   U18672 : NAND4_X1 port map( A1 => n17170, A2 => n17171, A3 => n17172, A4 => 
                           n17173, ZN => n17169);
   U18673 : NAND4_X1 port map( A1 => n17179, A2 => n17180, A3 => n17181, A4 => 
                           n17182, ZN => n17168);
   U18674 : OAI21_X1 port map( B1 => n4338, B2 => n16834, A => n17120, ZN => 
                           n5426);
   U18675 : OAI21_X1 port map( B1 => n17121, B2 => n17122, A => n16834, ZN => 
                           n17120);
   U18676 : NAND4_X1 port map( A1 => n17123, A2 => n17124, A3 => n17125, A4 => 
                           n17126, ZN => n17122);
   U18677 : NAND4_X1 port map( A1 => n17132, A2 => n17133, A3 => n17134, A4 => 
                           n17135, ZN => n17121);
   U18678 : OAI21_X1 port map( B1 => n4340, B2 => n16834, A => n17073, ZN => 
                           n5428);
   U18679 : OAI21_X1 port map( B1 => n17074, B2 => n17075, A => n16834, ZN => 
                           n17073);
   U18680 : NAND4_X1 port map( A1 => n17076, A2 => n17077, A3 => n17078, A4 => 
                           n17079, ZN => n17075);
   U18681 : NAND4_X1 port map( A1 => n17085, A2 => n17086, A3 => n17087, A4 => 
                           n17088, ZN => n17074);
   U18682 : OAI21_X1 port map( B1 => n4342, B2 => n16834, A => n17026, ZN => 
                           n5430);
   U18683 : OAI21_X1 port map( B1 => n17027, B2 => n17028, A => n16834, ZN => 
                           n17026);
   U18684 : NAND4_X1 port map( A1 => n17029, A2 => n17030, A3 => n17031, A4 => 
                           n17032, ZN => n17028);
   U18685 : NAND4_X1 port map( A1 => n17038, A2 => n17039, A3 => n17040, A4 => 
                           n17041, ZN => n17027);
   U18686 : OAI21_X1 port map( B1 => n4344, B2 => n16834, A => n16979, ZN => 
                           n5432);
   U18687 : OAI21_X1 port map( B1 => n16980, B2 => n16981, A => n16834, ZN => 
                           n16979);
   U18688 : NAND4_X1 port map( A1 => n16982, A2 => n16983, A3 => n16984, A4 => 
                           n16985, ZN => n16981);
   U18689 : NAND4_X1 port map( A1 => n16991, A2 => n16992, A3 => n16993, A4 => 
                           n16994, ZN => n16980);
   U18690 : OAI21_X1 port map( B1 => n4346, B2 => n16834, A => n16932, ZN => 
                           n5434);
   U18691 : OAI21_X1 port map( B1 => n16933, B2 => n16934, A => n16834, ZN => 
                           n16932);
   U18692 : NAND4_X1 port map( A1 => n16935, A2 => n16936, A3 => n16937, A4 => 
                           n16938, ZN => n16934);
   U18693 : NAND4_X1 port map( A1 => n16944, A2 => n16945, A3 => n16946, A4 => 
                           n16947, ZN => n16933);
   U18694 : OAI21_X1 port map( B1 => n4348, B2 => n16834, A => n16835, ZN => 
                           n5436);
   U18695 : OAI21_X1 port map( B1 => n16836, B2 => n16837, A => n16834, ZN => 
                           n16835);
   U18696 : NAND4_X1 port map( A1 => n16838, A2 => n16839, A3 => n16840, A4 => 
                           n16841, ZN => n16837);
   U18697 : NAND4_X1 port map( A1 => n16864, A2 => n16865, A3 => n16866, A4 => 
                           n16867, ZN => n16836);
   U18698 : AND2_X1 port map( A1 => n19677, A2 => ADD_RD1(2), ZN => n20751);
   U18699 : AND2_X1 port map( A1 => n19670, A2 => ADD_RD1(2), ZN => n20903);
   U18700 : AND2_X1 port map( A1 => n19662, A2 => ADD_RD1(2), ZN => n21038);
   U18701 : AND2_X1 port map( A1 => n18414, A2 => ADD_RD2(2), ZN => n21308);
   U18702 : AND2_X1 port map( A1 => n18405, A2 => ADD_RD2(2), ZN => n21460);
   U18703 : AND2_X1 port map( A1 => n18395, A2 => ADD_RD2(2), ZN => n21595);
   U18704 : AND2_X1 port map( A1 => n19662, A2 => ADD_RD1(2), ZN => n18465);
   U18705 : AND2_X1 port map( A1 => n19677, A2 => ADD_RD1(2), ZN => n18475);
   U18706 : AND2_X1 port map( A1 => n19670, A2 => ADD_RD1(2), ZN => n18481);
   U18707 : AND2_X1 port map( A1 => n18395, A2 => ADD_RD2(2), ZN => n16884);
   U18708 : AND2_X1 port map( A1 => n18414, A2 => ADD_RD2(2), ZN => n16896);
   U18709 : AND2_X1 port map( A1 => n18405, A2 => ADD_RD2(2), ZN => n16903);
   U18710 : AND2_X1 port map( A1 => n19663, A2 => ADD_RD1(2), ZN => n20687);
   U18711 : AND2_X1 port map( A1 => n18396, A2 => ADD_RD2(2), ZN => n21244);
   U18712 : AND2_X1 port map( A1 => n19663, A2 => ADD_RD1(2), ZN => n18471);
   U18713 : AND2_X1 port map( A1 => n18396, A2 => ADD_RD2(2), ZN => n16892);
   U18714 : INV_X1 port map( A => ADD_WR(0), ZN => n16795);
   U18715 : INV_X1 port map( A => ADD_WR(1), ZN => n16794);
   U18716 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n15645);
   U18717 : INV_X1 port map( A => n19632, ZN => n19631);
   U18718 : OAI222_X1 port map( A1 => n21161, A2 => n15927, B1 => n21174, B2 =>
                           n4510, C1 => n21177, C2 => n4478, ZN => n19632);
   U18719 : INV_X1 port map( A => n18359, ZN => n18358);
   U18720 : OAI222_X1 port map( A1 => n21718, A2 => n15927, B1 => n21731, B2 =>
                           n4510, C1 => n21734, C2 => n4478, ZN => n18359);
   U18721 : INV_X1 port map( A => n19621, ZN => n19620);
   U18722 : AOI221_X1 port map( B1 => n8573, B2 => n18441, C1 => n9021, C2 => 
                           n18442, A => n19622, ZN => n19621);
   U18723 : OAI22_X1 port map( A1 => n18445, A2 => n15469, B1 => n18444, B2 => 
                           n15503, ZN => n19622);
   U18724 : INV_X1 port map( A => n18348, ZN => n18347);
   U18725 : AOI221_X1 port map( B1 => n8573, B2 => n16859, C1 => n9021, C2 => 
                           n16860, A => n18349, ZN => n18348);
   U18726 : OAI22_X1 port map( A1 => n16863, A2 => n15469, B1 => n16862, B2 => 
                           n15503, ZN => n18349);
   U18727 : INV_X1 port map( A => ADD_WR(2), ZN => n16653);
   U18728 : INV_X1 port map( A => ADD_WR(5), ZN => n15644);
   U18729 : INV_X1 port map( A => ADD_WR(4), ZN => n15643);
   U18730 : INV_X1 port map( A => RESET, ZN => n15153);
   U18731 : INV_X1 port map( A => n20687, ZN => n20688);
   U18732 : INV_X1 port map( A => n20687, ZN => n20689);
   U18733 : INV_X1 port map( A => n20687, ZN => n20690);
   U18734 : INV_X1 port map( A => n20687, ZN => n20691);
   U18735 : INV_X1 port map( A => n20687, ZN => n20692);
   U18736 : INV_X1 port map( A => n20688, ZN => n20693);
   U18737 : INV_X1 port map( A => n20688, ZN => n20694);
   U18738 : INV_X1 port map( A => n20688, ZN => n20695);
   U18739 : INV_X1 port map( A => n20689, ZN => n20696);
   U18740 : INV_X1 port map( A => n20689, ZN => n20697);
   U18741 : INV_X1 port map( A => n20689, ZN => n20698);
   U18742 : INV_X1 port map( A => n20690, ZN => n20699);
   U18743 : INV_X1 port map( A => n20690, ZN => n20700);
   U18744 : INV_X1 port map( A => n20690, ZN => n20701);
   U18745 : INV_X1 port map( A => n20691, ZN => n20702);
   U18746 : INV_X1 port map( A => n20691, ZN => n20703);
   U18747 : INV_X1 port map( A => n20691, ZN => n20704);
   U18748 : INV_X1 port map( A => n20692, ZN => n20705);
   U18749 : INV_X1 port map( A => n20692, ZN => n20706);
   U18750 : INV_X1 port map( A => n20692, ZN => n20707);
   U18751 : INV_X1 port map( A => n20711, ZN => n20708);
   U18752 : INV_X1 port map( A => n18471, ZN => n20709);
   U18753 : INV_X1 port map( A => n18471, ZN => n20710);
   U18754 : INV_X1 port map( A => n18471, ZN => n20711);
   U18755 : INV_X1 port map( A => n20710, ZN => n20712);
   U18756 : INV_X1 port map( A => n20709, ZN => n20713);
   U18757 : INV_X1 port map( A => n20709, ZN => n20714);
   U18758 : INV_X1 port map( A => n20709, ZN => n20715);
   U18759 : INV_X1 port map( A => n20710, ZN => n20716);
   U18760 : INV_X1 port map( A => n20710, ZN => n20717);
   U18761 : INV_X1 port map( A => n20711, ZN => n20718);
   U18762 : INV_X1 port map( A => n20711, ZN => n20719);
   U18763 : INV_X1 port map( A => n18500, ZN => n20720);
   U18764 : INV_X1 port map( A => n18500, ZN => n20721);
   U18765 : INV_X1 port map( A => n20721, ZN => n20722);
   U18766 : INV_X1 port map( A => n20720, ZN => n20723);
   U18767 : INV_X1 port map( A => n20720, ZN => n20724);
   U18768 : INV_X1 port map( A => n20721, ZN => n20725);
   U18769 : INV_X1 port map( A => n20720, ZN => n20726);
   U18770 : INV_X1 port map( A => n20721, ZN => n20727);
   U18771 : INV_X1 port map( A => n20720, ZN => n20728);
   U18772 : INV_X1 port map( A => n18501, ZN => n20735);
   U18773 : INV_X1 port map( A => n18501, ZN => n20736);
   U18774 : INV_X1 port map( A => n20735, ZN => n20737);
   U18775 : INV_X1 port map( A => n20736, ZN => n20738);
   U18776 : INV_X1 port map( A => n20735, ZN => n20739);
   U18777 : INV_X1 port map( A => n20735, ZN => n20740);
   U18778 : INV_X1 port map( A => n20736, ZN => n20741);
   U18779 : INV_X1 port map( A => n20736, ZN => n20742);
   U18780 : INV_X1 port map( A => n20743, ZN => n20744);
   U18781 : INV_X1 port map( A => n20743, ZN => n20745);
   U18782 : INV_X1 port map( A => n20743, ZN => n20746);
   U18783 : INV_X1 port map( A => n20743, ZN => n20747);
   U18784 : INV_X1 port map( A => n20743, ZN => n20748);
   U18785 : INV_X1 port map( A => n20743, ZN => n20749);
   U18786 : INV_X1 port map( A => n20743, ZN => n20750);
   U18787 : INV_X1 port map( A => n20751, ZN => n20752);
   U18788 : INV_X1 port map( A => n20751, ZN => n20753);
   U18789 : INV_X1 port map( A => n20751, ZN => n20754);
   U18790 : INV_X1 port map( A => n20751, ZN => n20755);
   U18791 : INV_X1 port map( A => n20751, ZN => n20756);
   U18792 : INV_X1 port map( A => n20752, ZN => n20757);
   U18793 : INV_X1 port map( A => n20752, ZN => n20758);
   U18794 : INV_X1 port map( A => n20753, ZN => n20759);
   U18795 : INV_X1 port map( A => n20753, ZN => n20760);
   U18796 : INV_X1 port map( A => n20753, ZN => n20761);
   U18797 : INV_X1 port map( A => n20754, ZN => n20762);
   U18798 : INV_X1 port map( A => n20754, ZN => n20763);
   U18799 : INV_X1 port map( A => n20754, ZN => n20764);
   U18800 : INV_X1 port map( A => n20755, ZN => n20765);
   U18801 : INV_X1 port map( A => n20755, ZN => n20766);
   U18802 : INV_X1 port map( A => n20755, ZN => n20767);
   U18803 : INV_X1 port map( A => n20756, ZN => n20768);
   U18804 : INV_X1 port map( A => n20756, ZN => n20769);
   U18805 : INV_X1 port map( A => n20756, ZN => n20770);
   U18806 : INV_X1 port map( A => n18475, ZN => n20771);
   U18807 : INV_X1 port map( A => n18475, ZN => n20772);
   U18808 : INV_X1 port map( A => n18475, ZN => n20773);
   U18809 : INV_X1 port map( A => n18475, ZN => n20774);
   U18810 : INV_X1 port map( A => n20771, ZN => n20775);
   U18811 : INV_X1 port map( A => n20771, ZN => n20776);
   U18812 : INV_X1 port map( A => n20771, ZN => n20777);
   U18813 : INV_X1 port map( A => n20772, ZN => n20778);
   U18814 : INV_X1 port map( A => n20772, ZN => n20779);
   U18815 : INV_X1 port map( A => n20773, ZN => n20780);
   U18816 : INV_X1 port map( A => n20773, ZN => n20781);
   U18817 : INV_X1 port map( A => n20774, ZN => n20782);
   U18818 : INV_X1 port map( A => n20774, ZN => n20783);
   U18819 : INV_X1 port map( A => n20784, ZN => n20785);
   U18820 : INV_X1 port map( A => n20784, ZN => n20786);
   U18821 : INV_X1 port map( A => n20784, ZN => n20787);
   U18822 : INV_X1 port map( A => n20784, ZN => n20788);
   U18823 : INV_X1 port map( A => n20784, ZN => n20789);
   U18824 : INV_X1 port map( A => n20784, ZN => n20790);
   U18825 : INV_X1 port map( A => n20784, ZN => n20791);
   U18826 : INV_X1 port map( A => n18495, ZN => n20798);
   U18827 : INV_X1 port map( A => n18495, ZN => n20799);
   U18828 : INV_X1 port map( A => n20799, ZN => n20800);
   U18829 : INV_X1 port map( A => n20798, ZN => n20801);
   U18830 : INV_X1 port map( A => n20799, ZN => n20802);
   U18831 : INV_X1 port map( A => n20798, ZN => n20803);
   U18832 : INV_X1 port map( A => n20799, ZN => n20804);
   U18833 : INV_X1 port map( A => n20798, ZN => n20805);
   U18834 : INV_X1 port map( A => n20806, ZN => n20807);
   U18835 : INV_X1 port map( A => n20806, ZN => n20808);
   U18836 : INV_X1 port map( A => n20806, ZN => n20809);
   U18837 : INV_X1 port map( A => n20806, ZN => n20810);
   U18838 : INV_X1 port map( A => n20806, ZN => n20811);
   U18839 : INV_X1 port map( A => n20830, ZN => n20812);
   U18840 : INV_X1 port map( A => n20807, ZN => n20813);
   U18841 : INV_X1 port map( A => n20807, ZN => n20814);
   U18842 : INV_X1 port map( A => n20807, ZN => n20815);
   U18843 : INV_X1 port map( A => n20808, ZN => n20816);
   U18844 : INV_X1 port map( A => n20808, ZN => n20817);
   U18845 : INV_X1 port map( A => n20808, ZN => n20818);
   U18846 : INV_X1 port map( A => n20809, ZN => n20819);
   U18847 : INV_X1 port map( A => n20809, ZN => n20820);
   U18848 : INV_X1 port map( A => n20809, ZN => n20821);
   U18849 : INV_X1 port map( A => n20810, ZN => n20822);
   U18850 : INV_X1 port map( A => n20810, ZN => n20823);
   U18851 : INV_X1 port map( A => n20810, ZN => n20824);
   U18852 : INV_X1 port map( A => n20811, ZN => n20825);
   U18853 : INV_X1 port map( A => n20811, ZN => n20826);
   U18854 : INV_X1 port map( A => n20811, ZN => n20827);
   U18855 : INV_X1 port map( A => n18476, ZN => n20828);
   U18856 : INV_X1 port map( A => n18476, ZN => n20829);
   U18857 : INV_X1 port map( A => n18476, ZN => n20830);
   U18858 : INV_X1 port map( A => n20829, ZN => n20831);
   U18859 : INV_X1 port map( A => n20828, ZN => n20832);
   U18860 : INV_X1 port map( A => n20828, ZN => n20833);
   U18861 : INV_X1 port map( A => n20828, ZN => n20834);
   U18862 : INV_X1 port map( A => n20829, ZN => n20835);
   U18863 : INV_X1 port map( A => n20829, ZN => n20836);
   U18864 : INV_X1 port map( A => n20830, ZN => n20837);
   U18865 : INV_X1 port map( A => n20830, ZN => n20838);
   U18866 : INV_X1 port map( A => n20842, ZN => n20843);
   U18867 : INV_X1 port map( A => n20842, ZN => n20844);
   U18868 : INV_X1 port map( A => n20842, ZN => n20845);
   U18869 : INV_X1 port map( A => n20842, ZN => n20846);
   U18870 : INV_X1 port map( A => n20842, ZN => n20847);
   U18871 : INV_X1 port map( A => n20842, ZN => n20848);
   U18872 : INV_X1 port map( A => n20842, ZN => n20849);
   U18873 : INV_X1 port map( A => n20850, ZN => n20852);
   U18874 : INV_X1 port map( A => n20851, ZN => n20853);
   U18875 : INV_X1 port map( A => n20850, ZN => n20854);
   U18876 : INV_X1 port map( A => n20851, ZN => n20855);
   U18877 : INV_X1 port map( A => n20850, ZN => n20856);
   U18878 : INV_X1 port map( A => n20851, ZN => n20857);
   U18879 : INV_X1 port map( A => n20851, ZN => n20858);
   U18880 : INV_X1 port map( A => n18490, ZN => n20865);
   U18881 : INV_X1 port map( A => n20865, ZN => n20866);
   U18882 : INV_X1 port map( A => n20865, ZN => n20867);
   U18883 : INV_X1 port map( A => n20865, ZN => n20868);
   U18884 : INV_X1 port map( A => n20865, ZN => n20869);
   U18885 : INV_X1 port map( A => n20865, ZN => n20870);
   U18886 : INV_X1 port map( A => n20865, ZN => n20871);
   U18887 : INV_X1 port map( A => n20865, ZN => n20872);
   U18888 : INV_X1 port map( A => n18491, ZN => n20879);
   U18889 : INV_X1 port map( A => n18491, ZN => n20880);
   U18890 : INV_X1 port map( A => n20879, ZN => n20881);
   U18891 : INV_X1 port map( A => n20880, ZN => n20882);
   U18892 : INV_X1 port map( A => n20879, ZN => n20883);
   U18893 : INV_X1 port map( A => n20879, ZN => n20884);
   U18894 : INV_X1 port map( A => n20880, ZN => n20885);
   U18895 : INV_X1 port map( A => n20880, ZN => n20886);
   U18896 : INV_X1 port map( A => n20887, ZN => n20888);
   U18897 : INV_X1 port map( A => n20887, ZN => n20889);
   U18898 : INV_X1 port map( A => n20887, ZN => n20890);
   U18899 : INV_X1 port map( A => n20887, ZN => n20891);
   U18900 : INV_X1 port map( A => n20887, ZN => n20892);
   U18901 : INV_X1 port map( A => n20887, ZN => n20893);
   U18902 : INV_X1 port map( A => n20887, ZN => n20894);
   U18903 : INV_X1 port map( A => n20895, ZN => n20896);
   U18904 : INV_X1 port map( A => n20895, ZN => n20897);
   U18905 : INV_X1 port map( A => n20895, ZN => n20898);
   U18906 : INV_X1 port map( A => n20895, ZN => n20899);
   U18907 : INV_X1 port map( A => n20895, ZN => n20900);
   U18908 : INV_X1 port map( A => n20895, ZN => n20901);
   U18909 : INV_X1 port map( A => n20895, ZN => n20902);
   U18910 : INV_X1 port map( A => n20903, ZN => n20904);
   U18911 : INV_X1 port map( A => n20903, ZN => n20905);
   U18912 : INV_X1 port map( A => n20903, ZN => n20906);
   U18913 : INV_X1 port map( A => n20903, ZN => n20907);
   U18914 : INV_X1 port map( A => n20903, ZN => n20908);
   U18915 : INV_X1 port map( A => n20927, ZN => n20909);
   U18916 : INV_X1 port map( A => n20904, ZN => n20910);
   U18917 : INV_X1 port map( A => n20904, ZN => n20911);
   U18918 : INV_X1 port map( A => n20904, ZN => n20912);
   U18919 : INV_X1 port map( A => n20905, ZN => n20913);
   U18920 : INV_X1 port map( A => n20905, ZN => n20914);
   U18921 : INV_X1 port map( A => n20905, ZN => n20915);
   U18922 : INV_X1 port map( A => n20906, ZN => n20916);
   U18923 : INV_X1 port map( A => n20906, ZN => n20917);
   U18924 : INV_X1 port map( A => n20906, ZN => n20918);
   U18925 : INV_X1 port map( A => n20907, ZN => n20919);
   U18926 : INV_X1 port map( A => n20907, ZN => n20920);
   U18927 : INV_X1 port map( A => n20907, ZN => n20921);
   U18928 : INV_X1 port map( A => n20908, ZN => n20922);
   U18929 : INV_X1 port map( A => n20908, ZN => n20923);
   U18930 : INV_X1 port map( A => n20908, ZN => n20924);
   U18931 : INV_X1 port map( A => n18481, ZN => n20925);
   U18932 : INV_X1 port map( A => n18481, ZN => n20926);
   U18933 : INV_X1 port map( A => n18481, ZN => n20927);
   U18934 : INV_X1 port map( A => n20926, ZN => n20928);
   U18935 : INV_X1 port map( A => n20925, ZN => n20929);
   U18936 : INV_X1 port map( A => n20925, ZN => n20930);
   U18937 : INV_X1 port map( A => n20925, ZN => n20931);
   U18938 : INV_X1 port map( A => n20926, ZN => n20932);
   U18939 : INV_X1 port map( A => n20926, ZN => n20933);
   U18940 : INV_X1 port map( A => n20927, ZN => n20934);
   U18941 : INV_X1 port map( A => n20927, ZN => n20935);
   U18942 : INV_X1 port map( A => n18450, ZN => n20936);
   U18943 : INV_X1 port map( A => n18450, ZN => n20937);
   U18944 : INV_X1 port map( A => n20936, ZN => n20938);
   U18945 : INV_X1 port map( A => n20936, ZN => n20939);
   U18946 : INV_X1 port map( A => n20937, ZN => n20940);
   U18947 : INV_X1 port map( A => n20936, ZN => n20941);
   U18948 : INV_X1 port map( A => n20936, ZN => n20942);
   U18949 : INV_X1 port map( A => n20937, ZN => n20943);
   U18950 : INV_X1 port map( A => n20937, ZN => n20944);
   U18951 : INV_X1 port map( A => n20945, ZN => n20946);
   U18952 : INV_X1 port map( A => n20945, ZN => n20947);
   U18953 : INV_X1 port map( A => n20945, ZN => n20948);
   U18954 : INV_X1 port map( A => n20945, ZN => n20949);
   U18955 : INV_X1 port map( A => n20945, ZN => n20950);
   U18956 : INV_X1 port map( A => n20966, ZN => n20951);
   U18957 : INV_X1 port map( A => n20946, ZN => n20952);
   U18958 : INV_X1 port map( A => n20946, ZN => n20953);
   U18959 : INV_X1 port map( A => n20946, ZN => n20954);
   U18960 : INV_X1 port map( A => n20947, ZN => n20955);
   U18961 : INV_X1 port map( A => n20947, ZN => n20956);
   U18962 : INV_X1 port map( A => n20947, ZN => n20957);
   U18963 : INV_X1 port map( A => n20948, ZN => n20958);
   U18964 : INV_X1 port map( A => n20948, ZN => n20959);
   U18965 : INV_X1 port map( A => n20948, ZN => n20960);
   U18966 : INV_X1 port map( A => n20949, ZN => n20961);
   U18967 : INV_X1 port map( A => n20949, ZN => n20962);
   U18968 : INV_X1 port map( A => n20949, ZN => n20963);
   U18969 : INV_X1 port map( A => n20950, ZN => n20964);
   U18970 : INV_X1 port map( A => n18480, ZN => n20965);
   U18971 : INV_X1 port map( A => n18480, ZN => n20966);
   U18972 : INV_X1 port map( A => n18480, ZN => n20967);
   U18973 : INV_X1 port map( A => n18480, ZN => n20968);
   U18974 : INV_X1 port map( A => n20967, ZN => n20969);
   U18975 : INV_X1 port map( A => n20965, ZN => n20970);
   U18976 : INV_X1 port map( A => n20965, ZN => n20971);
   U18977 : INV_X1 port map( A => n20966, ZN => n20972);
   U18978 : INV_X1 port map( A => n20966, ZN => n20973);
   U18979 : INV_X1 port map( A => n20967, ZN => n20974);
   U18980 : INV_X1 port map( A => n20967, ZN => n20975);
   U18981 : INV_X1 port map( A => n20968, ZN => n20976);
   U18982 : INV_X1 port map( A => n20968, ZN => n20977);
   U18983 : INV_X1 port map( A => n20993, ZN => n20994);
   U18984 : INV_X1 port map( A => n20993, ZN => n20995);
   U18985 : INV_X1 port map( A => n20993, ZN => n20996);
   U18986 : INV_X1 port map( A => n20993, ZN => n20997);
   U18987 : INV_X1 port map( A => n20993, ZN => n20998);
   U18988 : INV_X1 port map( A => n20994, ZN => n20999);
   U18989 : INV_X1 port map( A => n20995, ZN => n21000);
   U18990 : INV_X1 port map( A => n20995, ZN => n21001);
   U18991 : INV_X1 port map( A => n20995, ZN => n21002);
   U18992 : INV_X1 port map( A => n20996, ZN => n21003);
   U18993 : INV_X1 port map( A => n20996, ZN => n21004);
   U18994 : INV_X1 port map( A => n20996, ZN => n21005);
   U18995 : INV_X1 port map( A => n20997, ZN => n21006);
   U18996 : INV_X1 port map( A => n20997, ZN => n21007);
   U18997 : INV_X1 port map( A => n20997, ZN => n21008);
   U18998 : INV_X1 port map( A => n20998, ZN => n21009);
   U18999 : INV_X1 port map( A => n20998, ZN => n21010);
   U19000 : INV_X1 port map( A => n20998, ZN => n21011);
   U19001 : INV_X1 port map( A => n21014, ZN => n21012);
   U19002 : INV_X1 port map( A => n18470, ZN => n21013);
   U19003 : INV_X1 port map( A => n18470, ZN => n21014);
   U19004 : INV_X1 port map( A => n18470, ZN => n21015);
   U19005 : INV_X1 port map( A => n18470, ZN => n21016);
   U19006 : INV_X1 port map( A => n21013, ZN => n21017);
   U19007 : INV_X1 port map( A => n21013, ZN => n21018);
   U19008 : INV_X1 port map( A => n21014, ZN => n21019);
   U19009 : INV_X1 port map( A => n21014, ZN => n21020);
   U19010 : INV_X1 port map( A => n21015, ZN => n21021);
   U19011 : INV_X1 port map( A => n21015, ZN => n21022);
   U19012 : INV_X1 port map( A => n21013, ZN => n21023);
   U19013 : INV_X1 port map( A => n21016, ZN => n21024);
   U19014 : INV_X1 port map( A => n21016, ZN => n21025);
   U19015 : INV_X1 port map( A => n21038, ZN => n21039);
   U19016 : INV_X1 port map( A => n21038, ZN => n21040);
   U19017 : INV_X1 port map( A => n21038, ZN => n21041);
   U19018 : INV_X1 port map( A => n21038, ZN => n21042);
   U19019 : INV_X1 port map( A => n21038, ZN => n21043);
   U19020 : INV_X1 port map( A => n21039, ZN => n21044);
   U19021 : INV_X1 port map( A => n21039, ZN => n21045);
   U19022 : INV_X1 port map( A => n21040, ZN => n21046);
   U19023 : INV_X1 port map( A => n21040, ZN => n21047);
   U19024 : INV_X1 port map( A => n21040, ZN => n21048);
   U19025 : INV_X1 port map( A => n21041, ZN => n21049);
   U19026 : INV_X1 port map( A => n21041, ZN => n21050);
   U19027 : INV_X1 port map( A => n21041, ZN => n21051);
   U19028 : INV_X1 port map( A => n21042, ZN => n21052);
   U19029 : INV_X1 port map( A => n21042, ZN => n21053);
   U19030 : INV_X1 port map( A => n21042, ZN => n21054);
   U19031 : INV_X1 port map( A => n21043, ZN => n21055);
   U19032 : INV_X1 port map( A => n21043, ZN => n21056);
   U19033 : INV_X1 port map( A => n21043, ZN => n21057);
   U19034 : INV_X1 port map( A => n18465, ZN => n21058);
   U19035 : INV_X1 port map( A => n18465, ZN => n21059);
   U19036 : INV_X1 port map( A => n18465, ZN => n21060);
   U19037 : INV_X1 port map( A => n18465, ZN => n21061);
   U19038 : INV_X1 port map( A => n21058, ZN => n21062);
   U19039 : INV_X1 port map( A => n21058, ZN => n21063);
   U19040 : INV_X1 port map( A => n21058, ZN => n21064);
   U19041 : INV_X1 port map( A => n21059, ZN => n21065);
   U19042 : INV_X1 port map( A => n21059, ZN => n21066);
   U19043 : INV_X1 port map( A => n21060, ZN => n21067);
   U19044 : INV_X1 port map( A => n21060, ZN => n21068);
   U19045 : INV_X1 port map( A => n21061, ZN => n21069);
   U19046 : INV_X1 port map( A => n21061, ZN => n21070);
   U19047 : INV_X1 port map( A => n21071, ZN => n21072);
   U19048 : INV_X1 port map( A => n21071, ZN => n21073);
   U19049 : INV_X1 port map( A => n21071, ZN => n21074);
   U19050 : INV_X1 port map( A => n21071, ZN => n21075);
   U19051 : INV_X1 port map( A => n21071, ZN => n21076);
   U19052 : INV_X1 port map( A => n21072, ZN => n21077);
   U19053 : INV_X1 port map( A => n21072, ZN => n21078);
   U19054 : INV_X1 port map( A => n21072, ZN => n21079);
   U19055 : INV_X1 port map( A => n21073, ZN => n21080);
   U19056 : INV_X1 port map( A => n21073, ZN => n21081);
   U19057 : INV_X1 port map( A => n21073, ZN => n21082);
   U19058 : INV_X1 port map( A => n21074, ZN => n21083);
   U19059 : INV_X1 port map( A => n21074, ZN => n21084);
   U19060 : INV_X1 port map( A => n21074, ZN => n21085);
   U19061 : INV_X1 port map( A => n21075, ZN => n21086);
   U19062 : INV_X1 port map( A => n21075, ZN => n21087);
   U19063 : INV_X1 port map( A => n21075, ZN => n21088);
   U19064 : INV_X1 port map( A => n21076, ZN => n21089);
   U19065 : INV_X1 port map( A => n21076, ZN => n21090);
   U19066 : INV_X1 port map( A => n21076, ZN => n21091);
   U19067 : INV_X1 port map( A => n21094, ZN => n21092);
   U19068 : INV_X1 port map( A => n18466, ZN => n21093);
   U19069 : INV_X1 port map( A => n18466, ZN => n21094);
   U19070 : INV_X1 port map( A => n18466, ZN => n21095);
   U19071 : INV_X1 port map( A => n21095, ZN => n21096);
   U19072 : INV_X1 port map( A => n21093, ZN => n21097);
   U19073 : INV_X1 port map( A => n21093, ZN => n21098);
   U19074 : INV_X1 port map( A => n21093, ZN => n21099);
   U19075 : INV_X1 port map( A => n21094, ZN => n21100);
   U19076 : INV_X1 port map( A => n21094, ZN => n21101);
   U19077 : INV_X1 port map( A => n21095, ZN => n21102);
   U19078 : INV_X1 port map( A => n21095, ZN => n21103);
   U19079 : INV_X1 port map( A => n18431, ZN => n21110);
   U19080 : INV_X1 port map( A => n18431, ZN => n21111);
   U19081 : INV_X1 port map( A => n21110, ZN => n21112);
   U19082 : INV_X1 port map( A => n21111, ZN => n21113);
   U19083 : INV_X1 port map( A => n21111, ZN => n21114);
   U19084 : INV_X1 port map( A => n21110, ZN => n21115);
   U19085 : INV_X1 port map( A => n21110, ZN => n21116);
   U19086 : INV_X1 port map( A => n21111, ZN => n21117);
   U19087 : INV_X1 port map( A => n18432, ZN => n21118);
   U19088 : INV_X1 port map( A => n18432, ZN => n21119);
   U19089 : INV_X1 port map( A => n21118, ZN => n21120);
   U19090 : INV_X1 port map( A => n21118, ZN => n21121);
   U19091 : INV_X1 port map( A => n21119, ZN => n21122);
   U19092 : INV_X1 port map( A => n21119, ZN => n21123);
   U19093 : INV_X1 port map( A => n21118, ZN => n21124);
   U19094 : INV_X1 port map( A => n21119, ZN => n21125);
   U19095 : INV_X1 port map( A => n21126, ZN => n21127);
   U19096 : INV_X1 port map( A => n21126, ZN => n21128);
   U19097 : INV_X1 port map( A => n21126, ZN => n21129);
   U19098 : INV_X1 port map( A => n21126, ZN => n21130);
   U19099 : INV_X1 port map( A => n21126, ZN => n21131);
   U19100 : INV_X1 port map( A => n21126, ZN => n21132);
   U19101 : INV_X1 port map( A => n21126, ZN => n21133);
   U19102 : INV_X1 port map( A => n21134, ZN => n21135);
   U19103 : INV_X1 port map( A => n21134, ZN => n21136);
   U19104 : INV_X1 port map( A => n21134, ZN => n21137);
   U19105 : INV_X1 port map( A => n21134, ZN => n21138);
   U19106 : INV_X1 port map( A => n21134, ZN => n21139);
   U19107 : INV_X1 port map( A => n21134, ZN => n21140);
   U19108 : INV_X1 port map( A => n21134, ZN => n21141);
   U19109 : INV_X1 port map( A => n18425, ZN => n21142);
   U19110 : INV_X1 port map( A => n18425, ZN => n21143);
   U19111 : INV_X1 port map( A => n21142, ZN => n21144);
   U19112 : INV_X1 port map( A => n21142, ZN => n21145);
   U19113 : INV_X1 port map( A => n21143, ZN => n21146);
   U19114 : INV_X1 port map( A => n21142, ZN => n21147);
   U19115 : INV_X1 port map( A => n21142, ZN => n21148);
   U19116 : INV_X1 port map( A => n21143, ZN => n21149);
   U19117 : INV_X1 port map( A => n21143, ZN => n21150);
   U19118 : INV_X1 port map( A => n18426, ZN => n21151);
   U19119 : INV_X1 port map( A => n18426, ZN => n21152);
   U19120 : INV_X1 port map( A => n21151, ZN => n21153);
   U19121 : INV_X1 port map( A => n21152, ZN => n21154);
   U19122 : INV_X1 port map( A => n21151, ZN => n21155);
   U19123 : INV_X1 port map( A => n21152, ZN => n21156);
   U19124 : INV_X1 port map( A => n21152, ZN => n21157);
   U19125 : INV_X1 port map( A => n21151, ZN => n21158);
   U19126 : INV_X1 port map( A => n21160, ZN => n21161);
   U19127 : INV_X1 port map( A => n21159, ZN => n21162);
   U19128 : INV_X1 port map( A => n21159, ZN => n21163);
   U19129 : INV_X1 port map( A => n21159, ZN => n21164);
   U19130 : INV_X1 port map( A => n21160, ZN => n21165);
   U19131 : INV_X1 port map( A => n21160, ZN => n21166);
   U19132 : INV_X1 port map( A => n21159, ZN => n21167);
   U19133 : INV_X1 port map( A => n21168, ZN => n21169);
   U19134 : INV_X1 port map( A => n21168, ZN => n21170);
   U19135 : INV_X1 port map( A => n21168, ZN => n21171);
   U19136 : INV_X1 port map( A => n21168, ZN => n21172);
   U19137 : INV_X1 port map( A => n21168, ZN => n21173);
   U19138 : INV_X1 port map( A => n21168, ZN => n21174);
   U19139 : INV_X1 port map( A => n21168, ZN => n21175);
   U19140 : INV_X1 port map( A => n21176, ZN => n21177);
   U19141 : INV_X1 port map( A => n21176, ZN => n21178);
   U19142 : INV_X1 port map( A => n21176, ZN => n21179);
   U19143 : INV_X1 port map( A => n21176, ZN => n21180);
   U19144 : INV_X1 port map( A => n21176, ZN => n21181);
   U19145 : INV_X1 port map( A => n21176, ZN => n21182);
   U19146 : INV_X1 port map( A => n21176, ZN => n21183);
   U19147 : INV_X1 port map( A => n21185, ZN => n21186);
   U19148 : INV_X1 port map( A => n21184, ZN => n21187);
   U19149 : INV_X1 port map( A => n21184, ZN => n21188);
   U19150 : INV_X1 port map( A => n21185, ZN => n21189);
   U19151 : INV_X1 port map( A => n21185, ZN => n21190);
   U19152 : INV_X1 port map( A => n21185, ZN => n21191);
   U19153 : INV_X1 port map( A => n21184, ZN => n21192);
   U19154 : INV_X1 port map( A => n21193, ZN => n21194);
   U19155 : INV_X1 port map( A => n21193, ZN => n21195);
   U19156 : INV_X1 port map( A => n21193, ZN => n21196);
   U19157 : INV_X1 port map( A => n21193, ZN => n21197);
   U19158 : INV_X1 port map( A => n21193, ZN => n21198);
   U19159 : INV_X1 port map( A => n21193, ZN => n21199);
   U19160 : INV_X1 port map( A => n21193, ZN => n21200);
   U19161 : INV_X1 port map( A => n18436, ZN => n21201);
   U19162 : INV_X1 port map( A => n18436, ZN => n21202);
   U19163 : INV_X1 port map( A => n21201, ZN => n21203);
   U19164 : INV_X1 port map( A => n21201, ZN => n21204);
   U19165 : INV_X1 port map( A => n21201, ZN => n21205);
   U19166 : INV_X1 port map( A => n21202, ZN => n21206);
   U19167 : INV_X1 port map( A => n21202, ZN => n21207);
   U19168 : INV_X1 port map( A => n21202, ZN => n21208);
   U19169 : INV_X1 port map( A => n18441, ZN => n21212);
   U19170 : INV_X1 port map( A => n21212, ZN => n21213);
   U19171 : INV_X1 port map( A => n21212, ZN => n21214);
   U19172 : INV_X1 port map( A => n21212, ZN => n21215);
   U19173 : INV_X1 port map( A => n21212, ZN => n21216);
   U19174 : INV_X1 port map( A => n21212, ZN => n21217);
   U19175 : INV_X1 port map( A => n21212, ZN => n21218);
   U19176 : INV_X1 port map( A => n21212, ZN => n21219);
   U19177 : INV_X1 port map( A => n18442, ZN => n21220);
   U19178 : INV_X1 port map( A => n21220, ZN => n21221);
   U19179 : INV_X1 port map( A => n21220, ZN => n21222);
   U19180 : INV_X1 port map( A => n21220, ZN => n21223);
   U19181 : INV_X1 port map( A => n21220, ZN => n21224);
   U19182 : INV_X1 port map( A => n21220, ZN => n21225);
   U19183 : INV_X1 port map( A => n21220, ZN => n21226);
   U19184 : INV_X1 port map( A => n21220, ZN => n21227);
   U19185 : INV_X1 port map( A => n21228, ZN => n21229);
   U19186 : INV_X1 port map( A => n21228, ZN => n21230);
   U19187 : INV_X1 port map( A => n21228, ZN => n21231);
   U19188 : INV_X1 port map( A => n21228, ZN => n21232);
   U19189 : INV_X1 port map( A => n21228, ZN => n21233);
   U19190 : INV_X1 port map( A => n21228, ZN => n21234);
   U19191 : INV_X1 port map( A => n21228, ZN => n21235);
   U19192 : INV_X1 port map( A => n21236, ZN => n21237);
   U19193 : INV_X1 port map( A => n21236, ZN => n21238);
   U19194 : INV_X1 port map( A => n21236, ZN => n21239);
   U19195 : INV_X1 port map( A => n21236, ZN => n21240);
   U19196 : INV_X1 port map( A => n21236, ZN => n21241);
   U19197 : INV_X1 port map( A => n21236, ZN => n21242);
   U19198 : INV_X1 port map( A => n21236, ZN => n21243);
   U19199 : INV_X1 port map( A => n21244, ZN => n21245);
   U19200 : INV_X1 port map( A => n21244, ZN => n21246);
   U19201 : INV_X1 port map( A => n21244, ZN => n21247);
   U19202 : INV_X1 port map( A => n21244, ZN => n21248);
   U19203 : INV_X1 port map( A => n21244, ZN => n21249);
   U19204 : INV_X1 port map( A => n21245, ZN => n21250);
   U19205 : INV_X1 port map( A => n21245, ZN => n21251);
   U19206 : INV_X1 port map( A => n21245, ZN => n21252);
   U19207 : INV_X1 port map( A => n21246, ZN => n21253);
   U19208 : INV_X1 port map( A => n21246, ZN => n21254);
   U19209 : INV_X1 port map( A => n21246, ZN => n21255);
   U19210 : INV_X1 port map( A => n21247, ZN => n21256);
   U19211 : INV_X1 port map( A => n21247, ZN => n21257);
   U19212 : INV_X1 port map( A => n21247, ZN => n21258);
   U19213 : INV_X1 port map( A => n21248, ZN => n21259);
   U19214 : INV_X1 port map( A => n21248, ZN => n21260);
   U19215 : INV_X1 port map( A => n21248, ZN => n21261);
   U19216 : INV_X1 port map( A => n21249, ZN => n21262);
   U19217 : INV_X1 port map( A => n21249, ZN => n21263);
   U19218 : INV_X1 port map( A => n21249, ZN => n21264);
   U19219 : INV_X1 port map( A => n21268, ZN => n21265);
   U19220 : INV_X1 port map( A => n16892, ZN => n21266);
   U19221 : INV_X1 port map( A => n16892, ZN => n21267);
   U19222 : INV_X1 port map( A => n16892, ZN => n21268);
   U19223 : INV_X1 port map( A => n21267, ZN => n21269);
   U19224 : INV_X1 port map( A => n21266, ZN => n21270);
   U19225 : INV_X1 port map( A => n21266, ZN => n21271);
   U19226 : INV_X1 port map( A => n21266, ZN => n21272);
   U19227 : INV_X1 port map( A => n21267, ZN => n21273);
   U19228 : INV_X1 port map( A => n21267, ZN => n21274);
   U19229 : INV_X1 port map( A => n21268, ZN => n21275);
   U19230 : INV_X1 port map( A => n21268, ZN => n21276);
   U19231 : INV_X1 port map( A => n16927, ZN => n21277);
   U19232 : INV_X1 port map( A => n16927, ZN => n21278);
   U19233 : INV_X1 port map( A => n21278, ZN => n21279);
   U19234 : INV_X1 port map( A => n21277, ZN => n21280);
   U19235 : INV_X1 port map( A => n21277, ZN => n21281);
   U19236 : INV_X1 port map( A => n21278, ZN => n21282);
   U19237 : INV_X1 port map( A => n21277, ZN => n21283);
   U19238 : INV_X1 port map( A => n21278, ZN => n21284);
   U19239 : INV_X1 port map( A => n21277, ZN => n21285);
   U19240 : INV_X1 port map( A => n16928, ZN => n21292);
   U19241 : INV_X1 port map( A => n16928, ZN => n21293);
   U19242 : INV_X1 port map( A => n21292, ZN => n21294);
   U19243 : INV_X1 port map( A => n21293, ZN => n21295);
   U19244 : INV_X1 port map( A => n21292, ZN => n21296);
   U19245 : INV_X1 port map( A => n21292, ZN => n21297);
   U19246 : INV_X1 port map( A => n21293, ZN => n21298);
   U19247 : INV_X1 port map( A => n21293, ZN => n21299);
   U19248 : INV_X1 port map( A => n21300, ZN => n21301);
   U19249 : INV_X1 port map( A => n21300, ZN => n21302);
   U19250 : INV_X1 port map( A => n21300, ZN => n21303);
   U19251 : INV_X1 port map( A => n21300, ZN => n21304);
   U19252 : INV_X1 port map( A => n21300, ZN => n21305);
   U19253 : INV_X1 port map( A => n21300, ZN => n21306);
   U19254 : INV_X1 port map( A => n21300, ZN => n21307);
   U19255 : INV_X1 port map( A => n21308, ZN => n21309);
   U19256 : INV_X1 port map( A => n21308, ZN => n21310);
   U19257 : INV_X1 port map( A => n21308, ZN => n21311);
   U19258 : INV_X1 port map( A => n21308, ZN => n21312);
   U19259 : INV_X1 port map( A => n21308, ZN => n21313);
   U19260 : INV_X1 port map( A => n21309, ZN => n21314);
   U19261 : INV_X1 port map( A => n21309, ZN => n21315);
   U19262 : INV_X1 port map( A => n21310, ZN => n21316);
   U19263 : INV_X1 port map( A => n21310, ZN => n21317);
   U19264 : INV_X1 port map( A => n21310, ZN => n21318);
   U19265 : INV_X1 port map( A => n21311, ZN => n21319);
   U19266 : INV_X1 port map( A => n21311, ZN => n21320);
   U19267 : INV_X1 port map( A => n21311, ZN => n21321);
   U19268 : INV_X1 port map( A => n21312, ZN => n21322);
   U19269 : INV_X1 port map( A => n21312, ZN => n21323);
   U19270 : INV_X1 port map( A => n21312, ZN => n21324);
   U19271 : INV_X1 port map( A => n21313, ZN => n21325);
   U19272 : INV_X1 port map( A => n21313, ZN => n21326);
   U19273 : INV_X1 port map( A => n21313, ZN => n21327);
   U19274 : INV_X1 port map( A => n16896, ZN => n21328);
   U19275 : INV_X1 port map( A => n16896, ZN => n21329);
   U19276 : INV_X1 port map( A => n16896, ZN => n21330);
   U19277 : INV_X1 port map( A => n16896, ZN => n21331);
   U19278 : INV_X1 port map( A => n21328, ZN => n21332);
   U19279 : INV_X1 port map( A => n21328, ZN => n21333);
   U19280 : INV_X1 port map( A => n21328, ZN => n21334);
   U19281 : INV_X1 port map( A => n21329, ZN => n21335);
   U19282 : INV_X1 port map( A => n21329, ZN => n21336);
   U19283 : INV_X1 port map( A => n21330, ZN => n21337);
   U19284 : INV_X1 port map( A => n21330, ZN => n21338);
   U19285 : INV_X1 port map( A => n21331, ZN => n21339);
   U19286 : INV_X1 port map( A => n21331, ZN => n21340);
   U19287 : INV_X1 port map( A => n21341, ZN => n21342);
   U19288 : INV_X1 port map( A => n21341, ZN => n21343);
   U19289 : INV_X1 port map( A => n21341, ZN => n21344);
   U19290 : INV_X1 port map( A => n21341, ZN => n21345);
   U19291 : INV_X1 port map( A => n21341, ZN => n21346);
   U19292 : INV_X1 port map( A => n21341, ZN => n21347);
   U19293 : INV_X1 port map( A => n21341, ZN => n21348);
   U19294 : INV_X1 port map( A => n16921, ZN => n21355);
   U19295 : INV_X1 port map( A => n16921, ZN => n21356);
   U19296 : INV_X1 port map( A => n21356, ZN => n21357);
   U19297 : INV_X1 port map( A => n21355, ZN => n21358);
   U19298 : INV_X1 port map( A => n21356, ZN => n21359);
   U19299 : INV_X1 port map( A => n21355, ZN => n21360);
   U19300 : INV_X1 port map( A => n21356, ZN => n21361);
   U19301 : INV_X1 port map( A => n21355, ZN => n21362);
   U19302 : INV_X1 port map( A => n21363, ZN => n21364);
   U19303 : INV_X1 port map( A => n21363, ZN => n21365);
   U19304 : INV_X1 port map( A => n21363, ZN => n21366);
   U19305 : INV_X1 port map( A => n21363, ZN => n21367);
   U19306 : INV_X1 port map( A => n21363, ZN => n21368);
   U19307 : INV_X1 port map( A => n21387, ZN => n21369);
   U19308 : INV_X1 port map( A => n21364, ZN => n21370);
   U19309 : INV_X1 port map( A => n21364, ZN => n21371);
   U19310 : INV_X1 port map( A => n21364, ZN => n21372);
   U19311 : INV_X1 port map( A => n21365, ZN => n21373);
   U19312 : INV_X1 port map( A => n21365, ZN => n21374);
   U19313 : INV_X1 port map( A => n21365, ZN => n21375);
   U19314 : INV_X1 port map( A => n21366, ZN => n21376);
   U19315 : INV_X1 port map( A => n21366, ZN => n21377);
   U19316 : INV_X1 port map( A => n21366, ZN => n21378);
   U19317 : INV_X1 port map( A => n21367, ZN => n21379);
   U19318 : INV_X1 port map( A => n21367, ZN => n21380);
   U19319 : INV_X1 port map( A => n21367, ZN => n21381);
   U19320 : INV_X1 port map( A => n21368, ZN => n21382);
   U19321 : INV_X1 port map( A => n21368, ZN => n21383);
   U19322 : INV_X1 port map( A => n21368, ZN => n21384);
   U19323 : INV_X1 port map( A => n16897, ZN => n21385);
   U19324 : INV_X1 port map( A => n16897, ZN => n21386);
   U19325 : INV_X1 port map( A => n16897, ZN => n21387);
   U19326 : INV_X1 port map( A => n21386, ZN => n21388);
   U19327 : INV_X1 port map( A => n21385, ZN => n21389);
   U19328 : INV_X1 port map( A => n21385, ZN => n21390);
   U19329 : INV_X1 port map( A => n21385, ZN => n21391);
   U19330 : INV_X1 port map( A => n21386, ZN => n21392);
   U19331 : INV_X1 port map( A => n21386, ZN => n21393);
   U19332 : INV_X1 port map( A => n21387, ZN => n21394);
   U19333 : INV_X1 port map( A => n21387, ZN => n21395);
   U19334 : INV_X1 port map( A => n21399, ZN => n21400);
   U19335 : INV_X1 port map( A => n21399, ZN => n21401);
   U19336 : INV_X1 port map( A => n21399, ZN => n21402);
   U19337 : INV_X1 port map( A => n21399, ZN => n21403);
   U19338 : INV_X1 port map( A => n21399, ZN => n21404);
   U19339 : INV_X1 port map( A => n21399, ZN => n21405);
   U19340 : INV_X1 port map( A => n21399, ZN => n21406);
   U19341 : INV_X1 port map( A => n21407, ZN => n21409);
   U19342 : INV_X1 port map( A => n21408, ZN => n21410);
   U19343 : INV_X1 port map( A => n21407, ZN => n21411);
   U19344 : INV_X1 port map( A => n21408, ZN => n21412);
   U19345 : INV_X1 port map( A => n21407, ZN => n21413);
   U19346 : INV_X1 port map( A => n21408, ZN => n21414);
   U19347 : INV_X1 port map( A => n21408, ZN => n21415);
   U19348 : INV_X1 port map( A => n16915, ZN => n21422);
   U19349 : INV_X1 port map( A => n21422, ZN => n21423);
   U19350 : INV_X1 port map( A => n21422, ZN => n21424);
   U19351 : INV_X1 port map( A => n21422, ZN => n21425);
   U19352 : INV_X1 port map( A => n21422, ZN => n21426);
   U19353 : INV_X1 port map( A => n21422, ZN => n21427);
   U19354 : INV_X1 port map( A => n21422, ZN => n21428);
   U19355 : INV_X1 port map( A => n21422, ZN => n21429);
   U19356 : INV_X1 port map( A => n16916, ZN => n21436);
   U19357 : INV_X1 port map( A => n16916, ZN => n21437);
   U19358 : INV_X1 port map( A => n21436, ZN => n21438);
   U19359 : INV_X1 port map( A => n21437, ZN => n21439);
   U19360 : INV_X1 port map( A => n21436, ZN => n21440);
   U19361 : INV_X1 port map( A => n21436, ZN => n21441);
   U19362 : INV_X1 port map( A => n21437, ZN => n21442);
   U19363 : INV_X1 port map( A => n21437, ZN => n21443);
   U19364 : INV_X1 port map( A => n21444, ZN => n21445);
   U19365 : INV_X1 port map( A => n21444, ZN => n21446);
   U19366 : INV_X1 port map( A => n21444, ZN => n21447);
   U19367 : INV_X1 port map( A => n21444, ZN => n21448);
   U19368 : INV_X1 port map( A => n21444, ZN => n21449);
   U19369 : INV_X1 port map( A => n21444, ZN => n21450);
   U19370 : INV_X1 port map( A => n21444, ZN => n21451);
   U19371 : INV_X1 port map( A => n21452, ZN => n21453);
   U19372 : INV_X1 port map( A => n21452, ZN => n21454);
   U19373 : INV_X1 port map( A => n21452, ZN => n21455);
   U19374 : INV_X1 port map( A => n21452, ZN => n21456);
   U19375 : INV_X1 port map( A => n21452, ZN => n21457);
   U19376 : INV_X1 port map( A => n21452, ZN => n21458);
   U19377 : INV_X1 port map( A => n21452, ZN => n21459);
   U19378 : INV_X1 port map( A => n21460, ZN => n21461);
   U19379 : INV_X1 port map( A => n21460, ZN => n21462);
   U19380 : INV_X1 port map( A => n21460, ZN => n21463);
   U19381 : INV_X1 port map( A => n21460, ZN => n21464);
   U19382 : INV_X1 port map( A => n21460, ZN => n21465);
   U19383 : INV_X1 port map( A => n21484, ZN => n21466);
   U19384 : INV_X1 port map( A => n21461, ZN => n21467);
   U19385 : INV_X1 port map( A => n21461, ZN => n21468);
   U19386 : INV_X1 port map( A => n21461, ZN => n21469);
   U19387 : INV_X1 port map( A => n21462, ZN => n21470);
   U19388 : INV_X1 port map( A => n21462, ZN => n21471);
   U19389 : INV_X1 port map( A => n21462, ZN => n21472);
   U19390 : INV_X1 port map( A => n21463, ZN => n21473);
   U19391 : INV_X1 port map( A => n21463, ZN => n21474);
   U19392 : INV_X1 port map( A => n21463, ZN => n21475);
   U19393 : INV_X1 port map( A => n21464, ZN => n21476);
   U19394 : INV_X1 port map( A => n21464, ZN => n21477);
   U19395 : INV_X1 port map( A => n21464, ZN => n21478);
   U19396 : INV_X1 port map( A => n21465, ZN => n21479);
   U19397 : INV_X1 port map( A => n21465, ZN => n21480);
   U19398 : INV_X1 port map( A => n21465, ZN => n21481);
   U19399 : INV_X1 port map( A => n16903, ZN => n21482);
   U19400 : INV_X1 port map( A => n16903, ZN => n21483);
   U19401 : INV_X1 port map( A => n16903, ZN => n21484);
   U19402 : INV_X1 port map( A => n21483, ZN => n21485);
   U19403 : INV_X1 port map( A => n21482, ZN => n21486);
   U19404 : INV_X1 port map( A => n21482, ZN => n21487);
   U19405 : INV_X1 port map( A => n21482, ZN => n21488);
   U19406 : INV_X1 port map( A => n21483, ZN => n21489);
   U19407 : INV_X1 port map( A => n21483, ZN => n21490);
   U19408 : INV_X1 port map( A => n21484, ZN => n21491);
   U19409 : INV_X1 port map( A => n21484, ZN => n21492);
   U19410 : INV_X1 port map( A => n16868, ZN => n21493);
   U19411 : INV_X1 port map( A => n16868, ZN => n21494);
   U19412 : INV_X1 port map( A => n21493, ZN => n21495);
   U19413 : INV_X1 port map( A => n21493, ZN => n21496);
   U19414 : INV_X1 port map( A => n21494, ZN => n21497);
   U19415 : INV_X1 port map( A => n21493, ZN => n21498);
   U19416 : INV_X1 port map( A => n21493, ZN => n21499);
   U19417 : INV_X1 port map( A => n21494, ZN => n21500);
   U19418 : INV_X1 port map( A => n21494, ZN => n21501);
   U19419 : INV_X1 port map( A => n21502, ZN => n21503);
   U19420 : INV_X1 port map( A => n21502, ZN => n21504);
   U19421 : INV_X1 port map( A => n21502, ZN => n21505);
   U19422 : INV_X1 port map( A => n21502, ZN => n21506);
   U19423 : INV_X1 port map( A => n21502, ZN => n21507);
   U19424 : INV_X1 port map( A => n21523, ZN => n21508);
   U19425 : INV_X1 port map( A => n21503, ZN => n21509);
   U19426 : INV_X1 port map( A => n21503, ZN => n21510);
   U19427 : INV_X1 port map( A => n21503, ZN => n21511);
   U19428 : INV_X1 port map( A => n21504, ZN => n21512);
   U19429 : INV_X1 port map( A => n21504, ZN => n21513);
   U19430 : INV_X1 port map( A => n21504, ZN => n21514);
   U19431 : INV_X1 port map( A => n21505, ZN => n21515);
   U19432 : INV_X1 port map( A => n21505, ZN => n21516);
   U19433 : INV_X1 port map( A => n21505, ZN => n21517);
   U19434 : INV_X1 port map( A => n21506, ZN => n21518);
   U19435 : INV_X1 port map( A => n21506, ZN => n21519);
   U19436 : INV_X1 port map( A => n21506, ZN => n21520);
   U19437 : INV_X1 port map( A => n21507, ZN => n21521);
   U19438 : INV_X1 port map( A => n16901, ZN => n21522);
   U19439 : INV_X1 port map( A => n16901, ZN => n21523);
   U19440 : INV_X1 port map( A => n16901, ZN => n21524);
   U19441 : INV_X1 port map( A => n16901, ZN => n21525);
   U19442 : INV_X1 port map( A => n21524, ZN => n21526);
   U19443 : INV_X1 port map( A => n21522, ZN => n21527);
   U19444 : INV_X1 port map( A => n21522, ZN => n21528);
   U19445 : INV_X1 port map( A => n21523, ZN => n21529);
   U19446 : INV_X1 port map( A => n21523, ZN => n21530);
   U19447 : INV_X1 port map( A => n21524, ZN => n21531);
   U19448 : INV_X1 port map( A => n21524, ZN => n21532);
   U19449 : INV_X1 port map( A => n21525, ZN => n21533);
   U19450 : INV_X1 port map( A => n21525, ZN => n21534);
   U19451 : INV_X1 port map( A => n21550, ZN => n21551);
   U19452 : INV_X1 port map( A => n21550, ZN => n21552);
   U19453 : INV_X1 port map( A => n21550, ZN => n21553);
   U19454 : INV_X1 port map( A => n21550, ZN => n21554);
   U19455 : INV_X1 port map( A => n21550, ZN => n21555);
   U19456 : INV_X1 port map( A => n21551, ZN => n21556);
   U19457 : INV_X1 port map( A => n21552, ZN => n21557);
   U19458 : INV_X1 port map( A => n21552, ZN => n21558);
   U19459 : INV_X1 port map( A => n21552, ZN => n21559);
   U19460 : INV_X1 port map( A => n21553, ZN => n21560);
   U19461 : INV_X1 port map( A => n21553, ZN => n21561);
   U19462 : INV_X1 port map( A => n21553, ZN => n21562);
   U19463 : INV_X1 port map( A => n21554, ZN => n21563);
   U19464 : INV_X1 port map( A => n21554, ZN => n21564);
   U19465 : INV_X1 port map( A => n21554, ZN => n21565);
   U19466 : INV_X1 port map( A => n21555, ZN => n21566);
   U19467 : INV_X1 port map( A => n21555, ZN => n21567);
   U19468 : INV_X1 port map( A => n21555, ZN => n21568);
   U19469 : INV_X1 port map( A => n21571, ZN => n21569);
   U19470 : INV_X1 port map( A => n16890, ZN => n21570);
   U19471 : INV_X1 port map( A => n16890, ZN => n21571);
   U19472 : INV_X1 port map( A => n16890, ZN => n21572);
   U19473 : INV_X1 port map( A => n16890, ZN => n21573);
   U19474 : INV_X1 port map( A => n21570, ZN => n21574);
   U19475 : INV_X1 port map( A => n21570, ZN => n21575);
   U19476 : INV_X1 port map( A => n21571, ZN => n21576);
   U19477 : INV_X1 port map( A => n21571, ZN => n21577);
   U19478 : INV_X1 port map( A => n21572, ZN => n21578);
   U19479 : INV_X1 port map( A => n21572, ZN => n21579);
   U19480 : INV_X1 port map( A => n21570, ZN => n21580);
   U19481 : INV_X1 port map( A => n21573, ZN => n21581);
   U19482 : INV_X1 port map( A => n21573, ZN => n21582);
   U19483 : INV_X1 port map( A => n21595, ZN => n21596);
   U19484 : INV_X1 port map( A => n21595, ZN => n21597);
   U19485 : INV_X1 port map( A => n21595, ZN => n21598);
   U19486 : INV_X1 port map( A => n21595, ZN => n21599);
   U19487 : INV_X1 port map( A => n21595, ZN => n21600);
   U19488 : INV_X1 port map( A => n21596, ZN => n21601);
   U19489 : INV_X1 port map( A => n21596, ZN => n21602);
   U19490 : INV_X1 port map( A => n21597, ZN => n21603);
   U19491 : INV_X1 port map( A => n21597, ZN => n21604);
   U19492 : INV_X1 port map( A => n21597, ZN => n21605);
   U19493 : INV_X1 port map( A => n21598, ZN => n21606);
   U19494 : INV_X1 port map( A => n21598, ZN => n21607);
   U19495 : INV_X1 port map( A => n21598, ZN => n21608);
   U19496 : INV_X1 port map( A => n21599, ZN => n21609);
   U19497 : INV_X1 port map( A => n21599, ZN => n21610);
   U19498 : INV_X1 port map( A => n21599, ZN => n21611);
   U19499 : INV_X1 port map( A => n21600, ZN => n21612);
   U19500 : INV_X1 port map( A => n21600, ZN => n21613);
   U19501 : INV_X1 port map( A => n21600, ZN => n21614);
   U19502 : INV_X1 port map( A => n16884, ZN => n21615);
   U19503 : INV_X1 port map( A => n16884, ZN => n21616);
   U19504 : INV_X1 port map( A => n16884, ZN => n21617);
   U19505 : INV_X1 port map( A => n16884, ZN => n21618);
   U19506 : INV_X1 port map( A => n21615, ZN => n21619);
   U19507 : INV_X1 port map( A => n21615, ZN => n21620);
   U19508 : INV_X1 port map( A => n21615, ZN => n21621);
   U19509 : INV_X1 port map( A => n21616, ZN => n21622);
   U19510 : INV_X1 port map( A => n21616, ZN => n21623);
   U19511 : INV_X1 port map( A => n21617, ZN => n21624);
   U19512 : INV_X1 port map( A => n21617, ZN => n21625);
   U19513 : INV_X1 port map( A => n21618, ZN => n21626);
   U19514 : INV_X1 port map( A => n21618, ZN => n21627);
   U19515 : INV_X1 port map( A => n21628, ZN => n21629);
   U19516 : INV_X1 port map( A => n21628, ZN => n21630);
   U19517 : INV_X1 port map( A => n21628, ZN => n21631);
   U19518 : INV_X1 port map( A => n21628, ZN => n21632);
   U19519 : INV_X1 port map( A => n21628, ZN => n21633);
   U19520 : INV_X1 port map( A => n21629, ZN => n21634);
   U19521 : INV_X1 port map( A => n21629, ZN => n21635);
   U19522 : INV_X1 port map( A => n21629, ZN => n21636);
   U19523 : INV_X1 port map( A => n21630, ZN => n21637);
   U19524 : INV_X1 port map( A => n21630, ZN => n21638);
   U19525 : INV_X1 port map( A => n21630, ZN => n21639);
   U19526 : INV_X1 port map( A => n21631, ZN => n21640);
   U19527 : INV_X1 port map( A => n21631, ZN => n21641);
   U19528 : INV_X1 port map( A => n21631, ZN => n21642);
   U19529 : INV_X1 port map( A => n21632, ZN => n21643);
   U19530 : INV_X1 port map( A => n21632, ZN => n21644);
   U19531 : INV_X1 port map( A => n21632, ZN => n21645);
   U19532 : INV_X1 port map( A => n21633, ZN => n21646);
   U19533 : INV_X1 port map( A => n21633, ZN => n21647);
   U19534 : INV_X1 port map( A => n21633, ZN => n21648);
   U19535 : INV_X1 port map( A => n21651, ZN => n21649);
   U19536 : INV_X1 port map( A => n16885, ZN => n21650);
   U19537 : INV_X1 port map( A => n16885, ZN => n21651);
   U19538 : INV_X1 port map( A => n16885, ZN => n21652);
   U19539 : INV_X1 port map( A => n21652, ZN => n21653);
   U19540 : INV_X1 port map( A => n21650, ZN => n21654);
   U19541 : INV_X1 port map( A => n21650, ZN => n21655);
   U19542 : INV_X1 port map( A => n21650, ZN => n21656);
   U19543 : INV_X1 port map( A => n21651, ZN => n21657);
   U19544 : INV_X1 port map( A => n21651, ZN => n21658);
   U19545 : INV_X1 port map( A => n21652, ZN => n21659);
   U19546 : INV_X1 port map( A => n21652, ZN => n21660);
   U19547 : INV_X1 port map( A => n16848, ZN => n21667);
   U19548 : INV_X1 port map( A => n16848, ZN => n21668);
   U19549 : INV_X1 port map( A => n21667, ZN => n21669);
   U19550 : INV_X1 port map( A => n21668, ZN => n21670);
   U19551 : INV_X1 port map( A => n21668, ZN => n21671);
   U19552 : INV_X1 port map( A => n21667, ZN => n21672);
   U19553 : INV_X1 port map( A => n21667, ZN => n21673);
   U19554 : INV_X1 port map( A => n21668, ZN => n21674);
   U19555 : INV_X1 port map( A => n16849, ZN => n21675);
   U19556 : INV_X1 port map( A => n16849, ZN => n21676);
   U19557 : INV_X1 port map( A => n21675, ZN => n21677);
   U19558 : INV_X1 port map( A => n21675, ZN => n21678);
   U19559 : INV_X1 port map( A => n21676, ZN => n21679);
   U19560 : INV_X1 port map( A => n21676, ZN => n21680);
   U19561 : INV_X1 port map( A => n21675, ZN => n21681);
   U19562 : INV_X1 port map( A => n21676, ZN => n21682);
   U19563 : INV_X1 port map( A => n21683, ZN => n21684);
   U19564 : INV_X1 port map( A => n21683, ZN => n21685);
   U19565 : INV_X1 port map( A => n21683, ZN => n21686);
   U19566 : INV_X1 port map( A => n21683, ZN => n21687);
   U19567 : INV_X1 port map( A => n21683, ZN => n21688);
   U19568 : INV_X1 port map( A => n21683, ZN => n21689);
   U19569 : INV_X1 port map( A => n21683, ZN => n21690);
   U19570 : INV_X1 port map( A => n21691, ZN => n21692);
   U19571 : INV_X1 port map( A => n21691, ZN => n21693);
   U19572 : INV_X1 port map( A => n21691, ZN => n21694);
   U19573 : INV_X1 port map( A => n21691, ZN => n21695);
   U19574 : INV_X1 port map( A => n21691, ZN => n21696);
   U19575 : INV_X1 port map( A => n21691, ZN => n21697);
   U19576 : INV_X1 port map( A => n21691, ZN => n21698);
   U19577 : INV_X1 port map( A => n16842, ZN => n21699);
   U19578 : INV_X1 port map( A => n16842, ZN => n21700);
   U19579 : INV_X1 port map( A => n21699, ZN => n21701);
   U19580 : INV_X1 port map( A => n21699, ZN => n21702);
   U19581 : INV_X1 port map( A => n21700, ZN => n21703);
   U19582 : INV_X1 port map( A => n21699, ZN => n21704);
   U19583 : INV_X1 port map( A => n21699, ZN => n21705);
   U19584 : INV_X1 port map( A => n21700, ZN => n21706);
   U19585 : INV_X1 port map( A => n21700, ZN => n21707);
   U19586 : INV_X1 port map( A => n16843, ZN => n21708);
   U19587 : INV_X1 port map( A => n16843, ZN => n21709);
   U19588 : INV_X1 port map( A => n21708, ZN => n21710);
   U19589 : INV_X1 port map( A => n21709, ZN => n21711);
   U19590 : INV_X1 port map( A => n21708, ZN => n21712);
   U19591 : INV_X1 port map( A => n21709, ZN => n21713);
   U19592 : INV_X1 port map( A => n21709, ZN => n21714);
   U19593 : INV_X1 port map( A => n21708, ZN => n21715);
   U19594 : INV_X1 port map( A => n21717, ZN => n21718);
   U19595 : INV_X1 port map( A => n21716, ZN => n21719);
   U19596 : INV_X1 port map( A => n21716, ZN => n21720);
   U19597 : INV_X1 port map( A => n21716, ZN => n21721);
   U19598 : INV_X1 port map( A => n21717, ZN => n21722);
   U19599 : INV_X1 port map( A => n21717, ZN => n21723);
   U19600 : INV_X1 port map( A => n21716, ZN => n21724);
   U19601 : INV_X1 port map( A => n21725, ZN => n21726);
   U19602 : INV_X1 port map( A => n21725, ZN => n21727);
   U19603 : INV_X1 port map( A => n21725, ZN => n21728);
   U19604 : INV_X1 port map( A => n21725, ZN => n21729);
   U19605 : INV_X1 port map( A => n21725, ZN => n21730);
   U19606 : INV_X1 port map( A => n21725, ZN => n21731);
   U19607 : INV_X1 port map( A => n21725, ZN => n21732);
   U19608 : INV_X1 port map( A => n21733, ZN => n21734);
   U19609 : INV_X1 port map( A => n21733, ZN => n21735);
   U19610 : INV_X1 port map( A => n21733, ZN => n21736);
   U19611 : INV_X1 port map( A => n21733, ZN => n21737);
   U19612 : INV_X1 port map( A => n21733, ZN => n21738);
   U19613 : INV_X1 port map( A => n21733, ZN => n21739);
   U19614 : INV_X1 port map( A => n21733, ZN => n21740);
   U19615 : INV_X1 port map( A => n21742, ZN => n21743);
   U19616 : INV_X1 port map( A => n21741, ZN => n21744);
   U19617 : INV_X1 port map( A => n21741, ZN => n21745);
   U19618 : INV_X1 port map( A => n21742, ZN => n21746);
   U19619 : INV_X1 port map( A => n21742, ZN => n21747);
   U19620 : INV_X1 port map( A => n21742, ZN => n21748);
   U19621 : INV_X1 port map( A => n21741, ZN => n21749);
   U19622 : INV_X1 port map( A => n21750, ZN => n21751);
   U19623 : INV_X1 port map( A => n21750, ZN => n21752);
   U19624 : INV_X1 port map( A => n21750, ZN => n21753);
   U19625 : INV_X1 port map( A => n21750, ZN => n21754);
   U19626 : INV_X1 port map( A => n21750, ZN => n21755);
   U19627 : INV_X1 port map( A => n21750, ZN => n21756);
   U19628 : INV_X1 port map( A => n21750, ZN => n21757);
   U19629 : INV_X1 port map( A => n16854, ZN => n21758);
   U19630 : INV_X1 port map( A => n16854, ZN => n21759);
   U19631 : INV_X1 port map( A => n21758, ZN => n21760);
   U19632 : INV_X1 port map( A => n21758, ZN => n21761);
   U19633 : INV_X1 port map( A => n21758, ZN => n21762);
   U19634 : INV_X1 port map( A => n21759, ZN => n21763);
   U19635 : INV_X1 port map( A => n21759, ZN => n21764);
   U19636 : INV_X1 port map( A => n21759, ZN => n21765);
   U19637 : INV_X1 port map( A => n16859, ZN => n21769);
   U19638 : INV_X1 port map( A => n21769, ZN => n21770);
   U19639 : INV_X1 port map( A => n21769, ZN => n21771);
   U19640 : INV_X1 port map( A => n21769, ZN => n21772);
   U19641 : INV_X1 port map( A => n21769, ZN => n21773);
   U19642 : INV_X1 port map( A => n21769, ZN => n21774);
   U19643 : INV_X1 port map( A => n21769, ZN => n21775);
   U19644 : INV_X1 port map( A => n21769, ZN => n21776);
   U19645 : INV_X1 port map( A => n16860, ZN => n21777);
   U19646 : INV_X1 port map( A => n21777, ZN => n21778);
   U19647 : INV_X1 port map( A => n21777, ZN => n21779);
   U19648 : INV_X1 port map( A => n21777, ZN => n21780);
   U19649 : INV_X1 port map( A => n21777, ZN => n21781);
   U19650 : INV_X1 port map( A => n21777, ZN => n21782);
   U19651 : INV_X1 port map( A => n21777, ZN => n21783);
   U19652 : INV_X1 port map( A => n21777, ZN => n21784);
   U19653 : INV_X1 port map( A => n21785, ZN => n21786);
   U19654 : INV_X1 port map( A => n21785, ZN => n21787);
   U19655 : INV_X1 port map( A => n21785, ZN => n21788);
   U19656 : INV_X1 port map( A => n21785, ZN => n21789);
   U19657 : INV_X1 port map( A => n21785, ZN => n21790);
   U19658 : INV_X1 port map( A => n21785, ZN => n21791);
   U19659 : INV_X1 port map( A => n21785, ZN => n21792);
   U19660 : INV_X1 port map( A => n21793, ZN => n21794);
   U19661 : INV_X1 port map( A => n21793, ZN => n21795);
   U19662 : INV_X1 port map( A => n21793, ZN => n21796);
   U19663 : INV_X1 port map( A => n21793, ZN => n21797);
   U19664 : INV_X1 port map( A => n21793, ZN => n21798);
   U19665 : INV_X1 port map( A => n21793, ZN => n21799);
   U19666 : INV_X1 port map( A => n21793, ZN => n21800);
   U19667 : CLKBUF_X1 port map( A => n15153, Z => n22370);
   U19668 : CLKBUF_X1 port map( A => n15153, Z => n22371);
   U19669 : CLKBUF_X1 port map( A => n15153, Z => n22372);
   U19670 : CLKBUF_X1 port map( A => n15150, Z => n22386);
   U19671 : CLKBUF_X1 port map( A => n15149, Z => n22392);
   U19672 : CLKBUF_X1 port map( A => n15148, Z => n22398);
   U19673 : CLKBUF_X1 port map( A => n15147, Z => n22404);
   U19674 : CLKBUF_X1 port map( A => n15146, Z => n22410);
   U19675 : CLKBUF_X1 port map( A => n15145, Z => n22416);
   U19676 : CLKBUF_X1 port map( A => n15144, Z => n22422);
   U19677 : CLKBUF_X1 port map( A => n15143, Z => n22428);
   U19678 : CLKBUF_X1 port map( A => n15142, Z => n22434);
   U19679 : CLKBUF_X1 port map( A => n15141, Z => n22440);
   U19680 : CLKBUF_X1 port map( A => n15140, Z => n22446);
   U19681 : CLKBUF_X1 port map( A => n15139, Z => n22452);
   U19682 : CLKBUF_X1 port map( A => n15138, Z => n22458);
   U19683 : CLKBUF_X1 port map( A => n15137, Z => n22464);
   U19684 : CLKBUF_X1 port map( A => n15136, Z => n22470);
   U19685 : CLKBUF_X1 port map( A => n15135, Z => n22476);
   U19686 : CLKBUF_X1 port map( A => n15134, Z => n22482);
   U19687 : CLKBUF_X1 port map( A => n15133, Z => n22488);
   U19688 : CLKBUF_X1 port map( A => n15132, Z => n22494);
   U19689 : CLKBUF_X1 port map( A => n15131, Z => n22500);
   U19690 : CLKBUF_X1 port map( A => n15130, Z => n22506);
   U19691 : CLKBUF_X1 port map( A => n15129, Z => n22512);
   U19692 : CLKBUF_X1 port map( A => n15128, Z => n22518);
   U19693 : CLKBUF_X1 port map( A => n15127, Z => n22524);
   U19694 : CLKBUF_X1 port map( A => n15126, Z => n22530);
   U19695 : CLKBUF_X1 port map( A => n15125, Z => n22536);
   U19696 : CLKBUF_X1 port map( A => n15124, Z => n22542);
   U19697 : CLKBUF_X1 port map( A => n15123, Z => n22548);
   U19698 : CLKBUF_X1 port map( A => n15122, Z => n22554);
   U19699 : CLKBUF_X1 port map( A => n15121, Z => n22560);
   U19700 : CLKBUF_X1 port map( A => n15120, Z => n22566);
   U19701 : CLKBUF_X1 port map( A => n15118, Z => n22581);

end SYN_BEHAVIORAL;
