
module FA_1071 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1070 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1069 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1068 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1067 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1066 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1065 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1064 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1063 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1062 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1061 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1060 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1059 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Co) );
endmodule


module FA_1058 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1057 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1056 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1055 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1054 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1053 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1052 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1051 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1050 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1049 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1048 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1047 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1046 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1045 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1044 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1043 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Co) );
endmodule


module FA_1042 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1041 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1040 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1039 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1038 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1037 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1036 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1035 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  AOI22_X1 U1 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
  INV_X1 U2 ( .A(n4), .ZN(Co) );
endmodule


module FA_1034 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1033 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1032 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1031 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1030 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1029 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1028 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1027 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1026 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1025 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1024 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1023 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1022 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1021 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1020 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1019 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1018 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1017 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1016 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1015 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1014 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1013 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1012 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1011 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1010 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1009 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module MUX21_GENERIC_N4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(n2), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n3), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n1), .ZN(Y[0]) );
  INV_X1 U4 ( .A(n5), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[3]), .A2(n4), .B1(SEL), .B2(B[3]), .ZN(n5) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n4), .B1(B[2]), .B2(SEL), .ZN(n3) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(SEL), .ZN(n2) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(SEL), .ZN(n1) );
  INV_X1 U9 ( .A(SEL), .ZN(n4) );
endmodule


module MUX21_GENERIC_N4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(n2), .ZN(Y[1]) );
  INV_X1 U2 ( .A(n3), .ZN(Y[2]) );
  INV_X1 U3 ( .A(n1), .ZN(Y[0]) );
  INV_X1 U4 ( .A(n5), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(A[3]), .A2(n4), .B1(SEL), .B2(B[3]), .ZN(n5) );
  AOI22_X1 U6 ( .A1(A[2]), .A2(n4), .B1(B[2]), .B2(SEL), .ZN(n3) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(SEL), .ZN(n2) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(SEL), .ZN(n1) );
  INV_X1 U9 ( .A(SEL), .ZN(n4) );
endmodule


module MUX21_GENERIC_N4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n1, n2, n3, n4, n5;

  INV_X1 U1 ( .A(SEL), .ZN(n4) );
  INV_X1 U2 ( .A(n2), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(A[1]), .A2(n4), .B1(B[1]), .B2(SEL), .ZN(n2) );
  INV_X1 U4 ( .A(n3), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(n4), .B1(B[2]), .B2(SEL), .ZN(n3) );
  INV_X1 U6 ( .A(n1), .ZN(Y[0]) );
  AOI22_X1 U7 ( .A1(A[0]), .A2(n4), .B1(B[0]), .B2(SEL), .ZN(n1) );
  INV_X1 U8 ( .A(n5), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n4), .B1(SEL), .B2(B[3]), .ZN(n5) );
endmodule


module MUX21_GENERIC_N4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   net167137, n1, n2;

  MUX2_X1 syn42 ( .A(A[3]), .B(B[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 syn40 ( .A(A[2]), .B(B[2]), .S(SEL), .Z(Y[2]) );
  INV_X1 U1 ( .A(SEL), .ZN(net167137) );
  INV_X1 U2 ( .A(n2), .ZN(Y[1]) );
  INV_X1 U3 ( .A(n1), .ZN(Y[0]) );
  AOI22_X1 U4 ( .A1(net167137), .A2(A[0]), .B1(SEL), .B2(B[0]), .ZN(n1) );
  AOI22_X1 U5 ( .A1(net167137), .A2(A[1]), .B1(SEL), .B2(B[1]), .ZN(n2) );
endmodule


module MUX21_GENERIC_N4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX2_X1 syn61 ( .A(A[3]), .B(B[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 syn57 ( .A(A[2]), .B(B[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U1 ( .A(A[0]), .B(B[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(A[1]), .B(B[1]), .S(SEL), .Z(Y[1]) );
endmodule


module MUX21_GENERIC_N4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX2_X1 syn61 ( .A(A[3]), .B(B[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 syn57 ( .A(A[2]), .B(B[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U1 ( .A(A[0]), .B(B[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(A[1]), .B(B[1]), .S(SEL), .Z(Y[1]) );
endmodule


module MUX21_GENERIC_N4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX2_X1 syn61 ( .A(A[3]), .B(B[3]), .S(SEL), .Z(Y[3]) );
  MUX2_X1 syn57 ( .A(A[2]), .B(B[2]), .S(SEL), .Z(Y[2]) );
  MUX2_X1 U1 ( .A(A[0]), .B(B[0]), .S(SEL), .Z(Y[0]) );
  MUX2_X1 U2 ( .A(A[1]), .B(B[1]), .S(SEL), .Z(Y[1]) );
endmodule


module RCA_generic_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1068 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1067 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1066 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1065 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1064 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1063 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1062 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1061 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1060 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1059 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1058 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1057 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1056 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1055 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1054 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1053 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1052 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1051 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1050 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1049 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1048 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1047 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1046 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1045 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1044 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1043 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1042 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1041 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1040 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1039 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1038 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1037 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1036 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1035 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1034 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1033 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1032 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1031 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1030 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1029 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1028 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1027 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1026 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1025 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1024 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1023 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1022 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1021 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1020 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1019 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1018 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1017 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1016 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1015 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1014 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1013 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_generic_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1012 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1011 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1010 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1009 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CARRY_SELECT_BLOCK_N4_7 ( A, B, C_in, O, C_o );
  input [3:0] A;
  input [3:0] B;
  output [3:0] O;
  input C_in;
  output C_o;

  wire   [3:0] mux_A;
  wire   [3:0] mux_B;

  RCA_generic_N4_14 carry_in_0 ( .A(A), .B(B), .Ci(1'b0), .S(mux_A) );
  RCA_generic_N4_13 carry_in_1 ( .A(A), .B(B), .Ci(1'b1), .S(mux_B) );
  MUX21_GENERIC_N4_7 mux_sum ( .A(mux_A), .B(mux_B), .SEL(C_in), .Y(O) );
endmodule


module CARRY_SELECT_BLOCK_N4_6 ( A, B, C_in, O, C_o );
  input [3:0] A;
  input [3:0] B;
  output [3:0] O;
  input C_in;
  output C_o;

  wire   [3:0] mux_A;
  wire   [3:0] mux_B;

  RCA_generic_N4_12 carry_in_0 ( .A(A), .B(B), .Ci(1'b0), .S(mux_A) );
  RCA_generic_N4_11 carry_in_1 ( .A(A), .B(B), .Ci(1'b1), .S(mux_B) );
  MUX21_GENERIC_N4_6 mux_sum ( .A(mux_A), .B(mux_B), .SEL(C_in), .Y(O) );
endmodule


module CARRY_SELECT_BLOCK_N4_5 ( A, B, C_in, O, C_o );
  input [3:0] A;
  input [3:0] B;
  output [3:0] O;
  input C_in;
  output C_o;

  wire   [3:0] mux_A;
  wire   [3:0] mux_B;

  RCA_generic_N4_10 carry_in_0 ( .A(A), .B(B), .Ci(1'b0), .S(mux_A) );
  RCA_generic_N4_9 carry_in_1 ( .A(A), .B(B), .Ci(1'b1), .S(mux_B) );
  MUX21_GENERIC_N4_5 mux_sum ( .A(mux_A), .B(mux_B), .SEL(C_in), .Y(O) );
endmodule


module CARRY_SELECT_BLOCK_N4_4 ( A, B, C_in, O, C_o );
  input [3:0] A;
  input [3:0] B;
  output [3:0] O;
  input C_in;
  output C_o;

  wire   [3:0] mux_A;
  wire   [3:0] mux_B;

  RCA_generic_N4_8 carry_in_0 ( .A(A), .B(B), .Ci(1'b0), .S(mux_A) );
  RCA_generic_N4_7 carry_in_1 ( .A(A), .B(B), .Ci(1'b1), .S(mux_B) );
  MUX21_GENERIC_N4_4 mux_sum ( .A(mux_A), .B(mux_B), .SEL(C_in), .Y(O) );
endmodule


module CARRY_SELECT_BLOCK_N4_3 ( A, B, C_in, O, C_o );
  input [3:0] A;
  input [3:0] B;
  output [3:0] O;
  input C_in;
  output C_o;

  wire   [3:0] mux_A;
  wire   [3:0] mux_B;

  RCA_generic_N4_6 carry_in_0 ( .A(A), .B(B), .Ci(1'b0), .S(mux_A) );
  RCA_generic_N4_5 carry_in_1 ( .A(A), .B(B), .Ci(1'b1), .S(mux_B) );
  MUX21_GENERIC_N4_3 mux_sum ( .A(mux_A), .B(mux_B), .SEL(C_in), .Y(O) );
endmodule


module CARRY_SELECT_BLOCK_N4_2 ( A, B, C_in, O, C_o );
  input [3:0] A;
  input [3:0] B;
  output [3:0] O;
  input C_in;
  output C_o;

  wire   [3:0] mux_A;
  wire   [3:0] mux_B;

  RCA_generic_N4_4 carry_in_0 ( .A(A), .B(B), .Ci(1'b0), .S(mux_A) );
  RCA_generic_N4_3 carry_in_1 ( .A(A), .B(B), .Ci(1'b1), .S(mux_B) );
  MUX21_GENERIC_N4_2 mux_sum ( .A(mux_A), .B(mux_B), .SEL(C_in), .Y(O) );
endmodule


module CARRY_SELECT_BLOCK_N4_1 ( A, B, C_in, O, C_o );
  input [3:0] A;
  input [3:0] B;
  output [3:0] O;
  input C_in;
  output C_o;

  wire   [3:0] mux_A;
  wire   [3:0] mux_B;

  RCA_generic_N4_2 carry_in_0 ( .A(A), .B(B), .Ci(1'b0), .S(mux_A) );
  RCA_generic_N4_1 carry_in_1 ( .A(A), .B(B), .Ci(1'b1), .S(mux_B) );
  MUX21_GENERIC_N4_1 mux_sum ( .A(mux_A), .B(mux_B), .SEL(C_in), .Y(O) );
endmodule


module PG_BLOCK_26 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AND2_X1 U2 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  AOI21_X1 U3 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
endmodule


module PG_BLOCK_25 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AOI21_X1 U2 ( .B1(Pi[1]), .B2(Gi[0]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
endmodule


module PG_BLOCK_24 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Go) );
  AND2_X1 U3 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
endmodule


module PG_BLOCK_23 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  AOI21_X1 U2 ( .B1(Pi[1]), .B2(Gi[0]), .A(Gi[1]), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Go) );
endmodule


module PG_BLOCK_22 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U2 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  INV_X1 U3 ( .A(n3), .ZN(Go) );
endmodule


module PG_BLOCK_21 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AOI21_X1 U2 ( .B1(Pi[1]), .B2(Gi[0]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
endmodule


module PG_BLOCK_20 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U2 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  INV_X1 U3 ( .A(n3), .ZN(Go) );
endmodule


module PG_BLOCK_19 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U2 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  INV_X1 U3 ( .A(n3), .ZN(Go) );
endmodule


module PG_BLOCK_18 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
endmodule


module PG_BLOCK_17 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  INV_X1 U2 ( .A(n3), .ZN(Go) );
  AOI21_X1 U3 ( .B1(Pi[1]), .B2(Gi[0]), .A(Gi[1]), .ZN(n3) );
endmodule


module PG_BLOCK_16 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
endmodule


module PG_BLOCK_15 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
endmodule


module PG_BLOCK_14 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
endmodule


module PG_BLOCK_13 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
endmodule


module PG_BLOCK_12 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Go) );
endmodule


module PG_BLOCK_11 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Go) );
endmodule


module PG_BLOCK_10 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Go) );
endmodule


module PG_BLOCK_9 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  INV_X1 U2 ( .A(n3), .ZN(Go) );
  AOI21_X1 U3 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
endmodule


module PG_BLOCK_8 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Go) );
endmodule


module PG_BLOCK_7 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  AND2_X1 U3 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
endmodule


module PG_BLOCK_6 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AOI21_X1 U1 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Go) );
  AND2_X1 U3 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
endmodule


module PG_BLOCK_5 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3, n4;

  INV_X1 U1 ( .A(Gi[1]), .ZN(n3) );
  AND2_X1 U2 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  NAND2_X1 U3 ( .A1(Gi[0]), .A2(Pi[1]), .ZN(n4) );
  NAND2_X1 U4 ( .A1(n3), .A2(n4), .ZN(Go) );
endmodule


module PG_BLOCK_4 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Go) );
endmodule


module PG_BLOCK_3 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  INV_X1 U2 ( .A(n3), .ZN(Go) );
  AOI21_X1 U3 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
endmodule


module PG_BLOCK_2 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  AOI21_X1 U2 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
  INV_X1 U3 ( .A(n3), .ZN(Go) );
endmodule


module PG_BLOCK_1 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n3;

  AND2_X1 U1 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  INV_X1 U2 ( .A(n3), .ZN(Go) );
  AOI21_X1 U3 ( .B1(Gi[0]), .B2(Pi[1]), .A(Gi[1]), .ZN(n3) );
endmodule


module G_BLOCK_8 ( Gi, Pi, Go );
  input [1:0] Gi;
  input Pi;
  output Go;
  wire   n3;

  AOI21_X1 U1 ( .B1(Pi), .B2(Gi[0]), .A(Gi[1]), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(Go) );
endmodule


module G_BLOCK_7 ( Gi, Pi, Go );
  input [1:0] Gi;
  input Pi;
  output Go;
  wire   n2, n3;

  INV_X1 U1 ( .A(Gi[1]), .ZN(n2) );
  NAND2_X1 U2 ( .A1(n3), .A2(n2), .ZN(Go) );
  NAND2_X1 U3 ( .A1(Gi[0]), .A2(Pi), .ZN(n3) );
endmodule


module G_BLOCK_6 ( Gi, Pi, Go );
  input [1:0] Gi;
  input Pi;
  output Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AOI21_X1 U2 ( .B1(Pi), .B2(Gi[0]), .A(Gi[1]), .ZN(n3) );
endmodule


module G_BLOCK_5 ( Gi, Pi, Go );
  input [1:0] Gi;
  input Pi;
  output Go;
  wire   n2, n3;

  NAND2_X1 U1 ( .A1(n3), .A2(n2), .ZN(Go) );
  INV_X1 U2 ( .A(Gi[1]), .ZN(n2) );
  NAND2_X1 U3 ( .A1(Gi[0]), .A2(Pi), .ZN(n3) );
endmodule


module G_BLOCK_4 ( Gi, Pi, Go );
  input [1:0] Gi;
  input Pi;
  output Go;
  wire   n2, n3;

  INV_X1 U1 ( .A(Gi[1]), .ZN(n2) );
  NAND2_X1 U2 ( .A1(Gi[0]), .A2(Pi), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n3), .A2(n2), .ZN(Go) );
endmodule


module G_BLOCK_3 ( Gi, Pi, Go );
  input [1:0] Gi;
  input Pi;
  output Go;
  wire   n2, n3;

  INV_X1 U1 ( .A(Gi[1]), .ZN(n2) );
  NAND2_X1 U2 ( .A1(n3), .A2(n2), .ZN(Go) );
  NAND2_X1 U3 ( .A1(Gi[0]), .A2(Pi), .ZN(n3) );
endmodule


module G_BLOCK_2 ( Gi, Pi, Go );
  input [1:0] Gi;
  input Pi;
  output Go;
  wire   n2, n3;

  NAND2_X1 U1 ( .A1(n3), .A2(n2), .ZN(Go) );
  INV_X1 U2 ( .A(Gi[1]), .ZN(n2) );
  NAND2_X1 U3 ( .A1(Gi[0]), .A2(Pi), .ZN(n3) );
endmodule


module G_BLOCK_1 ( Gi, Pi, Go );
  input [1:0] Gi;
  input Pi;
  output Go;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(Go) );
  AOI21_X1 U2 ( .B1(Pi), .B2(Gi[0]), .A(Gi[1]), .ZN(n3) );
endmodule


module FA_1008 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_GENERIC_N4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n10;

  INV_X1 U1 ( .A(SEL), .ZN(n7) );
  INV_X1 U2 ( .A(n9), .ZN(Y[1]) );
  AOI22_X1 U3 ( .A1(A[1]), .A2(n7), .B1(B[1]), .B2(SEL), .ZN(n9) );
  INV_X1 U4 ( .A(n8), .ZN(Y[2]) );
  AOI22_X1 U5 ( .A1(A[2]), .A2(n7), .B1(B[2]), .B2(SEL), .ZN(n8) );
  INV_X1 U6 ( .A(n10), .ZN(Y[0]) );
  AOI22_X1 U7 ( .A1(A[0]), .A2(n7), .B1(B[0]), .B2(SEL), .ZN(n10) );
  INV_X1 U8 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U9 ( .A1(A[3]), .A2(n7), .B1(SEL), .B2(B[3]), .ZN(n6) );
endmodule


module RCA_generic_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_1008 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_1071 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_1070 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1069 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CARRY_SELECT_BLOCK_N4_0 ( A, B, C_in, O, C_o );
  input [3:0] A;
  input [3:0] B;
  output [3:0] O;
  input C_in;
  output C_o;

  wire   [3:0] mux_A;
  wire   [3:0] mux_B;

  RCA_generic_N4_0 carry_in_0 ( .A(A), .B(B), .Ci(1'b0), .S(mux_A) );
  RCA_generic_N4_15 carry_in_1 ( .A(A), .B(B), .Ci(1'b1), .S(mux_B) );
  MUX21_GENERIC_N4_0 mux_sum ( .A(mux_A), .B(mux_B), .SEL(C_in), .Y(O) );
endmodule


module PG_BLOCK_0 ( Gi, Pi, Po, Go );
  input [1:0] Gi;
  input [1:0] Pi;
  output Po, Go;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(Go) );
  AND2_X1 U2 ( .A1(Pi[1]), .A2(Pi[0]), .ZN(Po) );
  AOI21_X1 U3 ( .B1(Pi[1]), .B2(Gi[0]), .A(Gi[1]), .ZN(n2) );
endmodule


module G_BLOCK_0 ( Gi, Pi, Go );
  input [1:0] Gi;
  input Pi;
  output Go;
  wire   n2;

  AOI21_X1 U1 ( .B1(Pi), .B2(Gi[0]), .A(Gi[1]), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(Go) );
endmodule


module SUM_GENERATOR_N32 ( A, B, C_in, O, C_o );
  input [31:0] A;
  input [31:0] B;
  input [8:0] C_in;
  output [31:0] O;
  output C_o;

  assign C_o = C_in[8];

  CARRY_SELECT_BLOCK_N4_0 csa_block_0 ( .A(A[3:0]), .B(B[3:0]), .C_in(C_in[0]), 
        .O(O[3:0]) );
  CARRY_SELECT_BLOCK_N4_7 csa_block_1 ( .A(A[7:4]), .B(B[7:4]), .C_in(C_in[1]), 
        .O(O[7:4]) );
  CARRY_SELECT_BLOCK_N4_6 csa_block_2 ( .A(A[11:8]), .B(B[11:8]), .C_in(
        C_in[2]), .O(O[11:8]) );
  CARRY_SELECT_BLOCK_N4_5 csa_block_3 ( .A(A[15:12]), .B(B[15:12]), .C_in(
        C_in[3]), .O(O[15:12]) );
  CARRY_SELECT_BLOCK_N4_4 csa_block_4 ( .A(A[19:16]), .B(B[19:16]), .C_in(
        C_in[4]), .O(O[19:16]) );
  CARRY_SELECT_BLOCK_N4_3 csa_block_5 ( .A(A[23:20]), .B(B[23:20]), .C_in(
        C_in[5]), .O(O[23:20]) );
  CARRY_SELECT_BLOCK_N4_2 csa_block_6 ( .A(A[27:24]), .B(B[27:24]), .C_in(
        C_in[6]), .O(O[27:24]) );
  CARRY_SELECT_BLOCK_N4_1 csa_block_7 ( .A(A[31:28]), .B(B[31:28]), .C_in(
        C_in[7]), .O(O[31:28]) );
endmodule


module CARRY_GENERATOR_N32 ( A, B, C_in, C_o );
  input [31:0] A;
  input [31:0] B;
  output [8:0] C_o;
  input C_in;
  wire   C_in, n22, n23, n24, G_10, \GG[2][7] , \GG[2][6] , \GG[1][7] ,
         \GG[1][5] , \GG[1][3] , \GG[0][7] , \GG[0][6] , \GG[0][5] ,
         \GG[0][4] , \GG[0][3] , \GG[0][2] , \GG[0][1] , \PP[2][7] ,
         \PP[2][6] , \PP[1][7] , \PP[1][5] , \PP[1][3] , \PP[0][7] ,
         \PP[0][6] , \PP[0][5] , \PP[0][4] , \PP[0][3] , \PP[0][2] ,
         \PP[0][1] , n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n16,
         n17, n18, n19;
  wire   [32:1] p;
  wire   [32:1] g;
  wire   [15:0] first_g;
  wire   [15:1] first_p;
  assign C_o[0] = C_in;

  G_BLOCK_0 g_i_0 ( .Gi({g[2], G_10}), .Pi(p[2]), .Go(first_g[0]) );
  PG_BLOCK_0 pg_i_1 ( .Gi(g[4:3]), .Pi(p[4:3]), .Po(first_p[1]), .Go(
        first_g[1]) );
  PG_BLOCK_26 pg_i_2 ( .Gi(g[6:5]), .Pi(p[6:5]), .Po(first_p[2]), .Go(
        first_g[2]) );
  PG_BLOCK_25 pg_i_3 ( .Gi(g[8:7]), .Pi(p[8:7]), .Po(first_p[3]), .Go(
        first_g[3]) );
  PG_BLOCK_24 pg_i_4 ( .Gi(g[10:9]), .Pi(p[10:9]), .Po(first_p[4]), .Go(
        first_g[4]) );
  PG_BLOCK_23 pg_i_5 ( .Gi(g[12:11]), .Pi(p[12:11]), .Po(first_p[5]), .Go(
        first_g[5]) );
  PG_BLOCK_22 pg_i_6 ( .Gi(g[14:13]), .Pi(p[14:13]), .Po(first_p[6]), .Go(
        first_g[6]) );
  PG_BLOCK_21 pg_i_7 ( .Gi(g[16:15]), .Pi(p[16:15]), .Po(first_p[7]), .Go(
        first_g[7]) );
  PG_BLOCK_20 pg_i_8 ( .Gi(g[18:17]), .Pi(p[18:17]), .Po(first_p[8]), .Go(
        first_g[8]) );
  PG_BLOCK_19 pg_i_9 ( .Gi(g[20:19]), .Pi(p[20:19]), .Po(first_p[9]), .Go(
        first_g[9]) );
  PG_BLOCK_18 pg_i_10 ( .Gi(g[22:21]), .Pi(p[22:21]), .Po(first_p[10]), .Go(
        first_g[10]) );
  PG_BLOCK_17 pg_i_11 ( .Gi(g[24:23]), .Pi(p[24:23]), .Po(first_p[11]), .Go(
        first_g[11]) );
  PG_BLOCK_16 pg_i_12 ( .Gi(g[26:25]), .Pi(p[26:25]), .Po(first_p[12]), .Go(
        first_g[12]) );
  PG_BLOCK_15 pg_i_13 ( .Gi(g[28:27]), .Pi(p[28:27]), .Po(first_p[13]), .Go(
        first_g[13]) );
  PG_BLOCK_14 pg_i_14 ( .Gi(g[30:29]), .Pi(p[30:29]), .Po(first_p[14]), .Go(
        first_g[14]) );
  PG_BLOCK_13 pg_i_15 ( .Gi(g[32:31]), .Pi(p[32:31]), .Po(first_p[15]), .Go(
        first_g[15]) );
  G_BLOCK_8 g_i_0_0 ( .Gi(first_g[1:0]), .Pi(first_p[1]), .Go(n24) );
  PG_BLOCK_12 pg_i_1_0 ( .Gi(first_g[3:2]), .Pi(first_p[3:2]), .Po(\PP[0][1] ), 
        .Go(\GG[0][1] ) );
  PG_BLOCK_11 pg_i_2_0 ( .Gi(first_g[5:4]), .Pi(first_p[5:4]), .Po(\PP[0][2] ), 
        .Go(\GG[0][2] ) );
  PG_BLOCK_10 pg_i_3_0 ( .Gi(first_g[7:6]), .Pi(first_p[7:6]), .Po(\PP[0][3] ), 
        .Go(\GG[0][3] ) );
  PG_BLOCK_9 pg_i_4_0 ( .Gi(first_g[9:8]), .Pi(first_p[9:8]), .Po(\PP[0][4] ), 
        .Go(\GG[0][4] ) );
  PG_BLOCK_8 pg_i_5_0 ( .Gi(first_g[11:10]), .Pi(first_p[11:10]), .Po(
        \PP[0][5] ), .Go(\GG[0][5] ) );
  PG_BLOCK_7 pg_i_6_0 ( .Gi(first_g[13:12]), .Pi(first_p[13:12]), .Po(
        \PP[0][6] ), .Go(\GG[0][6] ) );
  PG_BLOCK_6 pg_i_7_0 ( .Gi(first_g[15:14]), .Pi(first_p[15:14]), .Po(
        \PP[0][7] ), .Go(\GG[0][7] ) );
  G_BLOCK_7 g_i_0_1 ( .Gi({\GG[0][1] , n24}), .Pi(\PP[0][1] ), .Go(n23) );
  PG_BLOCK_5 pg_i_0_3 ( .Gi({\GG[0][3] , \GG[0][2] }), .Pi({\PP[0][3] , 
        \PP[0][2] }), .Po(\PP[1][3] ), .Go(\GG[1][3] ) );
  PG_BLOCK_4 pg_i_0_5 ( .Gi({\GG[0][5] , \GG[0][4] }), .Pi({\PP[0][5] , 
        \PP[0][4] }), .Po(\PP[1][5] ), .Go(\GG[1][5] ) );
  PG_BLOCK_3 pg_i_0_7 ( .Gi({\GG[0][7] , \GG[0][6] }), .Pi({\PP[0][7] , 
        \PP[0][6] }), .Po(\PP[1][7] ), .Go(\GG[1][7] ) );
  G_BLOCK_6 g_i_1_2 ( .Gi({\GG[0][2] , n23}), .Pi(\PP[0][2] ), .Go(C_o[3]) );
  G_BLOCK_5 g_i_1_3 ( .Gi({\GG[1][3] , n23}), .Pi(\PP[1][3] ), .Go(n22) );
  PG_BLOCK_2 pg_i_1_6 ( .Gi({\GG[0][6] , \GG[1][5] }), .Pi({\PP[0][6] , 
        \PP[1][5] }), .Po(\PP[2][6] ), .Go(\GG[2][6] ) );
  PG_BLOCK_1 pg_i_1_7 ( .Gi({\GG[1][7] , n14}), .Pi({\PP[1][7] , \PP[1][5] }), 
        .Po(\PP[2][7] ), .Go(\GG[2][7] ) );
  G_BLOCK_4 g_i_2_4 ( .Gi({\GG[0][4] , n22}), .Pi(\PP[0][4] ), .Go(C_o[5]) );
  G_BLOCK_3 g_i_2_5 ( .Gi({n14, n22}), .Pi(\PP[1][5] ), .Go(C_o[6]) );
  G_BLOCK_2 g_i_2_6 ( .Gi({\GG[2][6] , n22}), .Pi(\PP[2][6] ), .Go(C_o[7]) );
  G_BLOCK_1 g_i_2_7 ( .Gi({\GG[2][7] , C_o[4]}), .Pi(\PP[2][7] ), .Go(C_o[8])
         );
  XOR2_X1 U36 ( .A(B[8]), .B(A[8]), .Z(p[9]) );
  XOR2_X1 U38 ( .A(B[6]), .B(A[6]), .Z(p[7]) );
  XOR2_X1 U39 ( .A(B[5]), .B(A[5]), .Z(p[6]) );
  XOR2_X1 U40 ( .A(B[4]), .B(A[4]), .Z(p[5]) );
  XOR2_X1 U41 ( .A(B[3]), .B(A[3]), .Z(p[4]) );
  XOR2_X1 U42 ( .A(B[2]), .B(A[2]), .Z(p[3]) );
  XOR2_X1 U43 ( .A(B[31]), .B(A[31]), .Z(p[32]) );
  XOR2_X1 U44 ( .A(B[30]), .B(A[30]), .Z(p[31]) );
  XOR2_X1 U45 ( .A(B[29]), .B(A[29]), .Z(p[30]) );
  XOR2_X1 U46 ( .A(B[1]), .B(A[1]), .Z(p[2]) );
  XOR2_X1 U47 ( .A(B[28]), .B(A[28]), .Z(p[29]) );
  XOR2_X1 U48 ( .A(B[27]), .B(A[27]), .Z(p[28]) );
  XOR2_X1 U49 ( .A(B[26]), .B(A[26]), .Z(p[27]) );
  XOR2_X1 U50 ( .A(B[25]), .B(A[25]), .Z(p[26]) );
  XOR2_X1 U51 ( .A(B[24]), .B(A[24]), .Z(p[25]) );
  XOR2_X1 U52 ( .A(B[23]), .B(A[23]), .Z(p[24]) );
  XOR2_X1 U53 ( .A(B[22]), .B(A[22]), .Z(p[23]) );
  XOR2_X1 U54 ( .A(B[21]), .B(A[21]), .Z(p[22]) );
  XOR2_X1 U55 ( .A(B[20]), .B(A[20]), .Z(p[21]) );
  XOR2_X1 U56 ( .A(B[19]), .B(A[19]), .Z(p[20]) );
  XOR2_X1 U57 ( .A(B[18]), .B(A[18]), .Z(p[19]) );
  XOR2_X1 U58 ( .A(B[17]), .B(A[17]), .Z(p[18]) );
  XOR2_X1 U59 ( .A(B[16]), .B(A[16]), .Z(p[17]) );
  XOR2_X1 U61 ( .A(B[14]), .B(A[14]), .Z(p[15]) );
  XOR2_X1 U62 ( .A(B[13]), .B(A[13]), .Z(p[14]) );
  XOR2_X1 U63 ( .A(B[12]), .B(A[12]), .Z(p[13]) );
  XOR2_X1 U65 ( .A(B[10]), .B(A[10]), .Z(p[11]) );
  XOR2_X1 U66 ( .A(B[9]), .B(A[9]), .Z(p[10]) );
  BUF_X1 U1 ( .A(n23), .Z(C_o[2]) );
  BUF_X2 U2 ( .A(n22), .Z(C_o[4]) );
  AND2_X1 U3 ( .A1(B[14]), .A2(A[14]), .ZN(g[15]) );
  AND2_X1 U4 ( .A1(B[18]), .A2(A[18]), .ZN(g[19]) );
  AND2_X1 U5 ( .A1(B[19]), .A2(A[19]), .ZN(g[20]) );
  AND2_X1 U6 ( .A1(B[22]), .A2(A[22]), .ZN(g[23]) );
  AND2_X1 U7 ( .A1(B[23]), .A2(A[23]), .ZN(g[24]) );
  AND2_X1 U8 ( .A1(B[12]), .A2(A[12]), .ZN(g[13]) );
  AND2_X1 U9 ( .A1(B[13]), .A2(A[13]), .ZN(g[14]) );
  AND2_X1 U10 ( .A1(B[10]), .A2(A[10]), .ZN(g[11]) );
  AND2_X1 U11 ( .A1(B[11]), .A2(A[11]), .ZN(g[12]) );
  AND2_X1 U12 ( .A1(B[8]), .A2(A[8]), .ZN(g[9]) );
  AND2_X1 U13 ( .A1(B[9]), .A2(A[9]), .ZN(g[10]) );
  AND2_X1 U14 ( .A1(B[6]), .A2(A[6]), .ZN(g[7]) );
  AND2_X1 U15 ( .A1(B[7]), .A2(A[7]), .ZN(g[8]) );
  AND2_X1 U16 ( .A1(B[26]), .A2(A[26]), .ZN(g[27]) );
  AND2_X1 U17 ( .A1(B[27]), .A2(A[27]), .ZN(g[28]) );
  AND2_X1 U18 ( .A1(B[24]), .A2(A[24]), .ZN(g[25]) );
  AND2_X1 U19 ( .A1(B[25]), .A2(A[25]), .ZN(g[26]) );
  AND2_X1 U20 ( .A1(B[30]), .A2(A[30]), .ZN(g[31]) );
  AND2_X1 U21 ( .A1(B[31]), .A2(A[31]), .ZN(g[32]) );
  AND2_X1 U22 ( .A1(B[1]), .A2(A[1]), .ZN(g[2]) );
  AND2_X1 U23 ( .A1(B[16]), .A2(A[16]), .ZN(g[17]) );
  AND2_X1 U24 ( .A1(B[17]), .A2(A[17]), .ZN(g[18]) );
  AND2_X1 U25 ( .A1(B[29]), .A2(A[29]), .ZN(g[30]) );
  AND2_X1 U26 ( .A1(B[28]), .A2(A[28]), .ZN(g[29]) );
  AND2_X1 U27 ( .A1(B[2]), .A2(A[2]), .ZN(g[3]) );
  AND2_X1 U28 ( .A1(B[3]), .A2(A[3]), .ZN(g[4]) );
  AND2_X1 U29 ( .A1(B[20]), .A2(A[20]), .ZN(g[21]) );
  AND2_X1 U30 ( .A1(B[21]), .A2(A[21]), .ZN(g[22]) );
  AND2_X1 U31 ( .A1(B[4]), .A2(A[4]), .ZN(g[5]) );
  AND2_X1 U32 ( .A1(B[5]), .A2(A[5]), .ZN(g[6]) );
  INV_X1 U33 ( .A(A[0]), .ZN(n3) );
  BUF_X1 U34 ( .A(\GG[1][5] ), .Z(n14) );
  AND2_X1 U35 ( .A1(B[15]), .A2(A[15]), .ZN(g[16]) );
  NAND2_X1 U37 ( .A1(n7), .A2(B[15]), .ZN(n8) );
  NAND2_X1 U60 ( .A1(n6), .A2(A[15]), .ZN(n9) );
  NAND2_X1 U64 ( .A1(n9), .A2(n8), .ZN(p[16]) );
  INV_X1 U67 ( .A(B[15]), .ZN(n6) );
  INV_X1 U68 ( .A(A[15]), .ZN(n7) );
  NAND2_X1 U69 ( .A1(B[11]), .A2(n11), .ZN(n12) );
  NAND2_X1 U70 ( .A1(n10), .A2(A[11]), .ZN(n13) );
  NAND2_X1 U71 ( .A1(n12), .A2(n13), .ZN(p[12]) );
  INV_X1 U72 ( .A(B[11]), .ZN(n10) );
  INV_X1 U73 ( .A(A[11]), .ZN(n11) );
  NAND2_X1 U74 ( .A1(n17), .A2(B[7]), .ZN(n18) );
  NAND2_X1 U75 ( .A1(n16), .A2(A[7]), .ZN(n19) );
  NAND2_X1 U76 ( .A1(n18), .A2(n19), .ZN(p[8]) );
  INV_X1 U77 ( .A(B[7]), .ZN(n16) );
  INV_X1 U78 ( .A(A[7]), .ZN(n17) );
  OAI21_X1 U79 ( .B1(n3), .B2(n4), .A(n5), .ZN(G_10) );
  INV_X1 U80 ( .A(B[0]), .ZN(n4) );
  OAI21_X1 U81 ( .B1(A[0]), .B2(B[0]), .A(C_in), .ZN(n5) );
  CLKBUF_X1 U82 ( .A(n24), .Z(C_o[1]) );
endmodule


module P4ADD_N32 ( A, B, C_in, S, C_o );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input C_in;
  output C_o;
  wire   n1;
  wire   [8:0] carry;

  CARRY_GENERATOR_N32 carry_gen ( .A(A), .B(B), .C_in(C_in), .C_o(carry) );
  SUM_GENERATOR_N32 sum_gen ( .A({A[31:4], n1, A[2:0]}), .B(B), .C_in(carry), 
        .O(S), .C_o(C_o) );
  BUF_X1 U1 ( .A(A[3]), .Z(n1) );
endmodule

