
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_register_file_reg_size64_file_size32_1 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_register_file_reg_size64_file_size32_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_register_file_reg_size64_file_size32_1.all;

entity register_file_reg_size64_file_size32_1 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_reg_size64_file_size32_1;

architecture SYN_BEHAVIORAL of register_file_reg_size64_file_size32_1 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal OUT1_63_port, OUT1_62_port, OUT1_61_port, OUT1_60_port, OUT1_59_port,
      OUT1_58_port, OUT1_57_port, OUT1_56_port, OUT1_55_port, OUT1_54_port, 
      OUT1_53_port, OUT1_52_port, OUT1_51_port, OUT1_50_port, OUT1_49_port, 
      OUT1_48_port, OUT1_47_port, OUT1_46_port, OUT1_45_port, OUT1_44_port, 
      OUT1_43_port, OUT1_42_port, OUT1_41_port, OUT1_40_port, OUT1_39_port, 
      OUT1_38_port, OUT1_37_port, OUT1_36_port, OUT1_35_port, OUT1_34_port, 
      OUT1_33_port, OUT1_32_port, OUT1_31_port, OUT1_30_port, OUT1_29_port, 
      OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, OUT1_24_port, 
      OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, OUT1_19_port, 
      OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, OUT1_14_port, 
      OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, OUT1_9_port, 
      OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, OUT1_4_port, 
      OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port, OUT2_63_port, 
      OUT2_62_port, OUT2_61_port, OUT2_60_port, OUT2_59_port, OUT2_58_port, 
      OUT2_57_port, OUT2_56_port, OUT2_55_port, OUT2_54_port, OUT2_53_port, 
      OUT2_52_port, OUT2_51_port, OUT2_50_port, OUT2_49_port, OUT2_48_port, 
      OUT2_47_port, OUT2_46_port, OUT2_45_port, OUT2_44_port, OUT2_43_port, 
      OUT2_42_port, OUT2_41_port, OUT2_40_port, OUT2_39_port, OUT2_38_port, 
      OUT2_37_port, OUT2_36_port, OUT2_35_port, OUT2_34_port, OUT2_33_port, 
      OUT2_32_port, OUT2_31_port, OUT2_30_port, OUT2_29_port, OUT2_28_port, 
      OUT2_27_port, OUT2_26_port, OUT2_25_port, OUT2_24_port, OUT2_23_port, 
      OUT2_22_port, OUT2_21_port, OUT2_20_port, OUT2_19_port, OUT2_18_port, 
      OUT2_17_port, OUT2_16_port, OUT2_15_port, OUT2_14_port, OUT2_13_port, 
      OUT2_12_port, OUT2_11_port, OUT2_10_port, OUT2_9_port, OUT2_8_port, 
      OUT2_7_port, OUT2_6_port, OUT2_5_port, OUT2_4_port, OUT2_3_port, 
      OUT2_2_port, OUT2_1_port, OUT2_0_port, n4093, n4094, n4095, n4096, n4097,
      n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, 
      n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, 
      n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, 
      n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, 
      n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, 
      n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4157, n4158, 
      n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, 
      n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, 
      n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, 
      n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, 
      n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, 
      n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, 
      n4219, n4220, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, 
      n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, 
      n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, 
      n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, 
      n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, 
      n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, 
      n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, 
      n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, 
      n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, 
      n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, 
      n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, 
      n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, 
      n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, 
      n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, 
      n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, 
      n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, 
      n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, 
      n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, 
      n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, 
      n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, 
      n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, 
      n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, 
      n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, 
      n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, 
      n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, 
      n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, 
      n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, 
      n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, 
      n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, 
      n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, 
      n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, 
      n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, 
      n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, 
      n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, 
      n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, 
      n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, 
      n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, 
      n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, 
      n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, 
      n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, 
      n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, 
      n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, 
      n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, 
      n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, 
      n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, 
      n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, 
      n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, 
      n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, 
      n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, 
      n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, 
      n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, 
      n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, 
      n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, 
      n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, 
      n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, 
      n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, 
      n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, 
      n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, 
      n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, 
      n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, 
      n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, 
      n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, 
      n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, 
      n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, 
      n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, 
      n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, 
      n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, 
      n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, 
      n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, 
      n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, 
      n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, 
      n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, 
      n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, 
      n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, 
      n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, 
      n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, 
      n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, 
      n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, 
      n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, 
      n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, 
      n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, 
      n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, 
      n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, 
      n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, 
      n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, 
      n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, 
      n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, 
      n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, 
      n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, 
      n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, 
      n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, 
      n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, 
      n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, 
      n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, 
      n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, 
      n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, 
      n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, 
      n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, 
      n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, 
      n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, 
      n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, 
      n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, 
      n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, 
      n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, 
      n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, 
      n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, 
      n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, 
      n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, 
      n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, 
      n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, 
      n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, 
      n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, 
      n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, 
      n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, 
      n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, 
      n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, 
      n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, 
      n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, 
      n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, 
      n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, 
      n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, 
      n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, 
      n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, 
      n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, 
      n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, 
      n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, 
      n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, 
      n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, 
      n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, 
      n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, 
      n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, 
      n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, 
      n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, 
      n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, 
      n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, 
      n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, 
      n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, 
      n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, 
      n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, 
      n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, 
      n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, 
      n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, 
      n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, 
      n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, 
      n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, 
      n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, 
      n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, 
      n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, 
      n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, 
      n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, 
      n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, 
      n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, 
      n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, 
      n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, 
      n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, 
      n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, 
      n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, 
      n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, 
      n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, 
      n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, 
      n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, 
      n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, 
      n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, 
      n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, 
      n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, 
      n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, 
      n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, 
      n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, 
      n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, 
      n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, 
      n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, 
      n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, 
      n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, 
      n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, 
      n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, 
      n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, 
      n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, 
      n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, 
      n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, 
      n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, 
      n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, 
      n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, 
      n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, 
      n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, 
      n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, 
      n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, 
      n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, 
      n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, 
      n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, 
      n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, 
      n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, 
      n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, 
      n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, 
      n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, 
      n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, 
      n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, 
      n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, 
      n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, 
      n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, 
      n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, 
      n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, 
      n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, 
      n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, 
      n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, 
      n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, 
      n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, 
      n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, 
      n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, 
      n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, 
      n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, 
      n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, 
      n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, 
      n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, 
      n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, 
      n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, 
      n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, 
      n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, 
      n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n8573, n8575, 
      n8576, n8577, n8579, n8580, n8581, n8583, n8584, n8585, n8587, n8588, 
      n8589, n8591, n8592, n8593, n8595, n8596, n8597, n8599, n8600, n8601, 
      n8603, n8604, n8605, n8607, n8608, n8609, n8611, n8612, n8613, n8615, 
      n8616, n8617, n8619, n8620, n8621, n8623, n8624, n8625, n8627, n8628, 
      n8629, n8631, n8632, n8633, n8635, n8636, n8637, n8639, n8640, n8641, 
      n8643, n8644, n8645, n8647, n8648, n8649, n8651, n8652, n8653, n8655, 
      n8656, n8657, n8659, n8660, n8661, n8663, n8664, n8665, n8667, n8668, 
      n8669, n8671, n8672, n8673, n8675, n8676, n8677, n8679, n8680, n8681, 
      n8683, n8684, n8685, n8687, n8688, n8689, n8691, n8692, n8693, n8695, 
      n8696, n8697, n8699, n8700, n8701, n8703, n8704, n8705, n8707, n8708, 
      n8709, n8711, n8712, n8713, n8715, n8716, n8717, n8719, n8720, n8721, 
      n8723, n8724, n8725, n8727, n8728, n8729, n8731, n8732, n8733, n8735, 
      n8736, n8737, n8739, n8740, n8741, n8743, n8744, n8745, n8747, n8748, 
      n8749, n8751, n8752, n8753, n8755, n8756, n8757, n8759, n8760, n8761, 
      n8763, n8764, n8765, n8767, n8768, n8769, n8771, n8772, n8773, n8775, 
      n8776, n8777, n8779, n8780, n8781, n8783, n8784, n8785, n8787, n8788, 
      n8789, n8791, n8792, n8793, n8795, n8796, n8797, n8799, n8800, n8801, 
      n8803, n8804, n8805, n8807, n8808, n8809, n8811, n8812, n8813, n8815, 
      n8816, n8817, n8819, n8820, n8821, n8823, n8824, n8825, n8827, n8828, 
      n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, 
      n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, 
      n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, 
      n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, 
      n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, 
      n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, 
      n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, 
      n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, 
      n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, 
      n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, 
      n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, 
      n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, 
      n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8959, 
      n8960, n8961, n8963, n8964, n8965, n8967, n8968, n8969, n8971, n8972, 
      n8973, n8975, n8976, n8977, n8979, n8980, n8981, n8983, n8984, n8985, 
      n8987, n8988, n8989, n8991, n8992, n8993, n8995, n8996, n8997, n8999, 
      n9000, n9001, n9003, n9004, n9005, n9007, n9008, n9009, n9011, n9012, 
      n9013, n9015, n9016, n9017, n9019, n9020, n9021, n9023, n9024, n9025, 
      n9027, n9028, n9029, n9031, n9032, n9033, n9035, n9036, n9037, n9039, 
      n9040, n9041, n9043, n9044, n9045, n9047, n9048, n9049, n9051, n9052, 
      n9053, n9055, n9056, n9057, n9059, n9060, n9061, n9063, n9064, n9065, 
      n9067, n9068, n9069, n9071, n9072, n9073, n9075, n9076, n9077, n9079, 
      n9080, n9081, n9083, n9084, n9085, n9087, n9088, n9089, n9091, n9092, 
      n9093, n9095, n9096, n9097, n9099, n9100, n9101, n9103, n9104, n9105, 
      n9107, n9108, n9109, n9111, n9112, n9113, n9115, n9116, n9117, n9119, 
      n9120, n9121, n9123, n9124, n9125, n9127, n9128, n9129, n9131, n9132, 
      n9133, n9135, n9136, n9137, n9139, n9140, n9141, n9143, n9144, n9145, 
      n9147, n9148, n9149, n9151, n9152, n9153, n9155, n9156, n9157, n9159, 
      n9160, n9161, n9163, n9164, n9165, n9167, n9168, n9169, n9171, n9172, 
      n9173, n9175, n9176, n9177, n9179, n9180, n9181, n9183, n9184, n9185, 
      n9187, n9188, n9189, n9191, n9192, n9193, n9195, n9196, n9197, n9199, 
      n9200, n9201, n9203, n9204, n9205, n9207, n9208, n9209, n9211, n9212, 
      n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947, 
      n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955, n13956, 
      n13957, n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965, 
      n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973, n13974, 
      n13975, n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983, 
      n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992, 
      n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000, n14001, 
      n14002, n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010, 
      n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019, 
      n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027, n14028, 
      n14029, n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037, 
      n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045, n14046, 
      n14047, n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055, 
      n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064, 
      n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072, n14073, 
      n14074, n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082, 
      n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091, 
      n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099, n14100, 
      n14101, n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109, 
      n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117, n14118, 
      n14119, n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127, 
      n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136, 
      n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144, n14145, 
      n14146, n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154, 
      n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163, 
      n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171, n14172, 
      n14173, n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181, 
      n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189, n14190, 
      n14191, n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199, 
      n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208, 
      n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216, n14217, 
      n14218, n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226, 
      n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235, 
      n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243, n14244, 
      n14245, n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253, 
      n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261, n14262, 
      n14263, n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271, 
      n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280, 
      n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288, n14289, 
      n14290, n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298, 
      n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307, 
      n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315, n14316, 
      n14317, n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325, 
      n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333, n14334, 
      n14335, n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343, 
      n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352, 
      n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360, n14361, 
      n14362, n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370, 
      n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379, 
      n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387, n14388, 
      n14389, n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397, 
      n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405, n14406, 
      n14407, n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415, 
      n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424, 
      n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432, n14433, 
      n14434, n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442, 
      n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451, 
      n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459, n14460, 
      n14461, n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469, 
      n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477, n14478, 
      n14479, n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487, 
      n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496, 
      n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504, n14505, 
      n14506, n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514, 
      n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523, 
      n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531, n14532, 
      n14533, n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541, 
      n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549, n14550, 
      n14551, n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559, 
      n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568, 
      n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576, n14577, 
      n14578, n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586, 
      n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595, 
      n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603, n14604, 
      n14605, n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613, 
      n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621, n14622, 
      n14623, n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631, 
      n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640, 
      n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648, n14649, 
      n14650, n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658, 
      n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667, 
      n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675, n14676, 
      n14677, n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685, 
      n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693, n14694, 
      n14695, n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703, 
      n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712, 
      n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720, n14721, 
      n14722, n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730, 
      n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739, 
      n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747, n14748, 
      n14749, n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757, 
      n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765, n14766, 
      n14767, n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775, 
      n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784, 
      n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792, n14793, 
      n14794, n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802, 
      n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811, 
      n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819, n14820, 
      n14821, n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829, 
      n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837, n14838, 
      n14839, n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847, 
      n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856, 
      n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864, n14865, 
      n14866, n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874, 
      n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883, 
      n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891, n14892, 
      n14893, n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901, 
      n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909, n14910, 
      n14911, n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919, 
      n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928, 
      n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936, n14937, 
      n14938, n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946, 
      n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955, 
      n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963, n14964, 
      n14965, n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973, 
      n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981, n14982, 
      n14983, n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991, 
      n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000, 
      n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008, n15009, 
      n15010, n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018, 
      n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027, 
      n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035, n15036, 
      n15037, n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045, 
      n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053, n15054, 
      n15055, n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063, 
      n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072, 
      n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080, n15081, 
      n15082, n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090, 
      n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099, 
      n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107, n15108, 
      n15109, n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117, 
      n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125, n15126, 
      n15127, n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135, 
      n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144, 
      n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152, n15153, 
      n15154, n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162, 
      n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171, 
      n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179, n15180, 
      n15181, n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189, 
      n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197, n15198, 
      n15199, n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207, 
      n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216, 
      n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224, n15225, 
      n15226, n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234, 
      n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243, 
      n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251, n15252, 
      n15253, n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261, 
      n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269, n15270, 
      n15271, n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279, 
      n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288, 
      n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296, n15297, 
      n15298, n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306, 
      n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315, 
      n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323, n15324, 
      n15325, n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333, 
      n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341, n15342, 
      n15343, n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351, 
      n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360, 
      n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368, n15369, 
      n15370, n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378, 
      n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387, 
      n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395, n15396, 
      n15397, n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405, 
      n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413, n15414, 
      n15415, n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423, 
      n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432, 
      n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440, n15441, 
      n15442, n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450, 
      n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459, 
      n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467, n15468, 
      n15469, n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477, 
      n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485, n15486, 
      n15487, n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495, 
      n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504, 
      n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512, n15513, 
      n15514, n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522, 
      n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531, 
      n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539, n15540, 
      n15541, n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549, 
      n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557, n15558, 
      n15559, n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567, 
      n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576, 
      n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584, n15585, 
      n15586, n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594, 
      n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603, 
      n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611, n15612, 
      n15613, n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621, 
      n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629, n15630, 
      n15631, n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639, 
      n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648, 
      n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656, n15657, 
      n15658, n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666, 
      n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675, 
      n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683, n15684, 
      n15685, n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693, 
      n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701, n15702, 
      n15703, n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711, 
      n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720, 
      n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728, n15729, 
      n15730, n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738, 
      n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747, 
      n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755, n15756, 
      n15757, n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765, 
      n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773, n15774, 
      n15775, n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783, 
      n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792, 
      n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800, n15801, 
      n15802, n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810, 
      n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819, 
      n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827, n15828, 
      n15829, n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837, 
      n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845, n15846, 
      n15847, n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855, 
      n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864, 
      n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872, n15873, 
      n15874, n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882, 
      n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891, 
      n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899, n15900, 
      n15901, n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909, 
      n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917, n15918, 
      n15919, n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927, 
      n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936, 
      n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944, n15945, 
      n15946, n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954, 
      n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963, 
      n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971, n15972, 
      n15973, n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981, 
      n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989, n15990, 
      n15991, n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999, 
      n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008, 
      n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016, n16017, 
      n16018, n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026, 
      n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035, 
      n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043, n16044, 
      n16045, n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053, 
      n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061, n16062, 
      n16063, n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071, 
      n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080, 
      n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088, n16089, 
      n16090, n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098, 
      n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107, 
      n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115, n16116, 
      n16117, n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125, 
      n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133, n16134, 
      n16135, n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143, 
      n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152, 
      n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160, n16161, 
      n16162, n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170, 
      n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179, 
      n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187, n16188, 
      n16189, n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197, 
      n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205, n16206, 
      n16207, n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215, 
      n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224, 
      n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232, n16233, 
      n16234, n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242, 
      n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251, 
      n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259, n16260, 
      n16261, n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269, 
      n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277, n16278, 
      n16279, n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287, 
      n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296, 
      n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304, n16305, 
      n16306, n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314, 
      n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323, 
      n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331, n16332, 
      n16333, n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341, 
      n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349, n16350, 
      n16351, n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359, 
      n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368, 
      n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376, n16377, 
      n16378, n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386, 
      n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395, 
      n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403, n16404, 
      n16405, n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413, 
      n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421, n16422, 
      n16423, n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431, 
      n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440, 
      n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448, n16449, 
      n16450, n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458, 
      n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467, 
      n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475, n16476, 
      n16477, n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485, 
      n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493, n16494, 
      n16495, n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503, 
      n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512, 
      n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520, n16521, 
      n16522, n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530, 
      n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539, 
      n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547, n16548, 
      n16549, n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557, 
      n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565, n16566, 
      n16567, n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575, 
      n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584, 
      n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592, n16593, 
      n16594, n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602, 
      n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611, 
      n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619, n16620, 
      n16621, n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629, 
      n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637, n16638, 
      n16639, n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647, 
      n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656, 
      n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664, n16665, 
      n16666, n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674, 
      n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683, 
      n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691, n16692, 
      n16693, n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701, 
      n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709, n16710, 
      n16711, n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719, 
      n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728, 
      n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736, n16737, 
      n16738, n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746, 
      n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755, 
      n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763, n16764, 
      n16765, n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773, 
      n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781, n16782, 
      n16783, n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791, 
      n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800, 
      n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808, n16809, 
      n16810, n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818, 
      n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827, 
      n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835, n16836, 
      n16837, n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845, 
      n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853, n16854, 
      n16855, n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863, 
      n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872, 
      n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880, n16881, 
      n16882, n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890, 
      n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899, 
      n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907, n16908, 
      n16909, n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917, 
      n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925, n16926, 
      n16927, n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935, 
      n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944, 
      n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952, n16953, 
      n16954, n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962, 
      n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971, 
      n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979, n16980, 
      n16981, n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989, 
      n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997, n16998, 
      n16999, n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007, 
      n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016, 
      n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024, n17025, 
      n17026, n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034, 
      n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043, 
      n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051, n17052, 
      n17053, n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061, 
      n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069, n17070, 
      n17071, n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079, 
      n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088, 
      n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096, n17097, 
      n17098, n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106, 
      n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115, 
      n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123, n17124, 
      n17125, n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133, 
      n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141, n17142, 
      n17143, n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151, 
      n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160, 
      n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168, n17169, 
      n17170, n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178, 
      n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187, 
      n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195, n17196, 
      n17197, n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205, 
      n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213, n17214, 
      n17215, n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223, 
      n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232, 
      n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240, n17241, 
      n17242, n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250, 
      n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259, 
      n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267, n17268, 
      n17269, n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277, 
      n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285, n17286, 
      n17287, n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295, 
      n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304, 
      n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312, n17313, 
      n17314, n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322, 
      n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331, 
      n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339, n17340, 
      n17341, n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349, 
      n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357, n17358, 
      n17359, n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367, 
      n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376, 
      n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384, n17385, 
      n17386, n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394, 
      n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403, 
      n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411, n17412, 
      n17413, n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421, 
      n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429, n17430, 
      n17431, n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439, 
      n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448, 
      n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456, n17457, 
      n17458, n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466, 
      n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475, 
      n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483, n17484, 
      n17485, n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493, 
      n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501, n17502, 
      n17503, n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511, 
      n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520, 
      n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528, n17529, 
      n17530, n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538, 
      n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547, 
      n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555, n17556, 
      n17557, n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565, 
      n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573, n17574, 
      n17575, n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583, 
      n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592, 
      n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600, n17601, 
      n17602, n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610, 
      n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619, 
      n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627, n17628, 
      n17629, n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637, 
      n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645, n17646, 
      n17647, n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655, 
      n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664, 
      n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672, n17673, 
      n17674, n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682, 
      n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691, 
      n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699, n17700, 
      n17701, n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709, 
      n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717, n17718, 
      n17719, n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727, 
      n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736, 
      n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744, n17745, 
      n17746, n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754, 
      n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763, 
      n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771, n17772, 
      n17773, n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781, 
      n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789, n17790, 
      n17791, n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799, 
      n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808, 
      n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816, n17817, 
      n17818, n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826, 
      n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835, 
      n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843, n17844, 
      n17845, n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853, 
      n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861, n17862, 
      n17863, n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871, 
      n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880, 
      n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888, n17889, 
      n17890, n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898, 
      n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907, 
      n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915, n17916, 
      n17917, n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925, 
      n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933, n17934, 
      n17935, n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943, 
      n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952, 
      n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960, n17961, 
      n17962, n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970, 
      n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979, 
      n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987, n17988, 
      n17989, n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997, 
      n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005, n18006, 
      n18007, n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015, 
      n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024, 
      n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032, n18033, 
      n18034, n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042, 
      n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051, 
      n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059, n18060, 
      n18061, n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069, 
      n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077, n18078, 
      n18079, n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087, 
      n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096, 
      n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104, n18105, 
      n18106, n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114, 
      n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123, 
      n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131, n18132, 
      n18133, n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141, 
      n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149, n18150, 
      n18151, n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159, 
      n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168, 
      n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176, n18177, 
      n18178, n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186, 
      n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195, 
      n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203, n18204, 
      n18205, n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213, 
      n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221, n18222, 
      n18223, n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231, 
      n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240, 
      n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248, n18249, 
      n18250, n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258, 
      n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267, 
      n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275, n18276, 
      n18277, n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285, 
      n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293, n18294, 
      n18295, n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303, 
      n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312, 
      n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320, n18321, 
      n18322, n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330, 
      n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339, 
      n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347, n18348, 
      n18349, n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357, 
      n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365, n18366, 
      n18367, n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375, 
      n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384, 
      n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392, n18393, 
      n18394, n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402, 
      n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411, 
      n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419, n18420, 
      n18421, n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429, 
      n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437, n18438, 
      n18439, n18440, n18441, n18442, n18443, n18444, n18445, n18446, n18447, 
      n18448, n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456, 
      n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464, n18465, 
      n18466, n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474, 
      n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483, 
      n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491, n18492, 
      n18493, n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501, 
      n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509, n18510, 
      n18511, n18512, n18513, n18514, n18515, n18516, n18517, n18518, n18519, 
      n18520, n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528, 
      n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536, n18537, 
      n18538, n18539, n18540, n18541, n18544, n18545, n18548, n18549, n18550, 
      n18551, n18554, n18555, n18559, n18561, n18564, n18565, n18568, n18569, 
      n18570, n18571, n18574, n18575, n18579, n18581, n18584, n18585, n18588, 
      n18589, n18590, n18591, n18594, n18595, n18599, n18601, n18604, n18605, 
      n18608, n18609, n18610, n18611, n18614, n18615, n18619, n18621, n18624, 
      n18625, n18628, n18629, n18630, n18631, n18634, n18635, n18639, n18641, 
      n18644, n18645, n18648, n18649, n18650, n18651, n18654, n18655, n18659, 
      n18661, n18664, n18665, n18668, n18669, n18670, n18671, n18674, n18675, 
      n18679, n18681, n18684, n18685, n18688, n18689, n18690, n18691, n18694, 
      n18695, n18699, n18701, n18704, n18705, n18708, n18709, n18710, n18711, 
      n18714, n18715, n18719, n18721, n18724, n18725, n18728, n18729, n18730, 
      n18731, n18734, n18735, n18739, n18741, n18744, n18745, n18748, n18749, 
      n18750, n18751, n18754, n18755, n18759, n18761, n18764, n18765, n18768, 
      n18769, n18770, n18771, n18774, n18775, n18779, n18781, n18784, n18785, 
      n18788, n18789, n18790, n18791, n18794, n18795, n18799, n18801, n18804, 
      n18805, n18808, n18809, n18810, n18811, n18814, n18815, n18819, n18821, 
      n18824, n18825, n18828, n18829, n18830, n18831, n18834, n18835, n18839, 
      n18841, n18844, n18845, n18848, n18849, n18850, n18851, n18854, n18855, 
      n18859, n18861, n18864, n18865, n18868, n18869, n18870, n18871, n18874, 
      n18875, n18879, n18881, n18884, n18885, n18888, n18889, n18890, n18891, 
      n18894, n18895, n18899, n18901, n18904, n18905, n18908, n18909, n18910, 
      n18911, n18914, n18915, n18919, n18921, n18924, n18925, n18928, n18929, 
      n18930, n18931, n18934, n18935, n18939, n18941, n18944, n18945, n18948, 
      n18949, n18950, n18951, n18954, n18955, n18959, n18961, n18964, n18965, 
      n18968, n18969, n18970, n18971, n18974, n18975, n18979, n18981, n18984, 
      n18985, n18988, n18989, n18990, n18991, n18994, n18995, n18999, n19001, 
      n19004, n19005, n19008, n19009, n19010, n19011, n19014, n19015, n19019, 
      n19021, n19024, n19025, n19028, n19029, n19030, n19031, n19034, n19035, 
      n19039, n19041, n19044, n19045, n19048, n19049, n19050, n19051, n19054, 
      n19055, n19059, n19061, n19064, n19065, n19068, n19069, n19070, n19071, 
      n19074, n19075, n19079, n19081, n19084, n19085, n19088, n19089, n19090, 
      n19091, n19094, n19095, n19099, n19101, n19104, n19105, n19108, n19109, 
      n19110, n19111, n19114, n19115, n19119, n19121, n19124, n19125, n19128, 
      n19129, n19130, n19131, n19134, n19135, n19139, n19141, n19144, n19145, 
      n19148, n19149, n19150, n19151, n19154, n19155, n19159, n19161, n19164, 
      n19165, n19168, n19169, n19170, n19171, n19174, n19175, n19179, n19181, 
      n19184, n19185, n19188, n19189, n19190, n19191, n19194, n19195, n19199, 
      n19201, n19204, n19205, n19208, n19209, n19210, n19211, n19214, n19215, 
      n19219, n19221, n19224, n19225, n19228, n19229, n19230, n19231, n19234, 
      n19235, n19239, n19241, n19244, n19245, n19248, n19249, n19250, n19251, 
      n19254, n19255, n19259, n19261, n19264, n19265, n19268, n19269, n19270, 
      n19271, n19274, n19275, n19279, n19281, n19284, n19285, n19288, n19289, 
      n19290, n19291, n19294, n19295, n19299, n19301, n19304, n19305, n19308, 
      n19309, n19310, n19311, n19314, n19315, n19319, n19321, n19324, n19325, 
      n19328, n19329, n19330, n19331, n19334, n19335, n19339, n19341, n19344, 
      n19345, n19348, n19349, n19350, n19351, n19354, n19355, n19359, n19361, 
      n19364, n19365, n19368, n19369, n19370, n19371, n19374, n19375, n19379, 
      n19381, n19384, n19385, n19388, n19389, n19390, n19391, n19394, n19395, 
      n19399, n19401, n19404, n19405, n19408, n19409, n19410, n19411, n19414, 
      n19415, n19419, n19421, n19424, n19425, n19428, n19429, n19430, n19431, 
      n19434, n19435, n19439, n19441, n19444, n19445, n19448, n19449, n19450, 
      n19451, n19454, n19455, n19459, n19461, n19464, n19465, n19468, n19469, 
      n19470, n19471, n19474, n19475, n19479, n19481, n19484, n19485, n19488, 
      n19489, n19490, n19491, n19494, n19495, n19499, n19501, n19504, n19505, 
      n19508, n19509, n19510, n19511, n19514, n19515, n19519, n19521, n19524, 
      n19525, n19528, n19529, n19530, n19531, n19534, n19535, n19539, n19541, 
      n19544, n19545, n19548, n19549, n19550, n19551, n19554, n19555, n19559, 
      n19561, n19564, n19565, n19568, n19569, n19570, n19571, n19574, n19575, 
      n19579, n19581, n19584, n19585, n19588, n19589, n19590, n19591, n19594, 
      n19595, n19599, n19601, n19604, n19605, n19608, n19609, n19610, n19611, 
      n19614, n19615, n19619, n19621, n19624, n19625, n19628, n19629, n19630, 
      n19631, n19634, n19635, n19639, n19641, n19644, n19645, n19648, n19649, 
      n19650, n19651, n19654, n19655, n19659, n19661, n19664, n19665, n19668, 
      n19669, n19670, n19671, n19674, n19675, n19679, n19681, n19684, n19685, 
      n19688, n19689, n19690, n19691, n19694, n19695, n19699, n19701, n19704, 
      n19705, n19708, n19709, n19710, n19711, n19714, n19715, n19719, n19721, 
      n19724, n19725, n19728, n19729, n19730, n19731, n19734, n19735, n19739, 
      n19741, n19744, n19745, n19748, n19749, n19750, n19751, n19754, n19755, 
      n19759, n19761, n19764, n19765, n19768, n19769, n19770, n19771, n19774, 
      n19775, n19779, n19781, n19784, n19785, n19788, n19789, n19790, n19791, 
      n19794, n19795, n19799, n19801, n19804, n19805, n19808, n19809, n19810, 
      n19811, n19814, n19815, n19819, n19821, n19822, n19823, n19824, n19825, 
      n19826, n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834, 
      n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843, 
      n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851, n19852, 
      n19853, n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861, 
      n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869, n19870, 
      n19871, n19872, n19873, n19874, n19875, n19876, n19877, n19878, n19879, 
      n19880, n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888, 
      n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896, n19897, 
      n19898, n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906, 
      n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915, 
      n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923, n19924, 
      n19925, n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933, 
      n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941, n19942, 
      n19943, n19944, n19945, n19946, n19947, n19948, n19949, n19950, n19951, 
      n19952, n19953, n19954, n19955, n19956, n19957, n19958, n19959, n19960, 
      n19961, n19962, n19963, n19964, n19965, n19966, n19967, n19968, n19969, 
      n19970, n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978, 
      n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987, 
      n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995, n19996, 
      n19997, n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005, 
      n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013, n20014, 
      n20015, n20016, n20017, n20018, n20019, n20020, n20021, n20022, n20023, 
      n20024, n20025, n20026, n20027, n20028, n20029, n20030, n20031, n20032, 
      n20033, n20034, n20035, n20036, n20037, n20038, n20039, n20040, n20041, 
      n20042, n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050, 
      n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059, 
      n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067, n20068, 
      n20069, n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077, 
      n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085, n20086, 
      n20087, n20088, n20089, n20090, n20091, n20092, n20093, n20094, n20095, 
      n20096, n20097, n20098, n20099, n20100, n20101, n20102, n20103, n20104, 
      n20105, n20106, n20107, n20108, n20109, n20110, n20111, n20112, n20113, 
      n20114, n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122, 
      n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131, 
      n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139, n20140, 
      n20141, n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149, 
      n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157, n20158, 
      n20159, n20160, n20161, n20162, n20163, n20164, n20165, n20166, n20167, 
      n20168, n20169, n20170, n20171, n20172, n20173, n20174, n20175, n20176, 
      n20177, n20178, n20179, n20180, n20181, n20182, n20183, n20184, n20185, 
      n20186, n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194, 
      n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203, 
      n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211, n20212, 
      n20213, n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221, 
      n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229, n20230, 
      n20231, n20232, n20233, n20234, n20235, n20236, n20237, n20238, n20239, 
      n20240, n20241, n20242, n20243, n20244, n20245, n20246, n20247, n20248, 
      n20249, n20250, n20251, n20252, n20253, n20254, n20255, n20256, n20257, 
      n20258, n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266, 
      n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275, 
      n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283, n20284, 
      n20285, n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293, 
      n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301, n20302, 
      n20303, n20304, n20305, n20306, n20307, n20308, n20309, n20310, n20311, 
      n20312, n20313, n20314, n20315, n20316, n20317, n20318, n20319, n20320, 
      n20321, n20322, n20323, n20324, n20325, n20326, n20327, n20328, n20329, 
      n20330, n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338, 
      n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347, 
      n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355, n20356, 
      n20357, n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365, 
      n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373, n20374, 
      n20375, n20376, n20377, n20378, n20379, n20380, n20381, n20382, n20383, 
      n20384, n20385, n20386, n20387, n20388, n20389, n20390, n20391, n20392, 
      n20393, n20394, n20395, n20396, n20397, n20398, n20399, n20400, n20401, 
      n20402, n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410, 
      n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419, 
      n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427, n20428, 
      n20429, n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437, 
      n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445, n20446, 
      n20447, n20448, n20449, n20450, n20451, n20452, n20453, n20454, n20455, 
      n20456, n20457, n20458, n20459, n20460, n20461, n20462, n20463, n20464, 
      n20465, n20466, n20467, n20468, n20469, n20470, n20471, n20472, n20473, 
      n20474, n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482, 
      n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491, 
      n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499, n20500, 
      n20501, n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509, 
      n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517, n20518, 
      n20519, n20520, n20521, n20522, n20523, n20524, n20525, n20526, n20527, 
      n20528, n20529, n20530, n20531, n20532, n20533, n20534, n20535, n20536, 
      n20537, n20538, n20539, n20540, n20541, n20542, n20543, n20544, n20545, 
      n20546, n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554, 
      n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563, 
      n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571, n20572, 
      n20573, n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581, 
      n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589, n20590, 
      n20591, n20592, n20593, n20594, n20595, n20596, n20597, n20598, n20599, 
      n20600, n20601, n20602, n20603, n20604, n20605, n20606, n20607, n20608, 
      n20609, n20610, n20611, n20612, n20613, n20614, n20615, n20616, n20617, 
      n20618, n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626, 
      n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635, 
      n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643, n20644, 
      n20645, n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653, 
      n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661, n20662, 
      n20663, n20664, n20665, n20666, n20667, n20668, n20669, n20670, n20671, 
      n20672, n20673, n20674, n20675, n20676, n20677, n20678, n20679, n20680, 
      n20681, n20682, n20683, n20684, n20685, n20686, n20687, n20688, n20689, 
      n20690, n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698, 
      n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707, 
      n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715, n20716, 
      n20717, n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725, 
      n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733, n20734, 
      n20735, n20736, n20737, n20738, n20739, n20740, n20741, n20742, n20743, 
      n20744, n20745, n20746, n20747, n20748, n20749, n20750, n20751, n20752, 
      n20753, n20754, n20755, n20756, n20757, n20758, n20759, n20760, n20761, 
      n20762, n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770, 
      n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779, 
      n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787, n20788, 
      n20789, n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797, 
      n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805, n20806, 
      n20807, n20808, n20809, n20810, n20811, n20812, n20813, n20814, n20815, 
      n20816, n20817, n20818, n20819, n20820, n20821, n20822, n20823, n20824, 
      n20825, n20826, n20827, n20828, n20829, n20830, n20831, n20832, n20833, 
      n20834, n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842, 
      n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851, 
      n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859, n20860, 
      n20861, n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869, 
      n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877, n20878, 
      n20879, n20880, n20881, n20882, n20883, n20884, n20885, n20886, n20887, 
      n20888, n20889, n20890, n20891, n20892, n20893, n20894, n20895, n20896, 
      n20897, n20898, n20899, n20900, n20901, n20902, n20903, n20904, n20905, 
      n20906, n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914, 
      n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923, 
      n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931, n20932, 
      n20933, n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941, 
      n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949, n20950, 
      n20951, n20952, n20953, n20954, n20955, n20956, n20957, n20958, n20959, 
      n20960, n20961, n20962, n20963, n20964, n20965, n20966, n20967, n20968, 
      n20969, n20970, n20971, n20972, n20973, n20974, n20975, n20976, n20977, 
      n20978, n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986, 
      n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995, 
      n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003, n21004, 
      n21005, n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013, 
      n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021, n21022, 
      n21023, n21024, n21025, n21026, n21027, n21028, n21029, n21030, n21031, 
      n21032, n21033, n21034, n21035, n21036, n21037, n21038, n21039, n21040, 
      n21041, n21042, n21043, n21044, n21045, n21046, n21047, n21048, n21049, 
      n21050, n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058, 
      n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067, 
      n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075, n21076, 
      n21077, n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085, 
      n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093, n21094, 
      n21095, n21096, n21097, n21098, n21099, n21100, n21101, n21102, n21103, 
      n21104, n21105, n21106, n21107, n21108, n21109, n21110, n21111, n21112, 
      n21113, n21114, n21115, n21116, n21117, n21118, n21119, n21120, n21121, 
      n21122, n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130, 
      n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139, 
      n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147, n21148, 
      n21149, n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157, 
      n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165, n21166, 
      n21167, n21168, n21169, n21170, n21171, n21172, n21173, n21174, n21175, 
      n21176, n21177, n21178, n21179, n21180, n21181, n21182, n21183, n21184, 
      n21185, n21186, n21187, n21188, n21189, n21190, n21191, n21192, n21193, 
      n21194, n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202, 
      n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211, 
      n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219, n21220, 
      n21221, n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229, 
      n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237, n21238, 
      n21239, n21240, n21241, n21242, n21243, n21244, n21245, n21246, n21247, 
      n21248, n21249, n21250, n21251, n21252, n21253, n21254, n21255, n21256, 
      n21257, n21258, n21259, n21260, n21261, n21262, n21263, n21264, n21265, 
      n21266, n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274, 
      n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283, 
      n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291, n21292, 
      n21293, n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301, 
      n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309, n21310, 
      n21311, n21312, n21313, n21314, n21315, n21316, n21317, n21318, n21319, 
      n21320, n21321, n21322, n21323, n21324, n21325, n21326, n21327, n21328, 
      n21329, n21330, n21331, n21332, n21333, n21334, n21335, n21336, n21337, 
      n21338, n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346, 
      n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355, 
      n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363, n21364, 
      n21365, n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373, 
      n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381, n21382, 
      n21383, n21384, n21385, n21386, n21387, n21388, n21389, n21390, n21391, 
      n21392, n21393, n21394, n21395, n21396, n21397, n21398, n21399, n21400, 
      n21401, n21402, n21403, n21404, n21405, n21406, n21407, n21408, n21409, 
      n21410, n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418, 
      n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427, 
      n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435, n21436, 
      n21437, n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445, 
      n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453, n21454, 
      n21455, n21456, n21457, n21458, n21459, n21460, n21461, n21462, n21463, 
      n21464, n21465, n21466, n21467, n21468, n21469, n21470, n21471, n21472, 
      n21473, n21474, n21475, n21476, n21477, n21478, n21479, n21480, n21481, 
      n21482, n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490, 
      n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499, 
      n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507, n21508, 
      n21509, n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517, 
      n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525, n21526, 
      n21527, n21528, n21529, n21530, n21531, n21532, n21533, n21534, n21535, 
      n21536, n21537, n21538, n21539, n21540, n21541, n21542, n21543, n21544, 
      n21545, n21546, n21547, n21548, n21549, n21550, n21551, n21552, n21553, 
      n21554, n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562, 
      n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571, 
      n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579, n21580, 
      n21581, n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589, 
      n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597, n21598, 
      n21599, n21600, n21601, n21602, n21603, n21604, n21605, n21606, n21607, 
      n21608, n21609, n21610, n21611, n21612, n21613, n21614, n21615, n21616, 
      n21617, n21618, n21619, n21620, n21621, n21622, n21623, n21624, n21625, 
      n21626, n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634, 
      n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643, 
      n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651, n21652, 
      n21653, n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661, 
      n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669, n21670, 
      n21671, n21672, n21673, n21674, n21675, n21676, n21677, n21678, n21679, 
      n21680, n21681, n21682, n21683, n21684, n21685, n21686, n21687, n21688, 
      n21689, n21690, n21691, n21692, n21693, n21694, n21695, n21696, n21697, 
      n21698, n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706, 
      n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715, 
      n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723, n21724, 
      n21725, n21726, n21727, n21728, n21729, n21730 : std_logic;

begin
   OUT1 <= ( OUT1_63_port, OUT1_62_port, OUT1_61_port, OUT1_60_port, 
      OUT1_59_port, OUT1_58_port, OUT1_57_port, OUT1_56_port, OUT1_55_port, 
      OUT1_54_port, OUT1_53_port, OUT1_52_port, OUT1_51_port, OUT1_50_port, 
      OUT1_49_port, OUT1_48_port, OUT1_47_port, OUT1_46_port, OUT1_45_port, 
      OUT1_44_port, OUT1_43_port, OUT1_42_port, OUT1_41_port, OUT1_40_port, 
      OUT1_39_port, OUT1_38_port, OUT1_37_port, OUT1_36_port, OUT1_35_port, 
      OUT1_34_port, OUT1_33_port, OUT1_32_port, OUT1_31_port, OUT1_30_port, 
      OUT1_29_port, OUT1_28_port, OUT1_27_port, OUT1_26_port, OUT1_25_port, 
      OUT1_24_port, OUT1_23_port, OUT1_22_port, OUT1_21_port, OUT1_20_port, 
      OUT1_19_port, OUT1_18_port, OUT1_17_port, OUT1_16_port, OUT1_15_port, 
      OUT1_14_port, OUT1_13_port, OUT1_12_port, OUT1_11_port, OUT1_10_port, 
      OUT1_9_port, OUT1_8_port, OUT1_7_port, OUT1_6_port, OUT1_5_port, 
      OUT1_4_port, OUT1_3_port, OUT1_2_port, OUT1_1_port, OUT1_0_port );
   OUT2 <= ( OUT2_63_port, OUT2_62_port, OUT2_61_port, OUT2_60_port, 
      OUT2_59_port, OUT2_58_port, OUT2_57_port, OUT2_56_port, OUT2_55_port, 
      OUT2_54_port, OUT2_53_port, OUT2_52_port, OUT2_51_port, OUT2_50_port, 
      OUT2_49_port, OUT2_48_port, OUT2_47_port, OUT2_46_port, OUT2_45_port, 
      OUT2_44_port, OUT2_43_port, OUT2_42_port, OUT2_41_port, OUT2_40_port, 
      OUT2_39_port, OUT2_38_port, OUT2_37_port, OUT2_36_port, OUT2_35_port, 
      OUT2_34_port, OUT2_33_port, OUT2_32_port, OUT2_31_port, OUT2_30_port, 
      OUT2_29_port, OUT2_28_port, OUT2_27_port, OUT2_26_port, OUT2_25_port, 
      OUT2_24_port, OUT2_23_port, OUT2_22_port, OUT2_21_port, OUT2_20_port, 
      OUT2_19_port, OUT2_18_port, OUT2_17_port, OUT2_16_port, OUT2_15_port, 
      OUT2_14_port, OUT2_13_port, OUT2_12_port, OUT2_11_port, OUT2_10_port, 
      OUT2_9_port, OUT2_8_port, OUT2_7_port, OUT2_6_port, OUT2_5_port, 
      OUT2_4_port, OUT2_3_port, OUT2_2_port, OUT2_1_port, OUT2_0_port );
   
   OUT1_reg_63_inst : DFF_X1 port map( D => n5435, CK => CLK, Q => OUT1_63_port
                           , QN => n4220);
   OUT1_reg_62_inst : DFF_X1 port map( D => n5433, CK => CLK, Q => OUT1_62_port
                           , QN => n4219);
   OUT1_reg_61_inst : DFF_X1 port map( D => n5431, CK => CLK, Q => OUT1_61_port
                           , QN => n4218);
   OUT1_reg_60_inst : DFF_X1 port map( D => n5429, CK => CLK, Q => OUT1_60_port
                           , QN => n4217);
   OUT1_reg_59_inst : DFF_X1 port map( D => n5427, CK => CLK, Q => OUT1_59_port
                           , QN => n4216);
   OUT1_reg_58_inst : DFF_X1 port map( D => n5425, CK => CLK, Q => OUT1_58_port
                           , QN => n4215);
   OUT1_reg_57_inst : DFF_X1 port map( D => n5423, CK => CLK, Q => OUT1_57_port
                           , QN => n4214);
   OUT1_reg_56_inst : DFF_X1 port map( D => n5421, CK => CLK, Q => OUT1_56_port
                           , QN => n4213);
   OUT1_reg_55_inst : DFF_X1 port map( D => n5419, CK => CLK, Q => OUT1_55_port
                           , QN => n4212);
   OUT1_reg_54_inst : DFF_X1 port map( D => n5417, CK => CLK, Q => OUT1_54_port
                           , QN => n4211);
   OUT1_reg_53_inst : DFF_X1 port map( D => n5415, CK => CLK, Q => OUT1_53_port
                           , QN => n4210);
   OUT1_reg_52_inst : DFF_X1 port map( D => n5413, CK => CLK, Q => OUT1_52_port
                           , QN => n4209);
   OUT1_reg_51_inst : DFF_X1 port map( D => n5411, CK => CLK, Q => OUT1_51_port
                           , QN => n4208);
   OUT1_reg_50_inst : DFF_X1 port map( D => n5409, CK => CLK, Q => OUT1_50_port
                           , QN => n4207);
   OUT1_reg_49_inst : DFF_X1 port map( D => n5407, CK => CLK, Q => OUT1_49_port
                           , QN => n4206);
   OUT1_reg_48_inst : DFF_X1 port map( D => n5405, CK => CLK, Q => OUT1_48_port
                           , QN => n4205);
   OUT1_reg_47_inst : DFF_X1 port map( D => n5403, CK => CLK, Q => OUT1_47_port
                           , QN => n4204);
   OUT1_reg_46_inst : DFF_X1 port map( D => n5401, CK => CLK, Q => OUT1_46_port
                           , QN => n4203);
   OUT1_reg_45_inst : DFF_X1 port map( D => n5399, CK => CLK, Q => OUT1_45_port
                           , QN => n4202);
   OUT1_reg_44_inst : DFF_X1 port map( D => n5397, CK => CLK, Q => OUT1_44_port
                           , QN => n4201);
   OUT1_reg_43_inst : DFF_X1 port map( D => n5395, CK => CLK, Q => OUT1_43_port
                           , QN => n4200);
   OUT1_reg_42_inst : DFF_X1 port map( D => n5393, CK => CLK, Q => OUT1_42_port
                           , QN => n4199);
   OUT1_reg_41_inst : DFF_X1 port map( D => n5391, CK => CLK, Q => OUT1_41_port
                           , QN => n4198);
   OUT1_reg_40_inst : DFF_X1 port map( D => n5389, CK => CLK, Q => OUT1_40_port
                           , QN => n4197);
   OUT1_reg_39_inst : DFF_X1 port map( D => n5387, CK => CLK, Q => OUT1_39_port
                           , QN => n4196);
   OUT1_reg_38_inst : DFF_X1 port map( D => n5385, CK => CLK, Q => OUT1_38_port
                           , QN => n4195);
   OUT1_reg_37_inst : DFF_X1 port map( D => n5383, CK => CLK, Q => OUT1_37_port
                           , QN => n4194);
   OUT1_reg_36_inst : DFF_X1 port map( D => n5381, CK => CLK, Q => OUT1_36_port
                           , QN => n4193);
   OUT1_reg_35_inst : DFF_X1 port map( D => n5379, CK => CLK, Q => OUT1_35_port
                           , QN => n4192);
   OUT1_reg_34_inst : DFF_X1 port map( D => n5377, CK => CLK, Q => OUT1_34_port
                           , QN => n4191);
   OUT1_reg_33_inst : DFF_X1 port map( D => n5375, CK => CLK, Q => OUT1_33_port
                           , QN => n4190);
   OUT1_reg_32_inst : DFF_X1 port map( D => n5373, CK => CLK, Q => OUT1_32_port
                           , QN => n4189);
   OUT1_reg_31_inst : DFF_X1 port map( D => n5371, CK => CLK, Q => OUT1_31_port
                           , QN => n4188);
   OUT1_reg_30_inst : DFF_X1 port map( D => n5369, CK => CLK, Q => OUT1_30_port
                           , QN => n4187);
   OUT1_reg_29_inst : DFF_X1 port map( D => n5367, CK => CLK, Q => OUT1_29_port
                           , QN => n4186);
   OUT1_reg_28_inst : DFF_X1 port map( D => n5365, CK => CLK, Q => OUT1_28_port
                           , QN => n4185);
   OUT1_reg_27_inst : DFF_X1 port map( D => n5363, CK => CLK, Q => OUT1_27_port
                           , QN => n4184);
   OUT1_reg_26_inst : DFF_X1 port map( D => n5361, CK => CLK, Q => OUT1_26_port
                           , QN => n4183);
   OUT1_reg_25_inst : DFF_X1 port map( D => n5359, CK => CLK, Q => OUT1_25_port
                           , QN => n4182);
   OUT1_reg_24_inst : DFF_X1 port map( D => n5357, CK => CLK, Q => OUT1_24_port
                           , QN => n4181);
   OUT1_reg_23_inst : DFF_X1 port map( D => n5355, CK => CLK, Q => OUT1_23_port
                           , QN => n4180);
   OUT1_reg_22_inst : DFF_X1 port map( D => n5353, CK => CLK, Q => OUT1_22_port
                           , QN => n4179);
   OUT1_reg_21_inst : DFF_X1 port map( D => n5351, CK => CLK, Q => OUT1_21_port
                           , QN => n4178);
   OUT1_reg_20_inst : DFF_X1 port map( D => n5349, CK => CLK, Q => OUT1_20_port
                           , QN => n4177);
   OUT1_reg_19_inst : DFF_X1 port map( D => n5347, CK => CLK, Q => OUT1_19_port
                           , QN => n4176);
   OUT1_reg_18_inst : DFF_X1 port map( D => n5345, CK => CLK, Q => OUT1_18_port
                           , QN => n4175);
   OUT1_reg_17_inst : DFF_X1 port map( D => n5343, CK => CLK, Q => OUT1_17_port
                           , QN => n4174);
   OUT1_reg_16_inst : DFF_X1 port map( D => n5341, CK => CLK, Q => OUT1_16_port
                           , QN => n4173);
   OUT1_reg_15_inst : DFF_X1 port map( D => n5339, CK => CLK, Q => OUT1_15_port
                           , QN => n4172);
   OUT1_reg_14_inst : DFF_X1 port map( D => n5337, CK => CLK, Q => OUT1_14_port
                           , QN => n4171);
   OUT1_reg_13_inst : DFF_X1 port map( D => n5335, CK => CLK, Q => OUT1_13_port
                           , QN => n4170);
   OUT1_reg_12_inst : DFF_X1 port map( D => n5333, CK => CLK, Q => OUT1_12_port
                           , QN => n4169);
   OUT1_reg_11_inst : DFF_X1 port map( D => n5331, CK => CLK, Q => OUT1_11_port
                           , QN => n4168);
   OUT1_reg_10_inst : DFF_X1 port map( D => n5329, CK => CLK, Q => OUT1_10_port
                           , QN => n4167);
   OUT1_reg_9_inst : DFF_X1 port map( D => n5327, CK => CLK, Q => OUT1_9_port, 
                           QN => n4166);
   OUT1_reg_8_inst : DFF_X1 port map( D => n5325, CK => CLK, Q => OUT1_8_port, 
                           QN => n4165);
   OUT1_reg_7_inst : DFF_X1 port map( D => n5323, CK => CLK, Q => OUT1_7_port, 
                           QN => n4164);
   OUT1_reg_6_inst : DFF_X1 port map( D => n5321, CK => CLK, Q => OUT1_6_port, 
                           QN => n4163);
   OUT1_reg_5_inst : DFF_X1 port map( D => n5319, CK => CLK, Q => OUT1_5_port, 
                           QN => n4162);
   OUT1_reg_4_inst : DFF_X1 port map( D => n5317, CK => CLK, Q => OUT1_4_port, 
                           QN => n4161);
   OUT1_reg_3_inst : DFF_X1 port map( D => n5315, CK => CLK, Q => OUT1_3_port, 
                           QN => n4160);
   OUT1_reg_2_inst : DFF_X1 port map( D => n5313, CK => CLK, Q => OUT1_2_port, 
                           QN => n4159);
   OUT1_reg_1_inst : DFF_X1 port map( D => n5311, CK => CLK, Q => OUT1_1_port, 
                           QN => n4158);
   OUT1_reg_0_inst : DFF_X1 port map( D => n5309, CK => CLK, Q => OUT1_0_port, 
                           QN => n4157);
   OUT2_reg_62_inst : DFF_X1 port map( D => n5307, CK => CLK, Q => OUT2_62_port
                           , QN => n4155);
   OUT2_reg_61_inst : DFF_X1 port map( D => n5306, CK => CLK, Q => OUT2_61_port
                           , QN => n4154);
   OUT2_reg_60_inst : DFF_X1 port map( D => n5305, CK => CLK, Q => OUT2_60_port
                           , QN => n4153);
   OUT2_reg_59_inst : DFF_X1 port map( D => n5304, CK => CLK, Q => OUT2_59_port
                           , QN => n4152);
   OUT2_reg_58_inst : DFF_X1 port map( D => n5303, CK => CLK, Q => OUT2_58_port
                           , QN => n4151);
   OUT2_reg_57_inst : DFF_X1 port map( D => n5302, CK => CLK, Q => OUT2_57_port
                           , QN => n4150);
   OUT2_reg_56_inst : DFF_X1 port map( D => n5301, CK => CLK, Q => OUT2_56_port
                           , QN => n4149);
   OUT2_reg_55_inst : DFF_X1 port map( D => n5300, CK => CLK, Q => OUT2_55_port
                           , QN => n4148);
   OUT2_reg_54_inst : DFF_X1 port map( D => n5299, CK => CLK, Q => OUT2_54_port
                           , QN => n4147);
   OUT2_reg_53_inst : DFF_X1 port map( D => n5298, CK => CLK, Q => OUT2_53_port
                           , QN => n4146);
   OUT2_reg_52_inst : DFF_X1 port map( D => n5297, CK => CLK, Q => OUT2_52_port
                           , QN => n4145);
   OUT2_reg_51_inst : DFF_X1 port map( D => n5296, CK => CLK, Q => OUT2_51_port
                           , QN => n4144);
   OUT2_reg_50_inst : DFF_X1 port map( D => n5295, CK => CLK, Q => OUT2_50_port
                           , QN => n4143);
   OUT2_reg_49_inst : DFF_X1 port map( D => n5294, CK => CLK, Q => OUT2_49_port
                           , QN => n4142);
   OUT2_reg_48_inst : DFF_X1 port map( D => n5293, CK => CLK, Q => OUT2_48_port
                           , QN => n4141);
   OUT2_reg_47_inst : DFF_X1 port map( D => n5292, CK => CLK, Q => OUT2_47_port
                           , QN => n4140);
   OUT2_reg_46_inst : DFF_X1 port map( D => n5291, CK => CLK, Q => OUT2_46_port
                           , QN => n4139);
   OUT2_reg_45_inst : DFF_X1 port map( D => n5290, CK => CLK, Q => OUT2_45_port
                           , QN => n4138);
   OUT2_reg_44_inst : DFF_X1 port map( D => n5289, CK => CLK, Q => OUT2_44_port
                           , QN => n4137);
   OUT2_reg_43_inst : DFF_X1 port map( D => n5288, CK => CLK, Q => OUT2_43_port
                           , QN => n4136);
   OUT2_reg_42_inst : DFF_X1 port map( D => n5287, CK => CLK, Q => OUT2_42_port
                           , QN => n4135);
   OUT2_reg_41_inst : DFF_X1 port map( D => n5286, CK => CLK, Q => OUT2_41_port
                           , QN => n4134);
   OUT2_reg_40_inst : DFF_X1 port map( D => n5285, CK => CLK, Q => OUT2_40_port
                           , QN => n4133);
   OUT2_reg_39_inst : DFF_X1 port map( D => n5284, CK => CLK, Q => OUT2_39_port
                           , QN => n4132);
   OUT2_reg_38_inst : DFF_X1 port map( D => n5283, CK => CLK, Q => OUT2_38_port
                           , QN => n4131);
   OUT2_reg_37_inst : DFF_X1 port map( D => n5282, CK => CLK, Q => OUT2_37_port
                           , QN => n4130);
   OUT2_reg_36_inst : DFF_X1 port map( D => n5281, CK => CLK, Q => OUT2_36_port
                           , QN => n4129);
   OUT2_reg_35_inst : DFF_X1 port map( D => n5280, CK => CLK, Q => OUT2_35_port
                           , QN => n4128);
   OUT2_reg_34_inst : DFF_X1 port map( D => n5279, CK => CLK, Q => OUT2_34_port
                           , QN => n4127);
   OUT2_reg_33_inst : DFF_X1 port map( D => n5278, CK => CLK, Q => OUT2_33_port
                           , QN => n4126);
   OUT2_reg_32_inst : DFF_X1 port map( D => n5277, CK => CLK, Q => OUT2_32_port
                           , QN => n4125);
   OUT2_reg_31_inst : DFF_X1 port map( D => n5276, CK => CLK, Q => OUT2_31_port
                           , QN => n4124);
   OUT2_reg_30_inst : DFF_X1 port map( D => n5275, CK => CLK, Q => OUT2_30_port
                           , QN => n4123);
   OUT2_reg_29_inst : DFF_X1 port map( D => n5274, CK => CLK, Q => OUT2_29_port
                           , QN => n4122);
   OUT2_reg_28_inst : DFF_X1 port map( D => n5273, CK => CLK, Q => OUT2_28_port
                           , QN => n4121);
   OUT2_reg_27_inst : DFF_X1 port map( D => n5272, CK => CLK, Q => OUT2_27_port
                           , QN => n4120);
   OUT2_reg_26_inst : DFF_X1 port map( D => n5271, CK => CLK, Q => OUT2_26_port
                           , QN => n4119);
   OUT2_reg_25_inst : DFF_X1 port map( D => n5270, CK => CLK, Q => OUT2_25_port
                           , QN => n4118);
   OUT2_reg_24_inst : DFF_X1 port map( D => n5269, CK => CLK, Q => OUT2_24_port
                           , QN => n4117);
   OUT2_reg_23_inst : DFF_X1 port map( D => n5268, CK => CLK, Q => OUT2_23_port
                           , QN => n4116);
   OUT2_reg_22_inst : DFF_X1 port map( D => n5267, CK => CLK, Q => OUT2_22_port
                           , QN => n4115);
   OUT2_reg_21_inst : DFF_X1 port map( D => n5266, CK => CLK, Q => OUT2_21_port
                           , QN => n4114);
   OUT2_reg_20_inst : DFF_X1 port map( D => n5265, CK => CLK, Q => OUT2_20_port
                           , QN => n4113);
   OUT2_reg_19_inst : DFF_X1 port map( D => n5264, CK => CLK, Q => OUT2_19_port
                           , QN => n4112);
   OUT2_reg_18_inst : DFF_X1 port map( D => n5263, CK => CLK, Q => OUT2_18_port
                           , QN => n4111);
   OUT2_reg_17_inst : DFF_X1 port map( D => n5262, CK => CLK, Q => OUT2_17_port
                           , QN => n4110);
   OUT2_reg_16_inst : DFF_X1 port map( D => n5261, CK => CLK, Q => OUT2_16_port
                           , QN => n4109);
   OUT2_reg_15_inst : DFF_X1 port map( D => n5260, CK => CLK, Q => OUT2_15_port
                           , QN => n4108);
   OUT2_reg_14_inst : DFF_X1 port map( D => n5259, CK => CLK, Q => OUT2_14_port
                           , QN => n4107);
   OUT2_reg_13_inst : DFF_X1 port map( D => n5258, CK => CLK, Q => OUT2_13_port
                           , QN => n4106);
   OUT2_reg_12_inst : DFF_X1 port map( D => n5257, CK => CLK, Q => OUT2_12_port
                           , QN => n4105);
   OUT2_reg_11_inst : DFF_X1 port map( D => n5256, CK => CLK, Q => OUT2_11_port
                           , QN => n4104);
   OUT2_reg_10_inst : DFF_X1 port map( D => n5255, CK => CLK, Q => OUT2_10_port
                           , QN => n4103);
   OUT2_reg_9_inst : DFF_X1 port map( D => n5254, CK => CLK, Q => OUT2_9_port, 
                           QN => n4102);
   OUT2_reg_8_inst : DFF_X1 port map( D => n5253, CK => CLK, Q => OUT2_8_port, 
                           QN => n4101);
   OUT2_reg_7_inst : DFF_X1 port map( D => n5252, CK => CLK, Q => OUT2_7_port, 
                           QN => n4100);
   OUT2_reg_6_inst : DFF_X1 port map( D => n5251, CK => CLK, Q => OUT2_6_port, 
                           QN => n4099);
   OUT2_reg_5_inst : DFF_X1 port map( D => n5250, CK => CLK, Q => OUT2_5_port, 
                           QN => n4098);
   OUT2_reg_4_inst : DFF_X1 port map( D => n5249, CK => CLK, Q => OUT2_4_port, 
                           QN => n4097);
   OUT2_reg_3_inst : DFF_X1 port map( D => n5248, CK => CLK, Q => OUT2_3_port, 
                           QN => n4096);
   OUT2_reg_2_inst : DFF_X1 port map( D => n5247, CK => CLK, Q => OUT2_2_port, 
                           QN => n4095);
   OUT2_reg_1_inst : DFF_X1 port map( D => n5246, CK => CLK, Q => OUT2_1_port, 
                           QN => n4094);
   OUT2_reg_0_inst : DFF_X1 port map( D => n5245, CK => CLK, Q => OUT2_0_port, 
                           QN => n4093);
   U13039 : NAND3_X1 port map( A1 => n14472, A2 => n14473, A3 => n14474, ZN => 
                           n14070);
   U13040 : NAND3_X1 port map( A1 => n14474, A2 => n14473, A3 => ADD_WR(0), ZN 
                           => n14138);
   U13041 : NAND3_X1 port map( A1 => n14474, A2 => n14472, A3 => ADD_WR(3), ZN 
                           => n14607);
   U13042 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n14474, A3 => ADD_WR(3), 
                           ZN => n14674);
   U13043 : NAND3_X1 port map( A1 => n14472, A2 => n14473, A3 => n15536, ZN => 
                           n15138);
   U13044 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n14473, A3 => n15536, ZN 
                           => n15205);
   U13045 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n14472, A3 => n15536, ZN 
                           => n15669);
   U13046 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => ADD_WR(0), A3 => n15536, 
                           ZN => n15736);
   U13047 : NAND3_X1 port map( A1 => WR, A2 => ENABLE, A3 => n18540, ZN => 
                           n15071);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n7420, CK => CLK, Q => n8575
                           , QN => n13940);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n7419, CK => CLK, Q => n8579
                           , QN => n13943);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n7418, CK => CLK, Q => n8583
                           , QN => n13945);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n7417, CK => CLK, Q => n8587
                           , QN => n13947);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n7292, CK => CLK, Q => 
                           n18551, QN => n14140);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n7291, CK => CLK, Q => 
                           n18571, QN => n14142);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n7290, CK => CLK, Q => 
                           n18591, QN => n14143);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n7289, CK => CLK, Q => 
                           n18611, QN => n14144);
   REGISTERS_reg_6_63_inst : DFF_X1 port map( D => n7036, CK => CLK, Q => 
                           n18555, QN => n14406);
   REGISTERS_reg_6_62_inst : DFF_X1 port map( D => n7035, CK => CLK, Q => 
                           n18575, QN => n14408);
   REGISTERS_reg_6_61_inst : DFF_X1 port map( D => n7034, CK => CLK, Q => 
                           n18595, QN => n14409);
   REGISTERS_reg_6_60_inst : DFF_X1 port map( D => n7033, CK => CLK, Q => 
                           n18615, QN => n14410);
   REGISTERS_reg_4_63_inst : DFF_X1 port map( D => n7164, CK => CLK, Q => 
                           n18545, QN => n14273);
   REGISTERS_reg_4_62_inst : DFF_X1 port map( D => n7163, CK => CLK, Q => 
                           n18565, QN => n14275);
   REGISTERS_reg_4_61_inst : DFF_X1 port map( D => n7162, CK => CLK, Q => 
                           n18585, QN => n14276);
   REGISTERS_reg_4_60_inst : DFF_X1 port map( D => n7161, CK => CLK, Q => 
                           n18605, QN => n14277);
   REGISTERS_reg_5_63_inst : DFF_X1 port map( D => n7100, CK => CLK, Q => 
                           n20717, QN => n14340);
   REGISTERS_reg_5_62_inst : DFF_X1 port map( D => n7099, CK => CLK, Q => 
                           n20716, QN => n14342);
   REGISTERS_reg_5_61_inst : DFF_X1 port map( D => n7098, CK => CLK, Q => 
                           n20715, QN => n14343);
   REGISTERS_reg_5_60_inst : DFF_X1 port map( D => n7097, CK => CLK, Q => 
                           n20714, QN => n14344);
   REGISTERS_reg_7_63_inst : DFF_X1 port map( D => n6972, CK => CLK, Q => 
                           n20713, QN => n14476);
   REGISTERS_reg_7_62_inst : DFF_X1 port map( D => n6971, CK => CLK, Q => 
                           n20712, QN => n14478);
   REGISTERS_reg_7_61_inst : DFF_X1 port map( D => n6970, CK => CLK, Q => 
                           n20711, QN => n14479);
   REGISTERS_reg_7_60_inst : DFF_X1 port map( D => n6969, CK => CLK, Q => 
                           n20710, QN => n14480);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n7228, CK => CLK, Q => 
                           n20709, QN => n14207);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n7227, CK => CLK, Q => 
                           n20708, QN => n14209);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n7226, CK => CLK, Q => 
                           n20707, QN => n14210);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n7225, CK => CLK, Q => 
                           n20706, QN => n14211);
   REGISTERS_reg_10_63_inst : DFF_X1 port map( D => n6780, CK => CLK, Q => 
                           n18559, QN => n14676);
   REGISTERS_reg_10_62_inst : DFF_X1 port map( D => n6779, CK => CLK, Q => 
                           n18579, QN => n14678);
   REGISTERS_reg_10_61_inst : DFF_X1 port map( D => n6778, CK => CLK, Q => 
                           n18599, QN => n14679);
   REGISTERS_reg_10_60_inst : DFF_X1 port map( D => n6777, CK => CLK, Q => 
                           n18619, QN => n14680);
   REGISTERS_reg_8_63_inst : DFF_X1 port map( D => n6908, CK => CLK, Q => n8960
                           , QN => n14542);
   REGISTERS_reg_8_62_inst : DFF_X1 port map( D => n6907, CK => CLK, Q => n8964
                           , QN => n14544);
   REGISTERS_reg_8_61_inst : DFF_X1 port map( D => n6906, CK => CLK, Q => n8968
                           , QN => n14545);
   REGISTERS_reg_8_60_inst : DFF_X1 port map( D => n6905, CK => CLK, Q => n8972
                           , QN => n14546);
   REGISTERS_reg_14_63_inst : DFF_X1 port map( D => n6524, CK => CLK, Q => 
                           n20705, QN => n14940);
   REGISTERS_reg_14_62_inst : DFF_X1 port map( D => n6523, CK => CLK, Q => 
                           n20704, QN => n14942);
   REGISTERS_reg_14_61_inst : DFF_X1 port map( D => n6522, CK => CLK, Q => 
                           n20703, QN => n14943);
   REGISTERS_reg_14_60_inst : DFF_X1 port map( D => n6521, CK => CLK, Q => 
                           n20702, QN => n14944);
   REGISTERS_reg_12_63_inst : DFF_X1 port map( D => n6652, CK => CLK, Q => 
                           n20701, QN => n14808);
   REGISTERS_reg_12_62_inst : DFF_X1 port map( D => n6651, CK => CLK, Q => 
                           n20700, QN => n14810);
   REGISTERS_reg_12_61_inst : DFF_X1 port map( D => n6650, CK => CLK, Q => 
                           n20699, QN => n14811);
   REGISTERS_reg_12_60_inst : DFF_X1 port map( D => n6649, CK => CLK, Q => 
                           n20698, QN => n14812);
   REGISTERS_reg_11_63_inst : DFF_X1 port map( D => n6716, CK => CLK, Q => 
                           n20697, QN => n14742);
   REGISTERS_reg_11_62_inst : DFF_X1 port map( D => n6715, CK => CLK, Q => 
                           n20696, QN => n14744);
   REGISTERS_reg_11_61_inst : DFF_X1 port map( D => n6714, CK => CLK, Q => 
                           n20695, QN => n14745);
   REGISTERS_reg_11_60_inst : DFF_X1 port map( D => n6713, CK => CLK, Q => 
                           n20694, QN => n14746);
   REGISTERS_reg_9_63_inst : DFF_X1 port map( D => n6844, CK => CLK, Q => n8959
                           , QN => n14609);
   REGISTERS_reg_9_62_inst : DFF_X1 port map( D => n6843, CK => CLK, Q => n8963
                           , QN => n14611);
   REGISTERS_reg_9_61_inst : DFF_X1 port map( D => n6842, CK => CLK, Q => n8967
                           , QN => n14612);
   REGISTERS_reg_9_60_inst : DFF_X1 port map( D => n6841, CK => CLK, Q => n8971
                           , QN => n14613);
   REGISTERS_reg_15_63_inst : DFF_X1 port map( D => n6460, CK => CLK, Q => 
                           n20693, QN => n15006);
   REGISTERS_reg_15_62_inst : DFF_X1 port map( D => n6459, CK => CLK, Q => 
                           n20692, QN => n15008);
   REGISTERS_reg_15_61_inst : DFF_X1 port map( D => n6458, CK => CLK, Q => 
                           n20691, QN => n15009);
   REGISTERS_reg_15_60_inst : DFF_X1 port map( D => n6457, CK => CLK, Q => 
                           n20690, QN => n15010);
   REGISTERS_reg_13_63_inst : DFF_X1 port map( D => n6588, CK => CLK, Q => 
                           n8576, QN => n14874);
   REGISTERS_reg_13_62_inst : DFF_X1 port map( D => n6587, CK => CLK, Q => 
                           n8580, QN => n14876);
   REGISTERS_reg_13_61_inst : DFF_X1 port map( D => n6586, CK => CLK, Q => 
                           n8584, QN => n14877);
   REGISTERS_reg_13_60_inst : DFF_X1 port map( D => n6585, CK => CLK, Q => 
                           n8588, QN => n14878);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n7356, CK => CLK, Q => 
                           n20689, QN => n14073);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n7355, CK => CLK, Q => 
                           n20688, QN => n14075);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n7354, CK => CLK, Q => 
                           n20687, QN => n14076);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n7353, CK => CLK, Q => 
                           n20686, QN => n14077);
   REGISTERS_reg_30_63_inst : DFF_X1 port map( D => n5500, CK => CLK, Q => 
                           n20685, QN => n16004);
   REGISTERS_reg_30_62_inst : DFF_X1 port map( D => n5499, CK => CLK, Q => 
                           n20684, QN => n16006);
   REGISTERS_reg_30_61_inst : DFF_X1 port map( D => n5498, CK => CLK, Q => 
                           n20683, QN => n16007);
   REGISTERS_reg_30_60_inst : DFF_X1 port map( D => n5497, CK => CLK, Q => 
                           n20682, QN => n16008);
   REGISTERS_reg_29_63_inst : DFF_X1 port map( D => n5564, CK => CLK, Q => 
                           n18548, QN => n15938);
   REGISTERS_reg_29_62_inst : DFF_X1 port map( D => n5563, CK => CLK, Q => 
                           n18568, QN => n15940);
   REGISTERS_reg_29_61_inst : DFF_X1 port map( D => n5562, CK => CLK, Q => 
                           n18588, QN => n15941);
   REGISTERS_reg_29_60_inst : DFF_X1 port map( D => n5561, CK => CLK, Q => 
                           n18608, QN => n15942);
   REGISTERS_reg_28_63_inst : DFF_X1 port map( D => n5628, CK => CLK, Q => 
                           n20681, QN => n15872);
   REGISTERS_reg_28_62_inst : DFF_X1 port map( D => n5627, CK => CLK, Q => 
                           n20680, QN => n15874);
   REGISTERS_reg_28_61_inst : DFF_X1 port map( D => n5626, CK => CLK, Q => 
                           n20679, QN => n15875);
   REGISTERS_reg_28_60_inst : DFF_X1 port map( D => n5625, CK => CLK, Q => 
                           n20678, QN => n15876);
   REGISTERS_reg_27_63_inst : DFF_X1 port map( D => n5692, CK => CLK, Q => 
                           n18550, QN => n15806);
   REGISTERS_reg_27_62_inst : DFF_X1 port map( D => n5691, CK => CLK, Q => 
                           n18570, QN => n15808);
   REGISTERS_reg_27_61_inst : DFF_X1 port map( D => n5690, CK => CLK, Q => 
                           n18590, QN => n15809);
   REGISTERS_reg_27_60_inst : DFF_X1 port map( D => n5689, CK => CLK, Q => 
                           n18610, QN => n15810);
   REGISTERS_reg_26_63_inst : DFF_X1 port map( D => n5756, CK => CLK, Q => 
                           n20677, QN => n15740);
   REGISTERS_reg_26_62_inst : DFF_X1 port map( D => n5755, CK => CLK, Q => 
                           n20676, QN => n15742);
   REGISTERS_reg_26_61_inst : DFF_X1 port map( D => n5754, CK => CLK, Q => 
                           n20675, QN => n15743);
   REGISTERS_reg_26_60_inst : DFF_X1 port map( D => n5753, CK => CLK, Q => 
                           n20674, QN => n15744);
   REGISTERS_reg_25_63_inst : DFF_X1 port map( D => n5820, CK => CLK, Q => 
                           n8957, QN => n15671);
   REGISTERS_reg_25_62_inst : DFF_X1 port map( D => n5819, CK => CLK, Q => 
                           n8961, QN => n15673);
   REGISTERS_reg_25_61_inst : DFF_X1 port map( D => n5818, CK => CLK, Q => 
                           n8965, QN => n15674);
   REGISTERS_reg_25_60_inst : DFF_X1 port map( D => n5817, CK => CLK, Q => 
                           n8969, QN => n15675);
   REGISTERS_reg_31_63_inst : DFF_X1 port map( D => n5436, CK => CLK, Q => 
                           n18544, QN => n16070);
   REGISTERS_reg_31_62_inst : DFF_X1 port map( D => n5434, CK => CLK, Q => 
                           n18564, QN => n16124);
   REGISTERS_reg_31_61_inst : DFF_X1 port map( D => n5432, CK => CLK, Q => 
                           n18584, QN => n16143);
   REGISTERS_reg_31_60_inst : DFF_X1 port map( D => n5430, CK => CLK, Q => 
                           n18604, QN => n16162);
   REGISTERS_reg_23_63_inst : DFF_X1 port map( D => n5948, CK => CLK, Q => 
                           n8829, QN => n15538);
   REGISTERS_reg_23_62_inst : DFF_X1 port map( D => n5947, CK => CLK, Q => 
                           n8831, QN => n15540);
   REGISTERS_reg_23_61_inst : DFF_X1 port map( D => n5946, CK => CLK, Q => 
                           n8833, QN => n15541);
   REGISTERS_reg_23_60_inst : DFF_X1 port map( D => n5945, CK => CLK, Q => 
                           n8835, QN => n15542);
   REGISTERS_reg_22_63_inst : DFF_X1 port map( D => n6012, CK => CLK, Q => 
                           n18549, QN => n15471);
   REGISTERS_reg_22_62_inst : DFF_X1 port map( D => n6011, CK => CLK, Q => 
                           n18569, QN => n15473);
   REGISTERS_reg_22_61_inst : DFF_X1 port map( D => n6010, CK => CLK, Q => 
                           n18589, QN => n15474);
   REGISTERS_reg_22_60_inst : DFF_X1 port map( D => n6009, CK => CLK, Q => 
                           n18609, QN => n15475);
   REGISTERS_reg_21_63_inst : DFF_X1 port map( D => n6076, CK => CLK, Q => 
                           n20673, QN => n15405);
   REGISTERS_reg_21_62_inst : DFF_X1 port map( D => n6075, CK => CLK, Q => 
                           n20672, QN => n15407);
   REGISTERS_reg_21_61_inst : DFF_X1 port map( D => n6074, CK => CLK, Q => 
                           n20671, QN => n15408);
   REGISTERS_reg_21_60_inst : DFF_X1 port map( D => n6073, CK => CLK, Q => 
                           n20670, QN => n15409);
   REGISTERS_reg_20_63_inst : DFF_X1 port map( D => n6140, CK => CLK, Q => 
                           n18541, QN => n15339);
   REGISTERS_reg_20_62_inst : DFF_X1 port map( D => n6139, CK => CLK, Q => 
                           n18561, QN => n15341);
   REGISTERS_reg_20_61_inst : DFF_X1 port map( D => n6138, CK => CLK, Q => 
                           n18581, QN => n15342);
   REGISTERS_reg_20_60_inst : DFF_X1 port map( D => n6137, CK => CLK, Q => 
                           n18601, QN => n15343);
   REGISTERS_reg_19_63_inst : DFF_X1 port map( D => n6204, CK => CLK, Q => 
                           n20669, QN => n15273);
   REGISTERS_reg_19_62_inst : DFF_X1 port map( D => n6203, CK => CLK, Q => 
                           n20668, QN => n15275);
   REGISTERS_reg_19_61_inst : DFF_X1 port map( D => n6202, CK => CLK, Q => 
                           n20667, QN => n15276);
   REGISTERS_reg_19_60_inst : DFF_X1 port map( D => n6201, CK => CLK, Q => 
                           n20666, QN => n15277);
   REGISTERS_reg_18_63_inst : DFF_X1 port map( D => n6268, CK => CLK, Q => 
                           n8830, QN => n15207);
   REGISTERS_reg_18_62_inst : DFF_X1 port map( D => n6267, CK => CLK, Q => 
                           n8832, QN => n15209);
   REGISTERS_reg_18_61_inst : DFF_X1 port map( D => n6266, CK => CLK, Q => 
                           n8834, QN => n15210);
   REGISTERS_reg_18_60_inst : DFF_X1 port map( D => n6265, CK => CLK, Q => 
                           n8836, QN => n15211);
   REGISTERS_reg_24_63_inst : DFF_X1 port map( D => n5884, CK => CLK, Q => 
                           n20665, QN => n15604);
   REGISTERS_reg_24_62_inst : DFF_X1 port map( D => n5883, CK => CLK, Q => 
                           n20664, QN => n15606);
   REGISTERS_reg_24_61_inst : DFF_X1 port map( D => n5882, CK => CLK, Q => 
                           n20663, QN => n15607);
   REGISTERS_reg_24_60_inst : DFF_X1 port map( D => n5881, CK => CLK, Q => 
                           n20662, QN => n15608);
   REGISTERS_reg_17_63_inst : DFF_X1 port map( D => n6332, CK => CLK, Q => 
                           n18554, QN => n15140);
   REGISTERS_reg_17_62_inst : DFF_X1 port map( D => n6331, CK => CLK, Q => 
                           n18574, QN => n15142);
   REGISTERS_reg_17_61_inst : DFF_X1 port map( D => n6330, CK => CLK, Q => 
                           n18594, QN => n15143);
   REGISTERS_reg_17_60_inst : DFF_X1 port map( D => n6329, CK => CLK, Q => 
                           n18614, QN => n15144);
   REGISTERS_reg_16_63_inst : DFF_X1 port map( D => n6396, CK => CLK, Q => 
                           n8573, QN => n15073);
   REGISTERS_reg_16_62_inst : DFF_X1 port map( D => n6395, CK => CLK, Q => 
                           n8577, QN => n15075);
   REGISTERS_reg_16_61_inst : DFF_X1 port map( D => n6394, CK => CLK, Q => 
                           n8581, QN => n15076);
   REGISTERS_reg_16_60_inst : DFF_X1 port map( D => n6393, CK => CLK, Q => 
                           n8585, QN => n15077);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n7416, CK => CLK, Q => n8591
                           , QN => n13949);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n7415, CK => CLK, Q => n8595
                           , QN => n13951);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n7414, CK => CLK, Q => n8599
                           , QN => n13953);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n7413, CK => CLK, Q => n8603
                           , QN => n13955);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n7412, CK => CLK, Q => n8607
                           , QN => n13957);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n7411, CK => CLK, Q => n8611
                           , QN => n13959);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n7410, CK => CLK, Q => n8615
                           , QN => n13961);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n7409, CK => CLK, Q => n8619
                           , QN => n13963);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n7408, CK => CLK, Q => n8623
                           , QN => n13965);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n7407, CK => CLK, Q => n8627
                           , QN => n13967);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n7406, CK => CLK, Q => n8631
                           , QN => n13969);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n7405, CK => CLK, Q => n8635
                           , QN => n13971);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n7404, CK => CLK, Q => n8639
                           , QN => n13973);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n7403, CK => CLK, Q => n8643
                           , QN => n13975);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n7402, CK => CLK, Q => n8647
                           , QN => n13977);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n7401, CK => CLK, Q => n8651
                           , QN => n13979);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n7400, CK => CLK, Q => n8655
                           , QN => n13981);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n7399, CK => CLK, Q => n8659
                           , QN => n13983);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n7398, CK => CLK, Q => n8663
                           , QN => n13985);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n7397, CK => CLK, Q => n8667
                           , QN => n13987);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n7396, CK => CLK, Q => n8671
                           , QN => n13989);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n7395, CK => CLK, Q => n8675
                           , QN => n13991);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n7394, CK => CLK, Q => n8679
                           , QN => n13993);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n7393, CK => CLK, Q => n8683
                           , QN => n13995);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n7392, CK => CLK, Q => n8687
                           , QN => n13997);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n7391, CK => CLK, Q => n8691
                           , QN => n13999);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n7390, CK => CLK, Q => n8695
                           , QN => n14001);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n7389, CK => CLK, Q => n8699
                           , QN => n14003);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n7388, CK => CLK, Q => n8703
                           , QN => n14005);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n7387, CK => CLK, Q => n8707
                           , QN => n14007);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n7386, CK => CLK, Q => n8711
                           , QN => n14009);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n7385, CK => CLK, Q => n8715
                           , QN => n14011);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n7384, CK => CLK, Q => n8719
                           , QN => n14013);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n7383, CK => CLK, Q => n8723
                           , QN => n14015);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n7382, CK => CLK, Q => n8727
                           , QN => n14017);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n7381, CK => CLK, Q => n8731
                           , QN => n14019);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n7380, CK => CLK, Q => n8735
                           , QN => n14021);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n7379, CK => CLK, Q => n8739
                           , QN => n14023);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n7378, CK => CLK, Q => n8743
                           , QN => n14025);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n7377, CK => CLK, Q => n8747
                           , QN => n14027);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n7376, CK => CLK, Q => n8751
                           , QN => n14029);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n7375, CK => CLK, Q => n8755
                           , QN => n14031);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n7374, CK => CLK, Q => n8759
                           , QN => n14033);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n7373, CK => CLK, Q => n8763
                           , QN => n14035);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n7372, CK => CLK, Q => n8767
                           , QN => n14037);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n7371, CK => CLK, Q => n8771
                           , QN => n14039);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n7370, CK => CLK, Q => n8775
                           , QN => n14041);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n7369, CK => CLK, Q => n8779
                           , QN => n14043);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n7368, CK => CLK, Q => n8783
                           , QN => n14045);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n7367, CK => CLK, Q => n8787
                           , QN => n14047);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n7366, CK => CLK, Q => n8791,
                           QN => n14049);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n7365, CK => CLK, Q => n8795,
                           QN => n14051);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n7364, CK => CLK, Q => n8799,
                           QN => n14053);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n7363, CK => CLK, Q => n8803,
                           QN => n14055);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n7362, CK => CLK, Q => n8807,
                           QN => n14057);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n7361, CK => CLK, Q => n8811,
                           QN => n14059);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n7360, CK => CLK, Q => n8815,
                           QN => n14061);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n7359, CK => CLK, Q => n8819,
                           QN => n14063);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n7358, CK => CLK, Q => n8823,
                           QN => n14065);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n7357, CK => CLK, Q => n8827,
                           QN => n14067);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n7288, CK => CLK, Q => 
                           n18631, QN => n14145);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n7287, CK => CLK, Q => 
                           n18651, QN => n14146);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n7286, CK => CLK, Q => 
                           n18671, QN => n14147);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n7285, CK => CLK, Q => 
                           n18691, QN => n14148);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n7284, CK => CLK, Q => 
                           n18711, QN => n14149);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n7283, CK => CLK, Q => 
                           n18731, QN => n14150);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n7282, CK => CLK, Q => 
                           n18751, QN => n14151);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n7281, CK => CLK, Q => 
                           n18771, QN => n14152);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n7280, CK => CLK, Q => 
                           n18791, QN => n14153);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n7279, CK => CLK, Q => 
                           n18811, QN => n14154);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n7278, CK => CLK, Q => 
                           n18831, QN => n14155);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n7277, CK => CLK, Q => 
                           n18851, QN => n14156);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n7276, CK => CLK, Q => 
                           n18871, QN => n14157);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n7275, CK => CLK, Q => 
                           n18891, QN => n14158);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n7274, CK => CLK, Q => 
                           n18911, QN => n14159);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n7273, CK => CLK, Q => 
                           n18931, QN => n14160);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n7272, CK => CLK, Q => 
                           n18951, QN => n14161);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n7271, CK => CLK, Q => 
                           n18971, QN => n14162);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n7270, CK => CLK, Q => 
                           n18991, QN => n14163);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n7269, CK => CLK, Q => 
                           n19011, QN => n14164);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n7268, CK => CLK, Q => 
                           n19031, QN => n14165);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n7267, CK => CLK, Q => 
                           n19051, QN => n14166);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n7266, CK => CLK, Q => 
                           n19071, QN => n14167);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n7265, CK => CLK, Q => 
                           n19091, QN => n14168);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n7264, CK => CLK, Q => 
                           n19111, QN => n14169);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n7263, CK => CLK, Q => 
                           n19131, QN => n14170);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n7262, CK => CLK, Q => 
                           n19151, QN => n14171);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n7261, CK => CLK, Q => 
                           n19171, QN => n14172);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n7260, CK => CLK, Q => 
                           n19191, QN => n14173);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n7259, CK => CLK, Q => 
                           n19211, QN => n14174);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n7258, CK => CLK, Q => 
                           n19231, QN => n14175);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n7257, CK => CLK, Q => 
                           n19251, QN => n14176);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n7256, CK => CLK, Q => 
                           n19271, QN => n14177);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n7255, CK => CLK, Q => 
                           n19291, QN => n14178);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n7254, CK => CLK, Q => 
                           n19311, QN => n14179);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n7253, CK => CLK, Q => 
                           n19331, QN => n14180);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n7252, CK => CLK, Q => 
                           n19351, QN => n14181);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n7251, CK => CLK, Q => 
                           n19371, QN => n14182);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n7250, CK => CLK, Q => 
                           n19391, QN => n14183);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n7249, CK => CLK, Q => 
                           n19411, QN => n14184);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n7248, CK => CLK, Q => 
                           n19431, QN => n14185);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n7247, CK => CLK, Q => 
                           n19451, QN => n14186);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n7246, CK => CLK, Q => 
                           n19471, QN => n14187);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n7245, CK => CLK, Q => 
                           n19491, QN => n14188);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n7244, CK => CLK, Q => 
                           n19511, QN => n14189);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n7243, CK => CLK, Q => 
                           n19531, QN => n14190);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n7242, CK => CLK, Q => 
                           n19551, QN => n14191);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n7241, CK => CLK, Q => 
                           n19571, QN => n14192);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n7240, CK => CLK, Q => 
                           n19591, QN => n14193);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n7239, CK => CLK, Q => 
                           n19611, QN => n14194);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n7238, CK => CLK, Q => n19631
                           , QN => n14195);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n7237, CK => CLK, Q => n19651
                           , QN => n14196);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n7236, CK => CLK, Q => n19671
                           , QN => n14197);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n7235, CK => CLK, Q => n19691
                           , QN => n14198);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n7234, CK => CLK, Q => n19711
                           , QN => n14199);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n7233, CK => CLK, Q => n19731
                           , QN => n14200);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n7232, CK => CLK, Q => n19751
                           , QN => n14201);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n7231, CK => CLK, Q => n19771
                           , QN => n14202);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n7230, CK => CLK, Q => n19791
                           , QN => n14203);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n7229, CK => CLK, Q => n19811
                           , QN => n14204);
   REGISTERS_reg_6_59_inst : DFF_X1 port map( D => n7032, CK => CLK, Q => 
                           n18635, QN => n14411);
   REGISTERS_reg_6_58_inst : DFF_X1 port map( D => n7031, CK => CLK, Q => 
                           n18655, QN => n14412);
   REGISTERS_reg_6_57_inst : DFF_X1 port map( D => n7030, CK => CLK, Q => 
                           n18675, QN => n14413);
   REGISTERS_reg_6_56_inst : DFF_X1 port map( D => n7029, CK => CLK, Q => 
                           n18695, QN => n14414);
   REGISTERS_reg_6_55_inst : DFF_X1 port map( D => n7028, CK => CLK, Q => 
                           n18715, QN => n14415);
   REGISTERS_reg_6_54_inst : DFF_X1 port map( D => n7027, CK => CLK, Q => 
                           n18735, QN => n14416);
   REGISTERS_reg_6_53_inst : DFF_X1 port map( D => n7026, CK => CLK, Q => 
                           n18755, QN => n14417);
   REGISTERS_reg_6_52_inst : DFF_X1 port map( D => n7025, CK => CLK, Q => 
                           n18775, QN => n14418);
   REGISTERS_reg_6_51_inst : DFF_X1 port map( D => n7024, CK => CLK, Q => 
                           n18795, QN => n14419);
   REGISTERS_reg_6_50_inst : DFF_X1 port map( D => n7023, CK => CLK, Q => 
                           n18815, QN => n14420);
   REGISTERS_reg_6_49_inst : DFF_X1 port map( D => n7022, CK => CLK, Q => 
                           n18835, QN => n14421);
   REGISTERS_reg_6_48_inst : DFF_X1 port map( D => n7021, CK => CLK, Q => 
                           n18855, QN => n14422);
   REGISTERS_reg_6_47_inst : DFF_X1 port map( D => n7020, CK => CLK, Q => 
                           n18875, QN => n14423);
   REGISTERS_reg_6_46_inst : DFF_X1 port map( D => n7019, CK => CLK, Q => 
                           n18895, QN => n14424);
   REGISTERS_reg_6_45_inst : DFF_X1 port map( D => n7018, CK => CLK, Q => 
                           n18915, QN => n14425);
   REGISTERS_reg_6_44_inst : DFF_X1 port map( D => n7017, CK => CLK, Q => 
                           n18935, QN => n14426);
   REGISTERS_reg_6_43_inst : DFF_X1 port map( D => n7016, CK => CLK, Q => 
                           n18955, QN => n14427);
   REGISTERS_reg_6_42_inst : DFF_X1 port map( D => n7015, CK => CLK, Q => 
                           n18975, QN => n14428);
   REGISTERS_reg_6_41_inst : DFF_X1 port map( D => n7014, CK => CLK, Q => 
                           n18995, QN => n14429);
   REGISTERS_reg_6_40_inst : DFF_X1 port map( D => n7013, CK => CLK, Q => 
                           n19015, QN => n14430);
   REGISTERS_reg_6_39_inst : DFF_X1 port map( D => n7012, CK => CLK, Q => 
                           n19035, QN => n14431);
   REGISTERS_reg_6_38_inst : DFF_X1 port map( D => n7011, CK => CLK, Q => 
                           n19055, QN => n14432);
   REGISTERS_reg_6_37_inst : DFF_X1 port map( D => n7010, CK => CLK, Q => 
                           n19075, QN => n14433);
   REGISTERS_reg_6_36_inst : DFF_X1 port map( D => n7009, CK => CLK, Q => 
                           n19095, QN => n14434);
   REGISTERS_reg_6_35_inst : DFF_X1 port map( D => n7008, CK => CLK, Q => 
                           n19115, QN => n14435);
   REGISTERS_reg_6_34_inst : DFF_X1 port map( D => n7007, CK => CLK, Q => 
                           n19135, QN => n14436);
   REGISTERS_reg_6_33_inst : DFF_X1 port map( D => n7006, CK => CLK, Q => 
                           n19155, QN => n14437);
   REGISTERS_reg_6_32_inst : DFF_X1 port map( D => n7005, CK => CLK, Q => 
                           n19175, QN => n14438);
   REGISTERS_reg_6_31_inst : DFF_X1 port map( D => n7004, CK => CLK, Q => 
                           n19195, QN => n14439);
   REGISTERS_reg_6_30_inst : DFF_X1 port map( D => n7003, CK => CLK, Q => 
                           n19215, QN => n14440);
   REGISTERS_reg_6_29_inst : DFF_X1 port map( D => n7002, CK => CLK, Q => 
                           n19235, QN => n14441);
   REGISTERS_reg_6_28_inst : DFF_X1 port map( D => n7001, CK => CLK, Q => 
                           n19255, QN => n14442);
   REGISTERS_reg_6_27_inst : DFF_X1 port map( D => n7000, CK => CLK, Q => 
                           n19275, QN => n14443);
   REGISTERS_reg_6_26_inst : DFF_X1 port map( D => n6999, CK => CLK, Q => 
                           n19295, QN => n14444);
   REGISTERS_reg_6_25_inst : DFF_X1 port map( D => n6998, CK => CLK, Q => 
                           n19315, QN => n14445);
   REGISTERS_reg_6_24_inst : DFF_X1 port map( D => n6997, CK => CLK, Q => 
                           n19335, QN => n14446);
   REGISTERS_reg_6_23_inst : DFF_X1 port map( D => n6996, CK => CLK, Q => 
                           n19355, QN => n14447);
   REGISTERS_reg_6_22_inst : DFF_X1 port map( D => n6995, CK => CLK, Q => 
                           n19375, QN => n14448);
   REGISTERS_reg_6_21_inst : DFF_X1 port map( D => n6994, CK => CLK, Q => 
                           n19395, QN => n14449);
   REGISTERS_reg_6_20_inst : DFF_X1 port map( D => n6993, CK => CLK, Q => 
                           n19415, QN => n14450);
   REGISTERS_reg_6_19_inst : DFF_X1 port map( D => n6992, CK => CLK, Q => 
                           n19435, QN => n14451);
   REGISTERS_reg_6_18_inst : DFF_X1 port map( D => n6991, CK => CLK, Q => 
                           n19455, QN => n14452);
   REGISTERS_reg_6_17_inst : DFF_X1 port map( D => n6990, CK => CLK, Q => 
                           n19475, QN => n14453);
   REGISTERS_reg_6_16_inst : DFF_X1 port map( D => n6989, CK => CLK, Q => 
                           n19495, QN => n14454);
   REGISTERS_reg_6_15_inst : DFF_X1 port map( D => n6988, CK => CLK, Q => 
                           n19515, QN => n14455);
   REGISTERS_reg_6_14_inst : DFF_X1 port map( D => n6987, CK => CLK, Q => 
                           n19535, QN => n14456);
   REGISTERS_reg_6_13_inst : DFF_X1 port map( D => n6986, CK => CLK, Q => 
                           n19555, QN => n14457);
   REGISTERS_reg_6_12_inst : DFF_X1 port map( D => n6985, CK => CLK, Q => 
                           n19575, QN => n14458);
   REGISTERS_reg_6_11_inst : DFF_X1 port map( D => n6984, CK => CLK, Q => 
                           n19595, QN => n14459);
   REGISTERS_reg_6_10_inst : DFF_X1 port map( D => n6983, CK => CLK, Q => 
                           n19615, QN => n14460);
   REGISTERS_reg_6_9_inst : DFF_X1 port map( D => n6982, CK => CLK, Q => n19635
                           , QN => n14461);
   REGISTERS_reg_6_8_inst : DFF_X1 port map( D => n6981, CK => CLK, Q => n19655
                           , QN => n14462);
   REGISTERS_reg_6_7_inst : DFF_X1 port map( D => n6980, CK => CLK, Q => n19675
                           , QN => n14463);
   REGISTERS_reg_6_6_inst : DFF_X1 port map( D => n6979, CK => CLK, Q => n19695
                           , QN => n14464);
   REGISTERS_reg_6_5_inst : DFF_X1 port map( D => n6978, CK => CLK, Q => n19715
                           , QN => n14465);
   REGISTERS_reg_6_4_inst : DFF_X1 port map( D => n6977, CK => CLK, Q => n19735
                           , QN => n14466);
   REGISTERS_reg_6_3_inst : DFF_X1 port map( D => n6976, CK => CLK, Q => n19755
                           , QN => n14467);
   REGISTERS_reg_6_2_inst : DFF_X1 port map( D => n6975, CK => CLK, Q => n19775
                           , QN => n14468);
   REGISTERS_reg_6_1_inst : DFF_X1 port map( D => n6974, CK => CLK, Q => n19795
                           , QN => n14469);
   REGISTERS_reg_6_0_inst : DFF_X1 port map( D => n6973, CK => CLK, Q => n19815
                           , QN => n14470);
   REGISTERS_reg_4_59_inst : DFF_X1 port map( D => n7160, CK => CLK, Q => 
                           n18625, QN => n14278);
   REGISTERS_reg_4_58_inst : DFF_X1 port map( D => n7159, CK => CLK, Q => 
                           n18645, QN => n14279);
   REGISTERS_reg_4_57_inst : DFF_X1 port map( D => n7158, CK => CLK, Q => 
                           n18665, QN => n14280);
   REGISTERS_reg_4_56_inst : DFF_X1 port map( D => n7157, CK => CLK, Q => 
                           n18685, QN => n14281);
   REGISTERS_reg_4_55_inst : DFF_X1 port map( D => n7156, CK => CLK, Q => 
                           n18705, QN => n14282);
   REGISTERS_reg_4_54_inst : DFF_X1 port map( D => n7155, CK => CLK, Q => 
                           n18725, QN => n14283);
   REGISTERS_reg_4_53_inst : DFF_X1 port map( D => n7154, CK => CLK, Q => 
                           n18745, QN => n14284);
   REGISTERS_reg_4_52_inst : DFF_X1 port map( D => n7153, CK => CLK, Q => 
                           n18765, QN => n14285);
   REGISTERS_reg_4_51_inst : DFF_X1 port map( D => n7152, CK => CLK, Q => 
                           n18785, QN => n14286);
   REGISTERS_reg_4_50_inst : DFF_X1 port map( D => n7151, CK => CLK, Q => 
                           n18805, QN => n14287);
   REGISTERS_reg_4_49_inst : DFF_X1 port map( D => n7150, CK => CLK, Q => 
                           n18825, QN => n14288);
   REGISTERS_reg_4_48_inst : DFF_X1 port map( D => n7149, CK => CLK, Q => 
                           n18845, QN => n14289);
   REGISTERS_reg_4_47_inst : DFF_X1 port map( D => n7148, CK => CLK, Q => 
                           n18865, QN => n14290);
   REGISTERS_reg_4_46_inst : DFF_X1 port map( D => n7147, CK => CLK, Q => 
                           n18885, QN => n14291);
   REGISTERS_reg_4_45_inst : DFF_X1 port map( D => n7146, CK => CLK, Q => 
                           n18905, QN => n14292);
   REGISTERS_reg_4_44_inst : DFF_X1 port map( D => n7145, CK => CLK, Q => 
                           n18925, QN => n14293);
   REGISTERS_reg_4_43_inst : DFF_X1 port map( D => n7144, CK => CLK, Q => 
                           n18945, QN => n14294);
   REGISTERS_reg_4_42_inst : DFF_X1 port map( D => n7143, CK => CLK, Q => 
                           n18965, QN => n14295);
   REGISTERS_reg_4_41_inst : DFF_X1 port map( D => n7142, CK => CLK, Q => 
                           n18985, QN => n14296);
   REGISTERS_reg_4_40_inst : DFF_X1 port map( D => n7141, CK => CLK, Q => 
                           n19005, QN => n14297);
   REGISTERS_reg_4_39_inst : DFF_X1 port map( D => n7140, CK => CLK, Q => 
                           n19025, QN => n14298);
   REGISTERS_reg_4_38_inst : DFF_X1 port map( D => n7139, CK => CLK, Q => 
                           n19045, QN => n14299);
   REGISTERS_reg_4_37_inst : DFF_X1 port map( D => n7138, CK => CLK, Q => 
                           n19065, QN => n14300);
   REGISTERS_reg_4_36_inst : DFF_X1 port map( D => n7137, CK => CLK, Q => 
                           n19085, QN => n14301);
   REGISTERS_reg_4_35_inst : DFF_X1 port map( D => n7136, CK => CLK, Q => 
                           n19105, QN => n14302);
   REGISTERS_reg_4_34_inst : DFF_X1 port map( D => n7135, CK => CLK, Q => 
                           n19125, QN => n14303);
   REGISTERS_reg_4_33_inst : DFF_X1 port map( D => n7134, CK => CLK, Q => 
                           n19145, QN => n14304);
   REGISTERS_reg_4_32_inst : DFF_X1 port map( D => n7133, CK => CLK, Q => 
                           n19165, QN => n14305);
   REGISTERS_reg_4_31_inst : DFF_X1 port map( D => n7132, CK => CLK, Q => 
                           n19185, QN => n14306);
   REGISTERS_reg_4_30_inst : DFF_X1 port map( D => n7131, CK => CLK, Q => 
                           n19205, QN => n14307);
   REGISTERS_reg_4_29_inst : DFF_X1 port map( D => n7130, CK => CLK, Q => 
                           n19225, QN => n14308);
   REGISTERS_reg_4_28_inst : DFF_X1 port map( D => n7129, CK => CLK, Q => 
                           n19245, QN => n14309);
   REGISTERS_reg_4_27_inst : DFF_X1 port map( D => n7128, CK => CLK, Q => 
                           n19265, QN => n14310);
   REGISTERS_reg_4_26_inst : DFF_X1 port map( D => n7127, CK => CLK, Q => 
                           n19285, QN => n14311);
   REGISTERS_reg_4_25_inst : DFF_X1 port map( D => n7126, CK => CLK, Q => 
                           n19305, QN => n14312);
   REGISTERS_reg_4_24_inst : DFF_X1 port map( D => n7125, CK => CLK, Q => 
                           n19325, QN => n14313);
   REGISTERS_reg_4_23_inst : DFF_X1 port map( D => n7124, CK => CLK, Q => 
                           n19345, QN => n14314);
   REGISTERS_reg_4_22_inst : DFF_X1 port map( D => n7123, CK => CLK, Q => 
                           n19365, QN => n14315);
   REGISTERS_reg_4_21_inst : DFF_X1 port map( D => n7122, CK => CLK, Q => 
                           n19385, QN => n14316);
   REGISTERS_reg_4_20_inst : DFF_X1 port map( D => n7121, CK => CLK, Q => 
                           n19405, QN => n14317);
   REGISTERS_reg_4_19_inst : DFF_X1 port map( D => n7120, CK => CLK, Q => 
                           n19425, QN => n14318);
   REGISTERS_reg_4_18_inst : DFF_X1 port map( D => n7119, CK => CLK, Q => 
                           n19445, QN => n14319);
   REGISTERS_reg_4_17_inst : DFF_X1 port map( D => n7118, CK => CLK, Q => 
                           n19465, QN => n14320);
   REGISTERS_reg_4_16_inst : DFF_X1 port map( D => n7117, CK => CLK, Q => 
                           n19485, QN => n14321);
   REGISTERS_reg_4_15_inst : DFF_X1 port map( D => n7116, CK => CLK, Q => 
                           n19505, QN => n14322);
   REGISTERS_reg_4_14_inst : DFF_X1 port map( D => n7115, CK => CLK, Q => 
                           n19525, QN => n14323);
   REGISTERS_reg_4_13_inst : DFF_X1 port map( D => n7114, CK => CLK, Q => 
                           n19545, QN => n14324);
   REGISTERS_reg_4_12_inst : DFF_X1 port map( D => n7113, CK => CLK, Q => 
                           n19565, QN => n14325);
   REGISTERS_reg_4_11_inst : DFF_X1 port map( D => n7112, CK => CLK, Q => 
                           n19585, QN => n14326);
   REGISTERS_reg_4_10_inst : DFF_X1 port map( D => n7111, CK => CLK, Q => 
                           n19605, QN => n14327);
   REGISTERS_reg_4_9_inst : DFF_X1 port map( D => n7110, CK => CLK, Q => n19625
                           , QN => n14328);
   REGISTERS_reg_4_8_inst : DFF_X1 port map( D => n7109, CK => CLK, Q => n19645
                           , QN => n14329);
   REGISTERS_reg_4_7_inst : DFF_X1 port map( D => n7108, CK => CLK, Q => n19665
                           , QN => n14330);
   REGISTERS_reg_4_6_inst : DFF_X1 port map( D => n7107, CK => CLK, Q => n19685
                           , QN => n14331);
   REGISTERS_reg_4_5_inst : DFF_X1 port map( D => n7106, CK => CLK, Q => n19705
                           , QN => n14332);
   REGISTERS_reg_4_4_inst : DFF_X1 port map( D => n7105, CK => CLK, Q => n19725
                           , QN => n14333);
   REGISTERS_reg_4_3_inst : DFF_X1 port map( D => n7104, CK => CLK, Q => n19745
                           , QN => n14334);
   REGISTERS_reg_4_2_inst : DFF_X1 port map( D => n7103, CK => CLK, Q => n19765
                           , QN => n14335);
   REGISTERS_reg_4_1_inst : DFF_X1 port map( D => n7102, CK => CLK, Q => n19785
                           , QN => n14336);
   REGISTERS_reg_4_0_inst : DFF_X1 port map( D => n7101, CK => CLK, Q => n19805
                           , QN => n14337);
   REGISTERS_reg_5_59_inst : DFF_X1 port map( D => n7096, CK => CLK, Q => 
                           n20661, QN => n14345);
   REGISTERS_reg_5_58_inst : DFF_X1 port map( D => n7095, CK => CLK, Q => 
                           n20660, QN => n14346);
   REGISTERS_reg_5_57_inst : DFF_X1 port map( D => n7094, CK => CLK, Q => 
                           n20659, QN => n14347);
   REGISTERS_reg_5_56_inst : DFF_X1 port map( D => n7093, CK => CLK, Q => 
                           n20658, QN => n14348);
   REGISTERS_reg_5_55_inst : DFF_X1 port map( D => n7092, CK => CLK, Q => 
                           n20657, QN => n14349);
   REGISTERS_reg_5_54_inst : DFF_X1 port map( D => n7091, CK => CLK, Q => 
                           n20656, QN => n14350);
   REGISTERS_reg_5_53_inst : DFF_X1 port map( D => n7090, CK => CLK, Q => 
                           n20655, QN => n14351);
   REGISTERS_reg_5_52_inst : DFF_X1 port map( D => n7089, CK => CLK, Q => 
                           n20654, QN => n14352);
   REGISTERS_reg_5_51_inst : DFF_X1 port map( D => n7088, CK => CLK, Q => 
                           n20653, QN => n14353);
   REGISTERS_reg_5_50_inst : DFF_X1 port map( D => n7087, CK => CLK, Q => 
                           n20652, QN => n14354);
   REGISTERS_reg_5_49_inst : DFF_X1 port map( D => n7086, CK => CLK, Q => 
                           n20651, QN => n14355);
   REGISTERS_reg_5_48_inst : DFF_X1 port map( D => n7085, CK => CLK, Q => 
                           n20650, QN => n14356);
   REGISTERS_reg_5_47_inst : DFF_X1 port map( D => n7084, CK => CLK, Q => 
                           n20649, QN => n14357);
   REGISTERS_reg_5_46_inst : DFF_X1 port map( D => n7083, CK => CLK, Q => 
                           n20648, QN => n14358);
   REGISTERS_reg_5_45_inst : DFF_X1 port map( D => n7082, CK => CLK, Q => 
                           n20647, QN => n14359);
   REGISTERS_reg_5_44_inst : DFF_X1 port map( D => n7081, CK => CLK, Q => 
                           n20646, QN => n14360);
   REGISTERS_reg_5_43_inst : DFF_X1 port map( D => n7080, CK => CLK, Q => 
                           n20645, QN => n14361);
   REGISTERS_reg_5_42_inst : DFF_X1 port map( D => n7079, CK => CLK, Q => 
                           n20644, QN => n14362);
   REGISTERS_reg_5_41_inst : DFF_X1 port map( D => n7078, CK => CLK, Q => 
                           n20643, QN => n14363);
   REGISTERS_reg_5_40_inst : DFF_X1 port map( D => n7077, CK => CLK, Q => 
                           n20642, QN => n14364);
   REGISTERS_reg_5_39_inst : DFF_X1 port map( D => n7076, CK => CLK, Q => 
                           n20641, QN => n14365);
   REGISTERS_reg_5_38_inst : DFF_X1 port map( D => n7075, CK => CLK, Q => 
                           n20640, QN => n14366);
   REGISTERS_reg_5_37_inst : DFF_X1 port map( D => n7074, CK => CLK, Q => 
                           n20639, QN => n14367);
   REGISTERS_reg_5_36_inst : DFF_X1 port map( D => n7073, CK => CLK, Q => 
                           n20638, QN => n14368);
   REGISTERS_reg_5_35_inst : DFF_X1 port map( D => n7072, CK => CLK, Q => 
                           n20637, QN => n14369);
   REGISTERS_reg_5_34_inst : DFF_X1 port map( D => n7071, CK => CLK, Q => 
                           n20636, QN => n14370);
   REGISTERS_reg_5_33_inst : DFF_X1 port map( D => n7070, CK => CLK, Q => 
                           n20635, QN => n14371);
   REGISTERS_reg_5_32_inst : DFF_X1 port map( D => n7069, CK => CLK, Q => 
                           n20634, QN => n14372);
   REGISTERS_reg_5_31_inst : DFF_X1 port map( D => n7068, CK => CLK, Q => 
                           n20633, QN => n14373);
   REGISTERS_reg_5_30_inst : DFF_X1 port map( D => n7067, CK => CLK, Q => 
                           n20632, QN => n14374);
   REGISTERS_reg_5_29_inst : DFF_X1 port map( D => n7066, CK => CLK, Q => 
                           n20631, QN => n14375);
   REGISTERS_reg_5_28_inst : DFF_X1 port map( D => n7065, CK => CLK, Q => 
                           n20630, QN => n14376);
   REGISTERS_reg_5_27_inst : DFF_X1 port map( D => n7064, CK => CLK, Q => 
                           n20629, QN => n14377);
   REGISTERS_reg_5_26_inst : DFF_X1 port map( D => n7063, CK => CLK, Q => 
                           n20628, QN => n14378);
   REGISTERS_reg_5_25_inst : DFF_X1 port map( D => n7062, CK => CLK, Q => 
                           n20627, QN => n14379);
   REGISTERS_reg_5_24_inst : DFF_X1 port map( D => n7061, CK => CLK, Q => 
                           n20626, QN => n14380);
   REGISTERS_reg_5_23_inst : DFF_X1 port map( D => n7060, CK => CLK, Q => 
                           n20625, QN => n14381);
   REGISTERS_reg_5_22_inst : DFF_X1 port map( D => n7059, CK => CLK, Q => 
                           n20624, QN => n14382);
   REGISTERS_reg_5_21_inst : DFF_X1 port map( D => n7058, CK => CLK, Q => 
                           n20623, QN => n14383);
   REGISTERS_reg_5_20_inst : DFF_X1 port map( D => n7057, CK => CLK, Q => 
                           n20622, QN => n14384);
   REGISTERS_reg_5_19_inst : DFF_X1 port map( D => n7056, CK => CLK, Q => 
                           n20621, QN => n14385);
   REGISTERS_reg_5_18_inst : DFF_X1 port map( D => n7055, CK => CLK, Q => 
                           n20620, QN => n14386);
   REGISTERS_reg_5_17_inst : DFF_X1 port map( D => n7054, CK => CLK, Q => 
                           n20619, QN => n14387);
   REGISTERS_reg_5_16_inst : DFF_X1 port map( D => n7053, CK => CLK, Q => 
                           n20618, QN => n14388);
   REGISTERS_reg_5_15_inst : DFF_X1 port map( D => n7052, CK => CLK, Q => 
                           n20617, QN => n14389);
   REGISTERS_reg_5_14_inst : DFF_X1 port map( D => n7051, CK => CLK, Q => 
                           n20616, QN => n14390);
   REGISTERS_reg_5_13_inst : DFF_X1 port map( D => n7050, CK => CLK, Q => 
                           n20615, QN => n14391);
   REGISTERS_reg_5_12_inst : DFF_X1 port map( D => n7049, CK => CLK, Q => 
                           n20614, QN => n14392);
   REGISTERS_reg_5_11_inst : DFF_X1 port map( D => n7048, CK => CLK, Q => 
                           n20613, QN => n14393);
   REGISTERS_reg_5_10_inst : DFF_X1 port map( D => n7047, CK => CLK, Q => 
                           n20612, QN => n14394);
   REGISTERS_reg_5_9_inst : DFF_X1 port map( D => n7046, CK => CLK, Q => n20611
                           , QN => n14395);
   REGISTERS_reg_5_8_inst : DFF_X1 port map( D => n7045, CK => CLK, Q => n20610
                           , QN => n14396);
   REGISTERS_reg_5_7_inst : DFF_X1 port map( D => n7044, CK => CLK, Q => n20609
                           , QN => n14397);
   REGISTERS_reg_5_6_inst : DFF_X1 port map( D => n7043, CK => CLK, Q => n20608
                           , QN => n14398);
   REGISTERS_reg_5_5_inst : DFF_X1 port map( D => n7042, CK => CLK, Q => n20607
                           , QN => n14399);
   REGISTERS_reg_5_4_inst : DFF_X1 port map( D => n7041, CK => CLK, Q => n20606
                           , QN => n14400);
   REGISTERS_reg_5_3_inst : DFF_X1 port map( D => n7040, CK => CLK, Q => n20605
                           , QN => n14401);
   REGISTERS_reg_5_2_inst : DFF_X1 port map( D => n7039, CK => CLK, Q => n20604
                           , QN => n14402);
   REGISTERS_reg_5_1_inst : DFF_X1 port map( D => n7038, CK => CLK, Q => n20603
                           , QN => n14403);
   REGISTERS_reg_5_0_inst : DFF_X1 port map( D => n7037, CK => CLK, Q => n20602
                           , QN => n14404);
   REGISTERS_reg_7_59_inst : DFF_X1 port map( D => n6968, CK => CLK, Q => 
                           n20601, QN => n14481);
   REGISTERS_reg_7_58_inst : DFF_X1 port map( D => n6967, CK => CLK, Q => 
                           n20600, QN => n14482);
   REGISTERS_reg_7_57_inst : DFF_X1 port map( D => n6966, CK => CLK, Q => 
                           n20599, QN => n14483);
   REGISTERS_reg_7_56_inst : DFF_X1 port map( D => n6965, CK => CLK, Q => 
                           n20598, QN => n14484);
   REGISTERS_reg_7_55_inst : DFF_X1 port map( D => n6964, CK => CLK, Q => 
                           n20597, QN => n14485);
   REGISTERS_reg_7_54_inst : DFF_X1 port map( D => n6963, CK => CLK, Q => 
                           n20596, QN => n14486);
   REGISTERS_reg_7_53_inst : DFF_X1 port map( D => n6962, CK => CLK, Q => 
                           n20595, QN => n14487);
   REGISTERS_reg_7_52_inst : DFF_X1 port map( D => n6961, CK => CLK, Q => 
                           n20594, QN => n14488);
   REGISTERS_reg_7_51_inst : DFF_X1 port map( D => n6960, CK => CLK, Q => 
                           n20593, QN => n14489);
   REGISTERS_reg_7_50_inst : DFF_X1 port map( D => n6959, CK => CLK, Q => 
                           n20592, QN => n14490);
   REGISTERS_reg_7_49_inst : DFF_X1 port map( D => n6958, CK => CLK, Q => 
                           n20591, QN => n14491);
   REGISTERS_reg_7_48_inst : DFF_X1 port map( D => n6957, CK => CLK, Q => 
                           n20590, QN => n14492);
   REGISTERS_reg_7_47_inst : DFF_X1 port map( D => n6956, CK => CLK, Q => 
                           n20589, QN => n14493);
   REGISTERS_reg_7_46_inst : DFF_X1 port map( D => n6955, CK => CLK, Q => 
                           n20588, QN => n14494);
   REGISTERS_reg_7_45_inst : DFF_X1 port map( D => n6954, CK => CLK, Q => 
                           n20587, QN => n14495);
   REGISTERS_reg_7_44_inst : DFF_X1 port map( D => n6953, CK => CLK, Q => 
                           n20586, QN => n14496);
   REGISTERS_reg_7_43_inst : DFF_X1 port map( D => n6952, CK => CLK, Q => 
                           n20585, QN => n14497);
   REGISTERS_reg_7_42_inst : DFF_X1 port map( D => n6951, CK => CLK, Q => 
                           n20584, QN => n14498);
   REGISTERS_reg_7_41_inst : DFF_X1 port map( D => n6950, CK => CLK, Q => 
                           n20583, QN => n14499);
   REGISTERS_reg_7_40_inst : DFF_X1 port map( D => n6949, CK => CLK, Q => 
                           n20582, QN => n14500);
   REGISTERS_reg_7_39_inst : DFF_X1 port map( D => n6948, CK => CLK, Q => 
                           n20581, QN => n14501);
   REGISTERS_reg_7_38_inst : DFF_X1 port map( D => n6947, CK => CLK, Q => 
                           n20580, QN => n14502);
   REGISTERS_reg_7_37_inst : DFF_X1 port map( D => n6946, CK => CLK, Q => 
                           n20579, QN => n14503);
   REGISTERS_reg_7_36_inst : DFF_X1 port map( D => n6945, CK => CLK, Q => 
                           n20578, QN => n14504);
   REGISTERS_reg_7_35_inst : DFF_X1 port map( D => n6944, CK => CLK, Q => 
                           n20577, QN => n14505);
   REGISTERS_reg_7_34_inst : DFF_X1 port map( D => n6943, CK => CLK, Q => 
                           n20576, QN => n14506);
   REGISTERS_reg_7_33_inst : DFF_X1 port map( D => n6942, CK => CLK, Q => 
                           n20575, QN => n14507);
   REGISTERS_reg_7_32_inst : DFF_X1 port map( D => n6941, CK => CLK, Q => 
                           n20574, QN => n14508);
   REGISTERS_reg_7_31_inst : DFF_X1 port map( D => n6940, CK => CLK, Q => 
                           n20573, QN => n14509);
   REGISTERS_reg_7_30_inst : DFF_X1 port map( D => n6939, CK => CLK, Q => 
                           n20572, QN => n14510);
   REGISTERS_reg_7_29_inst : DFF_X1 port map( D => n6938, CK => CLK, Q => 
                           n20571, QN => n14511);
   REGISTERS_reg_7_28_inst : DFF_X1 port map( D => n6937, CK => CLK, Q => 
                           n20570, QN => n14512);
   REGISTERS_reg_7_27_inst : DFF_X1 port map( D => n6936, CK => CLK, Q => 
                           n20569, QN => n14513);
   REGISTERS_reg_7_26_inst : DFF_X1 port map( D => n6935, CK => CLK, Q => 
                           n20568, QN => n14514);
   REGISTERS_reg_7_25_inst : DFF_X1 port map( D => n6934, CK => CLK, Q => 
                           n20567, QN => n14515);
   REGISTERS_reg_7_24_inst : DFF_X1 port map( D => n6933, CK => CLK, Q => 
                           n20566, QN => n14516);
   REGISTERS_reg_7_23_inst : DFF_X1 port map( D => n6932, CK => CLK, Q => 
                           n20565, QN => n14517);
   REGISTERS_reg_7_22_inst : DFF_X1 port map( D => n6931, CK => CLK, Q => 
                           n20564, QN => n14518);
   REGISTERS_reg_7_21_inst : DFF_X1 port map( D => n6930, CK => CLK, Q => 
                           n20563, QN => n14519);
   REGISTERS_reg_7_20_inst : DFF_X1 port map( D => n6929, CK => CLK, Q => 
                           n20562, QN => n14520);
   REGISTERS_reg_7_19_inst : DFF_X1 port map( D => n6928, CK => CLK, Q => 
                           n20561, QN => n14521);
   REGISTERS_reg_7_18_inst : DFF_X1 port map( D => n6927, CK => CLK, Q => 
                           n20560, QN => n14522);
   REGISTERS_reg_7_17_inst : DFF_X1 port map( D => n6926, CK => CLK, Q => 
                           n20559, QN => n14523);
   REGISTERS_reg_7_16_inst : DFF_X1 port map( D => n6925, CK => CLK, Q => 
                           n20558, QN => n14524);
   REGISTERS_reg_7_15_inst : DFF_X1 port map( D => n6924, CK => CLK, Q => 
                           n20557, QN => n14525);
   REGISTERS_reg_7_14_inst : DFF_X1 port map( D => n6923, CK => CLK, Q => 
                           n20556, QN => n14526);
   REGISTERS_reg_7_13_inst : DFF_X1 port map( D => n6922, CK => CLK, Q => 
                           n20555, QN => n14527);
   REGISTERS_reg_7_12_inst : DFF_X1 port map( D => n6921, CK => CLK, Q => 
                           n20554, QN => n14528);
   REGISTERS_reg_7_11_inst : DFF_X1 port map( D => n6920, CK => CLK, Q => 
                           n20553, QN => n14529);
   REGISTERS_reg_7_10_inst : DFF_X1 port map( D => n6919, CK => CLK, Q => 
                           n20552, QN => n14530);
   REGISTERS_reg_7_9_inst : DFF_X1 port map( D => n6918, CK => CLK, Q => n20551
                           , QN => n14531);
   REGISTERS_reg_7_8_inst : DFF_X1 port map( D => n6917, CK => CLK, Q => n20550
                           , QN => n14532);
   REGISTERS_reg_7_7_inst : DFF_X1 port map( D => n6916, CK => CLK, Q => n20549
                           , QN => n14533);
   REGISTERS_reg_7_6_inst : DFF_X1 port map( D => n6915, CK => CLK, Q => n20548
                           , QN => n14534);
   REGISTERS_reg_7_5_inst : DFF_X1 port map( D => n6914, CK => CLK, Q => n20547
                           , QN => n14535);
   REGISTERS_reg_7_4_inst : DFF_X1 port map( D => n6913, CK => CLK, Q => n20546
                           , QN => n14536);
   REGISTERS_reg_7_3_inst : DFF_X1 port map( D => n6912, CK => CLK, Q => n20545
                           , QN => n14537);
   REGISTERS_reg_7_2_inst : DFF_X1 port map( D => n6911, CK => CLK, Q => n20544
                           , QN => n14538);
   REGISTERS_reg_7_1_inst : DFF_X1 port map( D => n6910, CK => CLK, Q => n20543
                           , QN => n14539);
   REGISTERS_reg_7_0_inst : DFF_X1 port map( D => n6909, CK => CLK, Q => n20542
                           , QN => n14540);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n7224, CK => CLK, Q => 
                           n20541, QN => n14212);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n7223, CK => CLK, Q => 
                           n20540, QN => n14213);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n7222, CK => CLK, Q => 
                           n20539, QN => n14214);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n7221, CK => CLK, Q => 
                           n20538, QN => n14215);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n7220, CK => CLK, Q => 
                           n20537, QN => n14216);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n7219, CK => CLK, Q => 
                           n20536, QN => n14217);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n7218, CK => CLK, Q => 
                           n20535, QN => n14218);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n7217, CK => CLK, Q => 
                           n20534, QN => n14219);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n7216, CK => CLK, Q => 
                           n20533, QN => n14220);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n7215, CK => CLK, Q => 
                           n20532, QN => n14221);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n7214, CK => CLK, Q => 
                           n20531, QN => n14222);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n7213, CK => CLK, Q => 
                           n20530, QN => n14223);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n7212, CK => CLK, Q => 
                           n20529, QN => n14224);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n7211, CK => CLK, Q => 
                           n20528, QN => n14225);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n7210, CK => CLK, Q => 
                           n20527, QN => n14226);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n7209, CK => CLK, Q => 
                           n20526, QN => n14227);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n7208, CK => CLK, Q => 
                           n20525, QN => n14228);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n7207, CK => CLK, Q => 
                           n20524, QN => n14229);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n7206, CK => CLK, Q => 
                           n20523, QN => n14230);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n7205, CK => CLK, Q => 
                           n20522, QN => n14231);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n7204, CK => CLK, Q => 
                           n20521, QN => n14232);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n7203, CK => CLK, Q => 
                           n20520, QN => n14233);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n7202, CK => CLK, Q => 
                           n20519, QN => n14234);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n7201, CK => CLK, Q => 
                           n20518, QN => n14235);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n7200, CK => CLK, Q => 
                           n20517, QN => n14236);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n7199, CK => CLK, Q => 
                           n20516, QN => n14237);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n7198, CK => CLK, Q => 
                           n20515, QN => n14238);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n7197, CK => CLK, Q => 
                           n20514, QN => n14239);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n7196, CK => CLK, Q => 
                           n20513, QN => n14240);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n7195, CK => CLK, Q => 
                           n20512, QN => n14241);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n7194, CK => CLK, Q => 
                           n20511, QN => n14242);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n7193, CK => CLK, Q => 
                           n20510, QN => n14243);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n7192, CK => CLK, Q => 
                           n20509, QN => n14244);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n7191, CK => CLK, Q => 
                           n20508, QN => n14245);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n7190, CK => CLK, Q => 
                           n20507, QN => n14246);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n7189, CK => CLK, Q => 
                           n20506, QN => n14247);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n7188, CK => CLK, Q => 
                           n20505, QN => n14248);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n7187, CK => CLK, Q => 
                           n20504, QN => n14249);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n7186, CK => CLK, Q => 
                           n20503, QN => n14250);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n7185, CK => CLK, Q => 
                           n20502, QN => n14251);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n7184, CK => CLK, Q => 
                           n20501, QN => n14252);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n7183, CK => CLK, Q => 
                           n20500, QN => n14253);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n7182, CK => CLK, Q => 
                           n20499, QN => n14254);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n7181, CK => CLK, Q => 
                           n20498, QN => n14255);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n7180, CK => CLK, Q => 
                           n20497, QN => n14256);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n7179, CK => CLK, Q => 
                           n20496, QN => n14257);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n7178, CK => CLK, Q => 
                           n20495, QN => n14258);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n7177, CK => CLK, Q => 
                           n20494, QN => n14259);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n7176, CK => CLK, Q => 
                           n20493, QN => n14260);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n7175, CK => CLK, Q => 
                           n20492, QN => n14261);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n7174, CK => CLK, Q => n20491
                           , QN => n14262);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n7173, CK => CLK, Q => n20490
                           , QN => n14263);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n7172, CK => CLK, Q => n20489
                           , QN => n14264);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n7171, CK => CLK, Q => n20488
                           , QN => n14265);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n7170, CK => CLK, Q => n20487
                           , QN => n14266);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n7169, CK => CLK, Q => n20486
                           , QN => n14267);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n7168, CK => CLK, Q => n20485
                           , QN => n14268);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n7167, CK => CLK, Q => n20484
                           , QN => n14269);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n7166, CK => CLK, Q => n20483
                           , QN => n14270);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n7165, CK => CLK, Q => n20482
                           , QN => n14271);
   REGISTERS_reg_10_59_inst : DFF_X1 port map( D => n6776, CK => CLK, Q => 
                           n18639, QN => n14681);
   REGISTERS_reg_10_58_inst : DFF_X1 port map( D => n6775, CK => CLK, Q => 
                           n18659, QN => n14682);
   REGISTERS_reg_10_57_inst : DFF_X1 port map( D => n6774, CK => CLK, Q => 
                           n18679, QN => n14683);
   REGISTERS_reg_10_56_inst : DFF_X1 port map( D => n6773, CK => CLK, Q => 
                           n18699, QN => n14684);
   REGISTERS_reg_10_55_inst : DFF_X1 port map( D => n6772, CK => CLK, Q => 
                           n18719, QN => n14685);
   REGISTERS_reg_10_54_inst : DFF_X1 port map( D => n6771, CK => CLK, Q => 
                           n18739, QN => n14686);
   REGISTERS_reg_10_53_inst : DFF_X1 port map( D => n6770, CK => CLK, Q => 
                           n18759, QN => n14687);
   REGISTERS_reg_10_52_inst : DFF_X1 port map( D => n6769, CK => CLK, Q => 
                           n18779, QN => n14688);
   REGISTERS_reg_10_51_inst : DFF_X1 port map( D => n6768, CK => CLK, Q => 
                           n18799, QN => n14689);
   REGISTERS_reg_10_50_inst : DFF_X1 port map( D => n6767, CK => CLK, Q => 
                           n18819, QN => n14690);
   REGISTERS_reg_10_49_inst : DFF_X1 port map( D => n6766, CK => CLK, Q => 
                           n18839, QN => n14691);
   REGISTERS_reg_10_48_inst : DFF_X1 port map( D => n6765, CK => CLK, Q => 
                           n18859, QN => n14692);
   REGISTERS_reg_10_47_inst : DFF_X1 port map( D => n6764, CK => CLK, Q => 
                           n18879, QN => n14693);
   REGISTERS_reg_10_46_inst : DFF_X1 port map( D => n6763, CK => CLK, Q => 
                           n18899, QN => n14694);
   REGISTERS_reg_10_45_inst : DFF_X1 port map( D => n6762, CK => CLK, Q => 
                           n18919, QN => n14695);
   REGISTERS_reg_10_44_inst : DFF_X1 port map( D => n6761, CK => CLK, Q => 
                           n18939, QN => n14696);
   REGISTERS_reg_10_43_inst : DFF_X1 port map( D => n6760, CK => CLK, Q => 
                           n18959, QN => n14697);
   REGISTERS_reg_10_42_inst : DFF_X1 port map( D => n6759, CK => CLK, Q => 
                           n18979, QN => n14698);
   REGISTERS_reg_10_41_inst : DFF_X1 port map( D => n6758, CK => CLK, Q => 
                           n18999, QN => n14699);
   REGISTERS_reg_10_40_inst : DFF_X1 port map( D => n6757, CK => CLK, Q => 
                           n19019, QN => n14700);
   REGISTERS_reg_10_39_inst : DFF_X1 port map( D => n6756, CK => CLK, Q => 
                           n19039, QN => n14701);
   REGISTERS_reg_10_38_inst : DFF_X1 port map( D => n6755, CK => CLK, Q => 
                           n19059, QN => n14702);
   REGISTERS_reg_10_37_inst : DFF_X1 port map( D => n6754, CK => CLK, Q => 
                           n19079, QN => n14703);
   REGISTERS_reg_10_36_inst : DFF_X1 port map( D => n6753, CK => CLK, Q => 
                           n19099, QN => n14704);
   REGISTERS_reg_10_35_inst : DFF_X1 port map( D => n6752, CK => CLK, Q => 
                           n19119, QN => n14705);
   REGISTERS_reg_10_34_inst : DFF_X1 port map( D => n6751, CK => CLK, Q => 
                           n19139, QN => n14706);
   REGISTERS_reg_10_33_inst : DFF_X1 port map( D => n6750, CK => CLK, Q => 
                           n19159, QN => n14707);
   REGISTERS_reg_10_32_inst : DFF_X1 port map( D => n6749, CK => CLK, Q => 
                           n19179, QN => n14708);
   REGISTERS_reg_10_31_inst : DFF_X1 port map( D => n6748, CK => CLK, Q => 
                           n19199, QN => n14709);
   REGISTERS_reg_10_30_inst : DFF_X1 port map( D => n6747, CK => CLK, Q => 
                           n19219, QN => n14710);
   REGISTERS_reg_10_29_inst : DFF_X1 port map( D => n6746, CK => CLK, Q => 
                           n19239, QN => n14711);
   REGISTERS_reg_10_28_inst : DFF_X1 port map( D => n6745, CK => CLK, Q => 
                           n19259, QN => n14712);
   REGISTERS_reg_10_27_inst : DFF_X1 port map( D => n6744, CK => CLK, Q => 
                           n19279, QN => n14713);
   REGISTERS_reg_10_26_inst : DFF_X1 port map( D => n6743, CK => CLK, Q => 
                           n19299, QN => n14714);
   REGISTERS_reg_10_25_inst : DFF_X1 port map( D => n6742, CK => CLK, Q => 
                           n19319, QN => n14715);
   REGISTERS_reg_10_24_inst : DFF_X1 port map( D => n6741, CK => CLK, Q => 
                           n19339, QN => n14716);
   REGISTERS_reg_10_23_inst : DFF_X1 port map( D => n6740, CK => CLK, Q => 
                           n19359, QN => n14717);
   REGISTERS_reg_10_22_inst : DFF_X1 port map( D => n6739, CK => CLK, Q => 
                           n19379, QN => n14718);
   REGISTERS_reg_10_21_inst : DFF_X1 port map( D => n6738, CK => CLK, Q => 
                           n19399, QN => n14719);
   REGISTERS_reg_10_20_inst : DFF_X1 port map( D => n6737, CK => CLK, Q => 
                           n19419, QN => n14720);
   REGISTERS_reg_10_19_inst : DFF_X1 port map( D => n6736, CK => CLK, Q => 
                           n19439, QN => n14721);
   REGISTERS_reg_10_18_inst : DFF_X1 port map( D => n6735, CK => CLK, Q => 
                           n19459, QN => n14722);
   REGISTERS_reg_10_17_inst : DFF_X1 port map( D => n6734, CK => CLK, Q => 
                           n19479, QN => n14723);
   REGISTERS_reg_10_16_inst : DFF_X1 port map( D => n6733, CK => CLK, Q => 
                           n19499, QN => n14724);
   REGISTERS_reg_10_15_inst : DFF_X1 port map( D => n6732, CK => CLK, Q => 
                           n19519, QN => n14725);
   REGISTERS_reg_10_14_inst : DFF_X1 port map( D => n6731, CK => CLK, Q => 
                           n19539, QN => n14726);
   REGISTERS_reg_10_13_inst : DFF_X1 port map( D => n6730, CK => CLK, Q => 
                           n19559, QN => n14727);
   REGISTERS_reg_10_12_inst : DFF_X1 port map( D => n6729, CK => CLK, Q => 
                           n19579, QN => n14728);
   REGISTERS_reg_10_11_inst : DFF_X1 port map( D => n6728, CK => CLK, Q => 
                           n19599, QN => n14729);
   REGISTERS_reg_10_10_inst : DFF_X1 port map( D => n6727, CK => CLK, Q => 
                           n19619, QN => n14730);
   REGISTERS_reg_10_9_inst : DFF_X1 port map( D => n6726, CK => CLK, Q => 
                           n19639, QN => n14731);
   REGISTERS_reg_10_8_inst : DFF_X1 port map( D => n6725, CK => CLK, Q => 
                           n19659, QN => n14732);
   REGISTERS_reg_10_7_inst : DFF_X1 port map( D => n6724, CK => CLK, Q => 
                           n19679, QN => n14733);
   REGISTERS_reg_10_6_inst : DFF_X1 port map( D => n6723, CK => CLK, Q => 
                           n19699, QN => n14734);
   REGISTERS_reg_10_5_inst : DFF_X1 port map( D => n6722, CK => CLK, Q => 
                           n19719, QN => n14735);
   REGISTERS_reg_10_4_inst : DFF_X1 port map( D => n6721, CK => CLK, Q => 
                           n19739, QN => n14736);
   REGISTERS_reg_10_3_inst : DFF_X1 port map( D => n6720, CK => CLK, Q => 
                           n19759, QN => n14737);
   REGISTERS_reg_10_2_inst : DFF_X1 port map( D => n6719, CK => CLK, Q => 
                           n19779, QN => n14738);
   REGISTERS_reg_10_1_inst : DFF_X1 port map( D => n6718, CK => CLK, Q => 
                           n19799, QN => n14739);
   REGISTERS_reg_10_0_inst : DFF_X1 port map( D => n6717, CK => CLK, Q => 
                           n19819, QN => n14740);
   REGISTERS_reg_8_59_inst : DFF_X1 port map( D => n6904, CK => CLK, Q => n8976
                           , QN => n14547);
   REGISTERS_reg_8_58_inst : DFF_X1 port map( D => n6903, CK => CLK, Q => n8980
                           , QN => n14548);
   REGISTERS_reg_8_57_inst : DFF_X1 port map( D => n6902, CK => CLK, Q => n8984
                           , QN => n14549);
   REGISTERS_reg_8_56_inst : DFF_X1 port map( D => n6901, CK => CLK, Q => n8988
                           , QN => n14550);
   REGISTERS_reg_8_55_inst : DFF_X1 port map( D => n6900, CK => CLK, Q => n8992
                           , QN => n14551);
   REGISTERS_reg_8_54_inst : DFF_X1 port map( D => n6899, CK => CLK, Q => n8996
                           , QN => n14552);
   REGISTERS_reg_8_53_inst : DFF_X1 port map( D => n6898, CK => CLK, Q => n9000
                           , QN => n14553);
   REGISTERS_reg_8_52_inst : DFF_X1 port map( D => n6897, CK => CLK, Q => n9004
                           , QN => n14554);
   REGISTERS_reg_8_51_inst : DFF_X1 port map( D => n6896, CK => CLK, Q => n9008
                           , QN => n14555);
   REGISTERS_reg_8_50_inst : DFF_X1 port map( D => n6895, CK => CLK, Q => n9012
                           , QN => n14556);
   REGISTERS_reg_8_49_inst : DFF_X1 port map( D => n6894, CK => CLK, Q => n9016
                           , QN => n14557);
   REGISTERS_reg_8_48_inst : DFF_X1 port map( D => n6893, CK => CLK, Q => n9020
                           , QN => n14558);
   REGISTERS_reg_8_47_inst : DFF_X1 port map( D => n6892, CK => CLK, Q => n9024
                           , QN => n14559);
   REGISTERS_reg_8_46_inst : DFF_X1 port map( D => n6891, CK => CLK, Q => n9028
                           , QN => n14560);
   REGISTERS_reg_8_45_inst : DFF_X1 port map( D => n6890, CK => CLK, Q => n9032
                           , QN => n14561);
   REGISTERS_reg_8_44_inst : DFF_X1 port map( D => n6889, CK => CLK, Q => n9036
                           , QN => n14562);
   REGISTERS_reg_8_43_inst : DFF_X1 port map( D => n6888, CK => CLK, Q => n9040
                           , QN => n14563);
   REGISTERS_reg_8_42_inst : DFF_X1 port map( D => n6887, CK => CLK, Q => n9044
                           , QN => n14564);
   REGISTERS_reg_8_41_inst : DFF_X1 port map( D => n6886, CK => CLK, Q => n9048
                           , QN => n14565);
   REGISTERS_reg_8_40_inst : DFF_X1 port map( D => n6885, CK => CLK, Q => n9052
                           , QN => n14566);
   REGISTERS_reg_8_39_inst : DFF_X1 port map( D => n6884, CK => CLK, Q => n9056
                           , QN => n14567);
   REGISTERS_reg_8_38_inst : DFF_X1 port map( D => n6883, CK => CLK, Q => n9060
                           , QN => n14568);
   REGISTERS_reg_8_37_inst : DFF_X1 port map( D => n6882, CK => CLK, Q => n9064
                           , QN => n14569);
   REGISTERS_reg_8_36_inst : DFF_X1 port map( D => n6881, CK => CLK, Q => n9068
                           , QN => n14570);
   REGISTERS_reg_8_35_inst : DFF_X1 port map( D => n6880, CK => CLK, Q => n9072
                           , QN => n14571);
   REGISTERS_reg_8_34_inst : DFF_X1 port map( D => n6879, CK => CLK, Q => n9076
                           , QN => n14572);
   REGISTERS_reg_8_33_inst : DFF_X1 port map( D => n6878, CK => CLK, Q => n9080
                           , QN => n14573);
   REGISTERS_reg_8_32_inst : DFF_X1 port map( D => n6877, CK => CLK, Q => n9084
                           , QN => n14574);
   REGISTERS_reg_8_31_inst : DFF_X1 port map( D => n6876, CK => CLK, Q => n9088
                           , QN => n14575);
   REGISTERS_reg_8_30_inst : DFF_X1 port map( D => n6875, CK => CLK, Q => n9092
                           , QN => n14576);
   REGISTERS_reg_8_29_inst : DFF_X1 port map( D => n6874, CK => CLK, Q => n9096
                           , QN => n14577);
   REGISTERS_reg_8_28_inst : DFF_X1 port map( D => n6873, CK => CLK, Q => n9100
                           , QN => n14578);
   REGISTERS_reg_8_27_inst : DFF_X1 port map( D => n6872, CK => CLK, Q => n9104
                           , QN => n14579);
   REGISTERS_reg_8_26_inst : DFF_X1 port map( D => n6871, CK => CLK, Q => n9108
                           , QN => n14580);
   REGISTERS_reg_8_25_inst : DFF_X1 port map( D => n6870, CK => CLK, Q => n9112
                           , QN => n14581);
   REGISTERS_reg_8_24_inst : DFF_X1 port map( D => n6869, CK => CLK, Q => n9116
                           , QN => n14582);
   REGISTERS_reg_8_23_inst : DFF_X1 port map( D => n6868, CK => CLK, Q => n9120
                           , QN => n14583);
   REGISTERS_reg_8_22_inst : DFF_X1 port map( D => n6867, CK => CLK, Q => n9124
                           , QN => n14584);
   REGISTERS_reg_8_21_inst : DFF_X1 port map( D => n6866, CK => CLK, Q => n9128
                           , QN => n14585);
   REGISTERS_reg_8_20_inst : DFF_X1 port map( D => n6865, CK => CLK, Q => n9132
                           , QN => n14586);
   REGISTERS_reg_8_19_inst : DFF_X1 port map( D => n6864, CK => CLK, Q => n9136
                           , QN => n14587);
   REGISTERS_reg_8_18_inst : DFF_X1 port map( D => n6863, CK => CLK, Q => n9140
                           , QN => n14588);
   REGISTERS_reg_8_17_inst : DFF_X1 port map( D => n6862, CK => CLK, Q => n9144
                           , QN => n14589);
   REGISTERS_reg_8_16_inst : DFF_X1 port map( D => n6861, CK => CLK, Q => n9148
                           , QN => n14590);
   REGISTERS_reg_8_15_inst : DFF_X1 port map( D => n6860, CK => CLK, Q => n9152
                           , QN => n14591);
   REGISTERS_reg_8_14_inst : DFF_X1 port map( D => n6859, CK => CLK, Q => n9156
                           , QN => n14592);
   REGISTERS_reg_8_13_inst : DFF_X1 port map( D => n6858, CK => CLK, Q => n9160
                           , QN => n14593);
   REGISTERS_reg_8_12_inst : DFF_X1 port map( D => n6857, CK => CLK, Q => n9164
                           , QN => n14594);
   REGISTERS_reg_8_11_inst : DFF_X1 port map( D => n6856, CK => CLK, Q => n9168
                           , QN => n14595);
   REGISTERS_reg_8_10_inst : DFF_X1 port map( D => n6855, CK => CLK, Q => n9172
                           , QN => n14596);
   REGISTERS_reg_8_9_inst : DFF_X1 port map( D => n6854, CK => CLK, Q => n9176,
                           QN => n14597);
   REGISTERS_reg_8_8_inst : DFF_X1 port map( D => n6853, CK => CLK, Q => n9180,
                           QN => n14598);
   REGISTERS_reg_8_7_inst : DFF_X1 port map( D => n6852, CK => CLK, Q => n9184,
                           QN => n14599);
   REGISTERS_reg_8_6_inst : DFF_X1 port map( D => n6851, CK => CLK, Q => n9188,
                           QN => n14600);
   REGISTERS_reg_8_5_inst : DFF_X1 port map( D => n6850, CK => CLK, Q => n9192,
                           QN => n14601);
   REGISTERS_reg_8_4_inst : DFF_X1 port map( D => n6849, CK => CLK, Q => n9196,
                           QN => n14602);
   REGISTERS_reg_8_3_inst : DFF_X1 port map( D => n6848, CK => CLK, Q => n9200,
                           QN => n14603);
   REGISTERS_reg_8_2_inst : DFF_X1 port map( D => n6847, CK => CLK, Q => n9204,
                           QN => n14604);
   REGISTERS_reg_8_1_inst : DFF_X1 port map( D => n6846, CK => CLK, Q => n9208,
                           QN => n14605);
   REGISTERS_reg_8_0_inst : DFF_X1 port map( D => n6845, CK => CLK, Q => n9212,
                           QN => n14606);
   REGISTERS_reg_14_59_inst : DFF_X1 port map( D => n6520, CK => CLK, Q => 
                           n20481, QN => n14945);
   REGISTERS_reg_14_58_inst : DFF_X1 port map( D => n6519, CK => CLK, Q => 
                           n20480, QN => n14946);
   REGISTERS_reg_14_57_inst : DFF_X1 port map( D => n6518, CK => CLK, Q => 
                           n20479, QN => n14947);
   REGISTERS_reg_14_56_inst : DFF_X1 port map( D => n6517, CK => CLK, Q => 
                           n20478, QN => n14948);
   REGISTERS_reg_14_55_inst : DFF_X1 port map( D => n6516, CK => CLK, Q => 
                           n20477, QN => n14949);
   REGISTERS_reg_14_54_inst : DFF_X1 port map( D => n6515, CK => CLK, Q => 
                           n20476, QN => n14950);
   REGISTERS_reg_14_53_inst : DFF_X1 port map( D => n6514, CK => CLK, Q => 
                           n20475, QN => n14951);
   REGISTERS_reg_14_52_inst : DFF_X1 port map( D => n6513, CK => CLK, Q => 
                           n20474, QN => n14952);
   REGISTERS_reg_14_51_inst : DFF_X1 port map( D => n6512, CK => CLK, Q => 
                           n20473, QN => n14953);
   REGISTERS_reg_14_50_inst : DFF_X1 port map( D => n6511, CK => CLK, Q => 
                           n20472, QN => n14954);
   REGISTERS_reg_14_49_inst : DFF_X1 port map( D => n6510, CK => CLK, Q => 
                           n20471, QN => n14955);
   REGISTERS_reg_14_48_inst : DFF_X1 port map( D => n6509, CK => CLK, Q => 
                           n20470, QN => n14956);
   REGISTERS_reg_14_47_inst : DFF_X1 port map( D => n6508, CK => CLK, Q => 
                           n20469, QN => n14957);
   REGISTERS_reg_14_46_inst : DFF_X1 port map( D => n6507, CK => CLK, Q => 
                           n20468, QN => n14958);
   REGISTERS_reg_14_45_inst : DFF_X1 port map( D => n6506, CK => CLK, Q => 
                           n20467, QN => n14959);
   REGISTERS_reg_14_44_inst : DFF_X1 port map( D => n6505, CK => CLK, Q => 
                           n20466, QN => n14960);
   REGISTERS_reg_14_43_inst : DFF_X1 port map( D => n6504, CK => CLK, Q => 
                           n20465, QN => n14961);
   REGISTERS_reg_14_42_inst : DFF_X1 port map( D => n6503, CK => CLK, Q => 
                           n20464, QN => n14962);
   REGISTERS_reg_14_41_inst : DFF_X1 port map( D => n6502, CK => CLK, Q => 
                           n20463, QN => n14963);
   REGISTERS_reg_14_40_inst : DFF_X1 port map( D => n6501, CK => CLK, Q => 
                           n20462, QN => n14964);
   REGISTERS_reg_14_39_inst : DFF_X1 port map( D => n6500, CK => CLK, Q => 
                           n20461, QN => n14965);
   REGISTERS_reg_14_38_inst : DFF_X1 port map( D => n6499, CK => CLK, Q => 
                           n20460, QN => n14966);
   REGISTERS_reg_14_37_inst : DFF_X1 port map( D => n6498, CK => CLK, Q => 
                           n20459, QN => n14967);
   REGISTERS_reg_14_36_inst : DFF_X1 port map( D => n6497, CK => CLK, Q => 
                           n20458, QN => n14968);
   REGISTERS_reg_14_35_inst : DFF_X1 port map( D => n6496, CK => CLK, Q => 
                           n20457, QN => n14969);
   REGISTERS_reg_14_34_inst : DFF_X1 port map( D => n6495, CK => CLK, Q => 
                           n20456, QN => n14970);
   REGISTERS_reg_14_33_inst : DFF_X1 port map( D => n6494, CK => CLK, Q => 
                           n20455, QN => n14971);
   REGISTERS_reg_14_32_inst : DFF_X1 port map( D => n6493, CK => CLK, Q => 
                           n20454, QN => n14972);
   REGISTERS_reg_14_31_inst : DFF_X1 port map( D => n6492, CK => CLK, Q => 
                           n20453, QN => n14973);
   REGISTERS_reg_14_30_inst : DFF_X1 port map( D => n6491, CK => CLK, Q => 
                           n20452, QN => n14974);
   REGISTERS_reg_14_29_inst : DFF_X1 port map( D => n6490, CK => CLK, Q => 
                           n20451, QN => n14975);
   REGISTERS_reg_14_28_inst : DFF_X1 port map( D => n6489, CK => CLK, Q => 
                           n20450, QN => n14976);
   REGISTERS_reg_14_27_inst : DFF_X1 port map( D => n6488, CK => CLK, Q => 
                           n20449, QN => n14977);
   REGISTERS_reg_14_26_inst : DFF_X1 port map( D => n6487, CK => CLK, Q => 
                           n20448, QN => n14978);
   REGISTERS_reg_14_25_inst : DFF_X1 port map( D => n6486, CK => CLK, Q => 
                           n20447, QN => n14979);
   REGISTERS_reg_14_24_inst : DFF_X1 port map( D => n6485, CK => CLK, Q => 
                           n20446, QN => n14980);
   REGISTERS_reg_14_23_inst : DFF_X1 port map( D => n6484, CK => CLK, Q => 
                           n20445, QN => n14981);
   REGISTERS_reg_14_22_inst : DFF_X1 port map( D => n6483, CK => CLK, Q => 
                           n20444, QN => n14982);
   REGISTERS_reg_14_21_inst : DFF_X1 port map( D => n6482, CK => CLK, Q => 
                           n20443, QN => n14983);
   REGISTERS_reg_14_20_inst : DFF_X1 port map( D => n6481, CK => CLK, Q => 
                           n20442, QN => n14984);
   REGISTERS_reg_14_19_inst : DFF_X1 port map( D => n6480, CK => CLK, Q => 
                           n20441, QN => n14985);
   REGISTERS_reg_14_18_inst : DFF_X1 port map( D => n6479, CK => CLK, Q => 
                           n20440, QN => n14986);
   REGISTERS_reg_14_17_inst : DFF_X1 port map( D => n6478, CK => CLK, Q => 
                           n20439, QN => n14987);
   REGISTERS_reg_14_16_inst : DFF_X1 port map( D => n6477, CK => CLK, Q => 
                           n20438, QN => n14988);
   REGISTERS_reg_14_15_inst : DFF_X1 port map( D => n6476, CK => CLK, Q => 
                           n20437, QN => n14989);
   REGISTERS_reg_14_14_inst : DFF_X1 port map( D => n6475, CK => CLK, Q => 
                           n20436, QN => n14990);
   REGISTERS_reg_14_13_inst : DFF_X1 port map( D => n6474, CK => CLK, Q => 
                           n20435, QN => n14991);
   REGISTERS_reg_14_12_inst : DFF_X1 port map( D => n6473, CK => CLK, Q => 
                           n20434, QN => n14992);
   REGISTERS_reg_14_11_inst : DFF_X1 port map( D => n6472, CK => CLK, Q => 
                           n20433, QN => n14993);
   REGISTERS_reg_14_10_inst : DFF_X1 port map( D => n6471, CK => CLK, Q => 
                           n20432, QN => n14994);
   REGISTERS_reg_14_9_inst : DFF_X1 port map( D => n6470, CK => CLK, Q => 
                           n20431, QN => n14995);
   REGISTERS_reg_14_8_inst : DFF_X1 port map( D => n6469, CK => CLK, Q => 
                           n20430, QN => n14996);
   REGISTERS_reg_14_7_inst : DFF_X1 port map( D => n6468, CK => CLK, Q => 
                           n20429, QN => n14997);
   REGISTERS_reg_14_6_inst : DFF_X1 port map( D => n6467, CK => CLK, Q => 
                           n20428, QN => n14998);
   REGISTERS_reg_14_5_inst : DFF_X1 port map( D => n6466, CK => CLK, Q => 
                           n20427, QN => n14999);
   REGISTERS_reg_14_4_inst : DFF_X1 port map( D => n6465, CK => CLK, Q => 
                           n20426, QN => n15000);
   REGISTERS_reg_14_3_inst : DFF_X1 port map( D => n6464, CK => CLK, Q => 
                           n20425, QN => n15001);
   REGISTERS_reg_14_2_inst : DFF_X1 port map( D => n6463, CK => CLK, Q => 
                           n20424, QN => n15002);
   REGISTERS_reg_14_1_inst : DFF_X1 port map( D => n6462, CK => CLK, Q => 
                           n20423, QN => n15003);
   REGISTERS_reg_14_0_inst : DFF_X1 port map( D => n6461, CK => CLK, Q => 
                           n20422, QN => n15004);
   REGISTERS_reg_12_59_inst : DFF_X1 port map( D => n6648, CK => CLK, Q => 
                           n20421, QN => n14813);
   REGISTERS_reg_12_58_inst : DFF_X1 port map( D => n6647, CK => CLK, Q => 
                           n20420, QN => n14814);
   REGISTERS_reg_12_57_inst : DFF_X1 port map( D => n6646, CK => CLK, Q => 
                           n20419, QN => n14815);
   REGISTERS_reg_12_56_inst : DFF_X1 port map( D => n6645, CK => CLK, Q => 
                           n20418, QN => n14816);
   REGISTERS_reg_12_55_inst : DFF_X1 port map( D => n6644, CK => CLK, Q => 
                           n20417, QN => n14817);
   REGISTERS_reg_12_54_inst : DFF_X1 port map( D => n6643, CK => CLK, Q => 
                           n20416, QN => n14818);
   REGISTERS_reg_12_53_inst : DFF_X1 port map( D => n6642, CK => CLK, Q => 
                           n20415, QN => n14819);
   REGISTERS_reg_12_52_inst : DFF_X1 port map( D => n6641, CK => CLK, Q => 
                           n20414, QN => n14820);
   REGISTERS_reg_12_51_inst : DFF_X1 port map( D => n6640, CK => CLK, Q => 
                           n20413, QN => n14821);
   REGISTERS_reg_12_50_inst : DFF_X1 port map( D => n6639, CK => CLK, Q => 
                           n20412, QN => n14822);
   REGISTERS_reg_12_49_inst : DFF_X1 port map( D => n6638, CK => CLK, Q => 
                           n20411, QN => n14823);
   REGISTERS_reg_12_48_inst : DFF_X1 port map( D => n6637, CK => CLK, Q => 
                           n20410, QN => n14824);
   REGISTERS_reg_12_47_inst : DFF_X1 port map( D => n6636, CK => CLK, Q => 
                           n20409, QN => n14825);
   REGISTERS_reg_12_46_inst : DFF_X1 port map( D => n6635, CK => CLK, Q => 
                           n20408, QN => n14826);
   REGISTERS_reg_12_45_inst : DFF_X1 port map( D => n6634, CK => CLK, Q => 
                           n20407, QN => n14827);
   REGISTERS_reg_12_44_inst : DFF_X1 port map( D => n6633, CK => CLK, Q => 
                           n20406, QN => n14828);
   REGISTERS_reg_12_43_inst : DFF_X1 port map( D => n6632, CK => CLK, Q => 
                           n20405, QN => n14829);
   REGISTERS_reg_12_42_inst : DFF_X1 port map( D => n6631, CK => CLK, Q => 
                           n20404, QN => n14830);
   REGISTERS_reg_12_41_inst : DFF_X1 port map( D => n6630, CK => CLK, Q => 
                           n20403, QN => n14831);
   REGISTERS_reg_12_40_inst : DFF_X1 port map( D => n6629, CK => CLK, Q => 
                           n20402, QN => n14832);
   REGISTERS_reg_12_39_inst : DFF_X1 port map( D => n6628, CK => CLK, Q => 
                           n20401, QN => n14833);
   REGISTERS_reg_12_38_inst : DFF_X1 port map( D => n6627, CK => CLK, Q => 
                           n20400, QN => n14834);
   REGISTERS_reg_12_37_inst : DFF_X1 port map( D => n6626, CK => CLK, Q => 
                           n20399, QN => n14835);
   REGISTERS_reg_12_36_inst : DFF_X1 port map( D => n6625, CK => CLK, Q => 
                           n20398, QN => n14836);
   REGISTERS_reg_12_35_inst : DFF_X1 port map( D => n6624, CK => CLK, Q => 
                           n20397, QN => n14837);
   REGISTERS_reg_12_34_inst : DFF_X1 port map( D => n6623, CK => CLK, Q => 
                           n20396, QN => n14838);
   REGISTERS_reg_12_33_inst : DFF_X1 port map( D => n6622, CK => CLK, Q => 
                           n20395, QN => n14839);
   REGISTERS_reg_12_32_inst : DFF_X1 port map( D => n6621, CK => CLK, Q => 
                           n20394, QN => n14840);
   REGISTERS_reg_12_31_inst : DFF_X1 port map( D => n6620, CK => CLK, Q => 
                           n20393, QN => n14841);
   REGISTERS_reg_12_30_inst : DFF_X1 port map( D => n6619, CK => CLK, Q => 
                           n20392, QN => n14842);
   REGISTERS_reg_12_29_inst : DFF_X1 port map( D => n6618, CK => CLK, Q => 
                           n20391, QN => n14843);
   REGISTERS_reg_12_28_inst : DFF_X1 port map( D => n6617, CK => CLK, Q => 
                           n20390, QN => n14844);
   REGISTERS_reg_12_27_inst : DFF_X1 port map( D => n6616, CK => CLK, Q => 
                           n20389, QN => n14845);
   REGISTERS_reg_12_26_inst : DFF_X1 port map( D => n6615, CK => CLK, Q => 
                           n20388, QN => n14846);
   REGISTERS_reg_12_25_inst : DFF_X1 port map( D => n6614, CK => CLK, Q => 
                           n20387, QN => n14847);
   REGISTERS_reg_12_24_inst : DFF_X1 port map( D => n6613, CK => CLK, Q => 
                           n20386, QN => n14848);
   REGISTERS_reg_12_23_inst : DFF_X1 port map( D => n6612, CK => CLK, Q => 
                           n20385, QN => n14849);
   REGISTERS_reg_12_22_inst : DFF_X1 port map( D => n6611, CK => CLK, Q => 
                           n20384, QN => n14850);
   REGISTERS_reg_12_21_inst : DFF_X1 port map( D => n6610, CK => CLK, Q => 
                           n20383, QN => n14851);
   REGISTERS_reg_12_20_inst : DFF_X1 port map( D => n6609, CK => CLK, Q => 
                           n20382, QN => n14852);
   REGISTERS_reg_12_19_inst : DFF_X1 port map( D => n6608, CK => CLK, Q => 
                           n20381, QN => n14853);
   REGISTERS_reg_12_18_inst : DFF_X1 port map( D => n6607, CK => CLK, Q => 
                           n20380, QN => n14854);
   REGISTERS_reg_12_17_inst : DFF_X1 port map( D => n6606, CK => CLK, Q => 
                           n20379, QN => n14855);
   REGISTERS_reg_12_16_inst : DFF_X1 port map( D => n6605, CK => CLK, Q => 
                           n20378, QN => n14856);
   REGISTERS_reg_12_15_inst : DFF_X1 port map( D => n6604, CK => CLK, Q => 
                           n20377, QN => n14857);
   REGISTERS_reg_12_14_inst : DFF_X1 port map( D => n6603, CK => CLK, Q => 
                           n20376, QN => n14858);
   REGISTERS_reg_12_13_inst : DFF_X1 port map( D => n6602, CK => CLK, Q => 
                           n20375, QN => n14859);
   REGISTERS_reg_12_12_inst : DFF_X1 port map( D => n6601, CK => CLK, Q => 
                           n20374, QN => n14860);
   REGISTERS_reg_12_11_inst : DFF_X1 port map( D => n6600, CK => CLK, Q => 
                           n20373, QN => n14861);
   REGISTERS_reg_12_10_inst : DFF_X1 port map( D => n6599, CK => CLK, Q => 
                           n20372, QN => n14862);
   REGISTERS_reg_12_9_inst : DFF_X1 port map( D => n6598, CK => CLK, Q => 
                           n20371, QN => n14863);
   REGISTERS_reg_12_8_inst : DFF_X1 port map( D => n6597, CK => CLK, Q => 
                           n20370, QN => n14864);
   REGISTERS_reg_12_7_inst : DFF_X1 port map( D => n6596, CK => CLK, Q => 
                           n20369, QN => n14865);
   REGISTERS_reg_12_6_inst : DFF_X1 port map( D => n6595, CK => CLK, Q => 
                           n20368, QN => n14866);
   REGISTERS_reg_12_5_inst : DFF_X1 port map( D => n6594, CK => CLK, Q => 
                           n20367, QN => n14867);
   REGISTERS_reg_12_4_inst : DFF_X1 port map( D => n6593, CK => CLK, Q => 
                           n20366, QN => n14868);
   REGISTERS_reg_12_3_inst : DFF_X1 port map( D => n6592, CK => CLK, Q => 
                           n20365, QN => n14869);
   REGISTERS_reg_12_2_inst : DFF_X1 port map( D => n6591, CK => CLK, Q => 
                           n20364, QN => n14870);
   REGISTERS_reg_12_1_inst : DFF_X1 port map( D => n6590, CK => CLK, Q => 
                           n20363, QN => n14871);
   REGISTERS_reg_12_0_inst : DFF_X1 port map( D => n6589, CK => CLK, Q => 
                           n20362, QN => n14872);
   REGISTERS_reg_11_59_inst : DFF_X1 port map( D => n6712, CK => CLK, Q => 
                           n20361, QN => n14747);
   REGISTERS_reg_11_58_inst : DFF_X1 port map( D => n6711, CK => CLK, Q => 
                           n20360, QN => n14748);
   REGISTERS_reg_11_57_inst : DFF_X1 port map( D => n6710, CK => CLK, Q => 
                           n20359, QN => n14749);
   REGISTERS_reg_11_56_inst : DFF_X1 port map( D => n6709, CK => CLK, Q => 
                           n20358, QN => n14750);
   REGISTERS_reg_11_55_inst : DFF_X1 port map( D => n6708, CK => CLK, Q => 
                           n20357, QN => n14751);
   REGISTERS_reg_11_54_inst : DFF_X1 port map( D => n6707, CK => CLK, Q => 
                           n20356, QN => n14752);
   REGISTERS_reg_11_53_inst : DFF_X1 port map( D => n6706, CK => CLK, Q => 
                           n20355, QN => n14753);
   REGISTERS_reg_11_52_inst : DFF_X1 port map( D => n6705, CK => CLK, Q => 
                           n20354, QN => n14754);
   REGISTERS_reg_11_51_inst : DFF_X1 port map( D => n6704, CK => CLK, Q => 
                           n20353, QN => n14755);
   REGISTERS_reg_11_50_inst : DFF_X1 port map( D => n6703, CK => CLK, Q => 
                           n20352, QN => n14756);
   REGISTERS_reg_11_49_inst : DFF_X1 port map( D => n6702, CK => CLK, Q => 
                           n20351, QN => n14757);
   REGISTERS_reg_11_48_inst : DFF_X1 port map( D => n6701, CK => CLK, Q => 
                           n20350, QN => n14758);
   REGISTERS_reg_11_47_inst : DFF_X1 port map( D => n6700, CK => CLK, Q => 
                           n20349, QN => n14759);
   REGISTERS_reg_11_46_inst : DFF_X1 port map( D => n6699, CK => CLK, Q => 
                           n20348, QN => n14760);
   REGISTERS_reg_11_45_inst : DFF_X1 port map( D => n6698, CK => CLK, Q => 
                           n20347, QN => n14761);
   REGISTERS_reg_11_44_inst : DFF_X1 port map( D => n6697, CK => CLK, Q => 
                           n20346, QN => n14762);
   REGISTERS_reg_11_43_inst : DFF_X1 port map( D => n6696, CK => CLK, Q => 
                           n20345, QN => n14763);
   REGISTERS_reg_11_42_inst : DFF_X1 port map( D => n6695, CK => CLK, Q => 
                           n20344, QN => n14764);
   REGISTERS_reg_11_41_inst : DFF_X1 port map( D => n6694, CK => CLK, Q => 
                           n20343, QN => n14765);
   REGISTERS_reg_11_40_inst : DFF_X1 port map( D => n6693, CK => CLK, Q => 
                           n20342, QN => n14766);
   REGISTERS_reg_11_39_inst : DFF_X1 port map( D => n6692, CK => CLK, Q => 
                           n20341, QN => n14767);
   REGISTERS_reg_11_38_inst : DFF_X1 port map( D => n6691, CK => CLK, Q => 
                           n20340, QN => n14768);
   REGISTERS_reg_11_37_inst : DFF_X1 port map( D => n6690, CK => CLK, Q => 
                           n20339, QN => n14769);
   REGISTERS_reg_11_36_inst : DFF_X1 port map( D => n6689, CK => CLK, Q => 
                           n20338, QN => n14770);
   REGISTERS_reg_11_35_inst : DFF_X1 port map( D => n6688, CK => CLK, Q => 
                           n20337, QN => n14771);
   REGISTERS_reg_11_34_inst : DFF_X1 port map( D => n6687, CK => CLK, Q => 
                           n20336, QN => n14772);
   REGISTERS_reg_11_33_inst : DFF_X1 port map( D => n6686, CK => CLK, Q => 
                           n20335, QN => n14773);
   REGISTERS_reg_11_32_inst : DFF_X1 port map( D => n6685, CK => CLK, Q => 
                           n20334, QN => n14774);
   REGISTERS_reg_11_31_inst : DFF_X1 port map( D => n6684, CK => CLK, Q => 
                           n20333, QN => n14775);
   REGISTERS_reg_11_30_inst : DFF_X1 port map( D => n6683, CK => CLK, Q => 
                           n20332, QN => n14776);
   REGISTERS_reg_11_29_inst : DFF_X1 port map( D => n6682, CK => CLK, Q => 
                           n20331, QN => n14777);
   REGISTERS_reg_11_28_inst : DFF_X1 port map( D => n6681, CK => CLK, Q => 
                           n20330, QN => n14778);
   REGISTERS_reg_11_27_inst : DFF_X1 port map( D => n6680, CK => CLK, Q => 
                           n20329, QN => n14779);
   REGISTERS_reg_11_26_inst : DFF_X1 port map( D => n6679, CK => CLK, Q => 
                           n20328, QN => n14780);
   REGISTERS_reg_11_25_inst : DFF_X1 port map( D => n6678, CK => CLK, Q => 
                           n20327, QN => n14781);
   REGISTERS_reg_11_24_inst : DFF_X1 port map( D => n6677, CK => CLK, Q => 
                           n20326, QN => n14782);
   REGISTERS_reg_11_23_inst : DFF_X1 port map( D => n6676, CK => CLK, Q => 
                           n20325, QN => n14783);
   REGISTERS_reg_11_22_inst : DFF_X1 port map( D => n6675, CK => CLK, Q => 
                           n20324, QN => n14784);
   REGISTERS_reg_11_21_inst : DFF_X1 port map( D => n6674, CK => CLK, Q => 
                           n20323, QN => n14785);
   REGISTERS_reg_11_20_inst : DFF_X1 port map( D => n6673, CK => CLK, Q => 
                           n20322, QN => n14786);
   REGISTERS_reg_11_19_inst : DFF_X1 port map( D => n6672, CK => CLK, Q => 
                           n20321, QN => n14787);
   REGISTERS_reg_11_18_inst : DFF_X1 port map( D => n6671, CK => CLK, Q => 
                           n20320, QN => n14788);
   REGISTERS_reg_11_17_inst : DFF_X1 port map( D => n6670, CK => CLK, Q => 
                           n20319, QN => n14789);
   REGISTERS_reg_11_16_inst : DFF_X1 port map( D => n6669, CK => CLK, Q => 
                           n20318, QN => n14790);
   REGISTERS_reg_11_15_inst : DFF_X1 port map( D => n6668, CK => CLK, Q => 
                           n20317, QN => n14791);
   REGISTERS_reg_11_14_inst : DFF_X1 port map( D => n6667, CK => CLK, Q => 
                           n20316, QN => n14792);
   REGISTERS_reg_11_13_inst : DFF_X1 port map( D => n6666, CK => CLK, Q => 
                           n20315, QN => n14793);
   REGISTERS_reg_11_12_inst : DFF_X1 port map( D => n6665, CK => CLK, Q => 
                           n20314, QN => n14794);
   REGISTERS_reg_11_11_inst : DFF_X1 port map( D => n6664, CK => CLK, Q => 
                           n20313, QN => n14795);
   REGISTERS_reg_11_10_inst : DFF_X1 port map( D => n6663, CK => CLK, Q => 
                           n20312, QN => n14796);
   REGISTERS_reg_11_9_inst : DFF_X1 port map( D => n6662, CK => CLK, Q => 
                           n20311, QN => n14797);
   REGISTERS_reg_11_8_inst : DFF_X1 port map( D => n6661, CK => CLK, Q => 
                           n20310, QN => n14798);
   REGISTERS_reg_11_7_inst : DFF_X1 port map( D => n6660, CK => CLK, Q => 
                           n20309, QN => n14799);
   REGISTERS_reg_11_6_inst : DFF_X1 port map( D => n6659, CK => CLK, Q => 
                           n20308, QN => n14800);
   REGISTERS_reg_11_5_inst : DFF_X1 port map( D => n6658, CK => CLK, Q => 
                           n20307, QN => n14801);
   REGISTERS_reg_11_4_inst : DFF_X1 port map( D => n6657, CK => CLK, Q => 
                           n20306, QN => n14802);
   REGISTERS_reg_11_3_inst : DFF_X1 port map( D => n6656, CK => CLK, Q => 
                           n20305, QN => n14803);
   REGISTERS_reg_11_2_inst : DFF_X1 port map( D => n6655, CK => CLK, Q => 
                           n20304, QN => n14804);
   REGISTERS_reg_11_1_inst : DFF_X1 port map( D => n6654, CK => CLK, Q => 
                           n20303, QN => n14805);
   REGISTERS_reg_11_0_inst : DFF_X1 port map( D => n6653, CK => CLK, Q => 
                           n20302, QN => n14806);
   REGISTERS_reg_9_59_inst : DFF_X1 port map( D => n6840, CK => CLK, Q => n8975
                           , QN => n14614);
   REGISTERS_reg_9_58_inst : DFF_X1 port map( D => n6839, CK => CLK, Q => n8979
                           , QN => n14615);
   REGISTERS_reg_9_57_inst : DFF_X1 port map( D => n6838, CK => CLK, Q => n8983
                           , QN => n14616);
   REGISTERS_reg_9_56_inst : DFF_X1 port map( D => n6837, CK => CLK, Q => n8987
                           , QN => n14617);
   REGISTERS_reg_9_55_inst : DFF_X1 port map( D => n6836, CK => CLK, Q => n8991
                           , QN => n14618);
   REGISTERS_reg_9_54_inst : DFF_X1 port map( D => n6835, CK => CLK, Q => n8995
                           , QN => n14619);
   REGISTERS_reg_9_53_inst : DFF_X1 port map( D => n6834, CK => CLK, Q => n8999
                           , QN => n14620);
   REGISTERS_reg_9_52_inst : DFF_X1 port map( D => n6833, CK => CLK, Q => n9003
                           , QN => n14621);
   REGISTERS_reg_9_51_inst : DFF_X1 port map( D => n6832, CK => CLK, Q => n9007
                           , QN => n14622);
   REGISTERS_reg_9_50_inst : DFF_X1 port map( D => n6831, CK => CLK, Q => n9011
                           , QN => n14623);
   REGISTERS_reg_9_49_inst : DFF_X1 port map( D => n6830, CK => CLK, Q => n9015
                           , QN => n14624);
   REGISTERS_reg_9_48_inst : DFF_X1 port map( D => n6829, CK => CLK, Q => n9019
                           , QN => n14625);
   REGISTERS_reg_9_47_inst : DFF_X1 port map( D => n6828, CK => CLK, Q => n9023
                           , QN => n14626);
   REGISTERS_reg_9_46_inst : DFF_X1 port map( D => n6827, CK => CLK, Q => n9027
                           , QN => n14627);
   REGISTERS_reg_9_45_inst : DFF_X1 port map( D => n6826, CK => CLK, Q => n9031
                           , QN => n14628);
   REGISTERS_reg_9_44_inst : DFF_X1 port map( D => n6825, CK => CLK, Q => n9035
                           , QN => n14629);
   REGISTERS_reg_9_43_inst : DFF_X1 port map( D => n6824, CK => CLK, Q => n9039
                           , QN => n14630);
   REGISTERS_reg_9_42_inst : DFF_X1 port map( D => n6823, CK => CLK, Q => n9043
                           , QN => n14631);
   REGISTERS_reg_9_41_inst : DFF_X1 port map( D => n6822, CK => CLK, Q => n9047
                           , QN => n14632);
   REGISTERS_reg_9_40_inst : DFF_X1 port map( D => n6821, CK => CLK, Q => n9051
                           , QN => n14633);
   REGISTERS_reg_9_39_inst : DFF_X1 port map( D => n6820, CK => CLK, Q => n9055
                           , QN => n14634);
   REGISTERS_reg_9_38_inst : DFF_X1 port map( D => n6819, CK => CLK, Q => n9059
                           , QN => n14635);
   REGISTERS_reg_9_37_inst : DFF_X1 port map( D => n6818, CK => CLK, Q => n9063
                           , QN => n14636);
   REGISTERS_reg_9_36_inst : DFF_X1 port map( D => n6817, CK => CLK, Q => n9067
                           , QN => n14637);
   REGISTERS_reg_9_35_inst : DFF_X1 port map( D => n6816, CK => CLK, Q => n9071
                           , QN => n14638);
   REGISTERS_reg_9_34_inst : DFF_X1 port map( D => n6815, CK => CLK, Q => n9075
                           , QN => n14639);
   REGISTERS_reg_9_33_inst : DFF_X1 port map( D => n6814, CK => CLK, Q => n9079
                           , QN => n14640);
   REGISTERS_reg_9_32_inst : DFF_X1 port map( D => n6813, CK => CLK, Q => n9083
                           , QN => n14641);
   REGISTERS_reg_9_31_inst : DFF_X1 port map( D => n6812, CK => CLK, Q => n9087
                           , QN => n14642);
   REGISTERS_reg_9_30_inst : DFF_X1 port map( D => n6811, CK => CLK, Q => n9091
                           , QN => n14643);
   REGISTERS_reg_9_29_inst : DFF_X1 port map( D => n6810, CK => CLK, Q => n9095
                           , QN => n14644);
   REGISTERS_reg_9_28_inst : DFF_X1 port map( D => n6809, CK => CLK, Q => n9099
                           , QN => n14645);
   REGISTERS_reg_9_27_inst : DFF_X1 port map( D => n6808, CK => CLK, Q => n9103
                           , QN => n14646);
   REGISTERS_reg_9_26_inst : DFF_X1 port map( D => n6807, CK => CLK, Q => n9107
                           , QN => n14647);
   REGISTERS_reg_9_25_inst : DFF_X1 port map( D => n6806, CK => CLK, Q => n9111
                           , QN => n14648);
   REGISTERS_reg_9_24_inst : DFF_X1 port map( D => n6805, CK => CLK, Q => n9115
                           , QN => n14649);
   REGISTERS_reg_9_23_inst : DFF_X1 port map( D => n6804, CK => CLK, Q => n9119
                           , QN => n14650);
   REGISTERS_reg_9_22_inst : DFF_X1 port map( D => n6803, CK => CLK, Q => n9123
                           , QN => n14651);
   REGISTERS_reg_9_21_inst : DFF_X1 port map( D => n6802, CK => CLK, Q => n9127
                           , QN => n14652);
   REGISTERS_reg_9_20_inst : DFF_X1 port map( D => n6801, CK => CLK, Q => n9131
                           , QN => n14653);
   REGISTERS_reg_9_19_inst : DFF_X1 port map( D => n6800, CK => CLK, Q => n9135
                           , QN => n14654);
   REGISTERS_reg_9_18_inst : DFF_X1 port map( D => n6799, CK => CLK, Q => n9139
                           , QN => n14655);
   REGISTERS_reg_9_17_inst : DFF_X1 port map( D => n6798, CK => CLK, Q => n9143
                           , QN => n14656);
   REGISTERS_reg_9_16_inst : DFF_X1 port map( D => n6797, CK => CLK, Q => n9147
                           , QN => n14657);
   REGISTERS_reg_9_15_inst : DFF_X1 port map( D => n6796, CK => CLK, Q => n9151
                           , QN => n14658);
   REGISTERS_reg_9_14_inst : DFF_X1 port map( D => n6795, CK => CLK, Q => n9155
                           , QN => n14659);
   REGISTERS_reg_9_13_inst : DFF_X1 port map( D => n6794, CK => CLK, Q => n9159
                           , QN => n14660);
   REGISTERS_reg_9_12_inst : DFF_X1 port map( D => n6793, CK => CLK, Q => n9163
                           , QN => n14661);
   REGISTERS_reg_9_11_inst : DFF_X1 port map( D => n6792, CK => CLK, Q => n9167
                           , QN => n14662);
   REGISTERS_reg_9_10_inst : DFF_X1 port map( D => n6791, CK => CLK, Q => n9171
                           , QN => n14663);
   REGISTERS_reg_9_9_inst : DFF_X1 port map( D => n6790, CK => CLK, Q => n9175,
                           QN => n14664);
   REGISTERS_reg_9_8_inst : DFF_X1 port map( D => n6789, CK => CLK, Q => n9179,
                           QN => n14665);
   REGISTERS_reg_9_7_inst : DFF_X1 port map( D => n6788, CK => CLK, Q => n9183,
                           QN => n14666);
   REGISTERS_reg_9_6_inst : DFF_X1 port map( D => n6787, CK => CLK, Q => n9187,
                           QN => n14667);
   REGISTERS_reg_9_5_inst : DFF_X1 port map( D => n6786, CK => CLK, Q => n9191,
                           QN => n14668);
   REGISTERS_reg_9_4_inst : DFF_X1 port map( D => n6785, CK => CLK, Q => n9195,
                           QN => n14669);
   REGISTERS_reg_9_3_inst : DFF_X1 port map( D => n6784, CK => CLK, Q => n9199,
                           QN => n14670);
   REGISTERS_reg_9_2_inst : DFF_X1 port map( D => n6783, CK => CLK, Q => n9203,
                           QN => n14671);
   REGISTERS_reg_9_1_inst : DFF_X1 port map( D => n6782, CK => CLK, Q => n9207,
                           QN => n14672);
   REGISTERS_reg_9_0_inst : DFF_X1 port map( D => n6781, CK => CLK, Q => n9211,
                           QN => n14673);
   REGISTERS_reg_15_59_inst : DFF_X1 port map( D => n6456, CK => CLK, Q => 
                           n20301, QN => n15011);
   REGISTERS_reg_15_58_inst : DFF_X1 port map( D => n6455, CK => CLK, Q => 
                           n20300, QN => n15012);
   REGISTERS_reg_15_57_inst : DFF_X1 port map( D => n6454, CK => CLK, Q => 
                           n20299, QN => n15013);
   REGISTERS_reg_15_56_inst : DFF_X1 port map( D => n6453, CK => CLK, Q => 
                           n20298, QN => n15014);
   REGISTERS_reg_15_55_inst : DFF_X1 port map( D => n6452, CK => CLK, Q => 
                           n20297, QN => n15015);
   REGISTERS_reg_15_54_inst : DFF_X1 port map( D => n6451, CK => CLK, Q => 
                           n20296, QN => n15016);
   REGISTERS_reg_15_53_inst : DFF_X1 port map( D => n6450, CK => CLK, Q => 
                           n20295, QN => n15017);
   REGISTERS_reg_15_52_inst : DFF_X1 port map( D => n6449, CK => CLK, Q => 
                           n20294, QN => n15018);
   REGISTERS_reg_15_51_inst : DFF_X1 port map( D => n6448, CK => CLK, Q => 
                           n20293, QN => n15019);
   REGISTERS_reg_15_50_inst : DFF_X1 port map( D => n6447, CK => CLK, Q => 
                           n20292, QN => n15020);
   REGISTERS_reg_15_49_inst : DFF_X1 port map( D => n6446, CK => CLK, Q => 
                           n20291, QN => n15021);
   REGISTERS_reg_15_48_inst : DFF_X1 port map( D => n6445, CK => CLK, Q => 
                           n20290, QN => n15022);
   REGISTERS_reg_15_47_inst : DFF_X1 port map( D => n6444, CK => CLK, Q => 
                           n20289, QN => n15023);
   REGISTERS_reg_15_46_inst : DFF_X1 port map( D => n6443, CK => CLK, Q => 
                           n20288, QN => n15024);
   REGISTERS_reg_15_45_inst : DFF_X1 port map( D => n6442, CK => CLK, Q => 
                           n20287, QN => n15025);
   REGISTERS_reg_15_44_inst : DFF_X1 port map( D => n6441, CK => CLK, Q => 
                           n20286, QN => n15026);
   REGISTERS_reg_15_43_inst : DFF_X1 port map( D => n6440, CK => CLK, Q => 
                           n20285, QN => n15027);
   REGISTERS_reg_15_42_inst : DFF_X1 port map( D => n6439, CK => CLK, Q => 
                           n20284, QN => n15028);
   REGISTERS_reg_15_41_inst : DFF_X1 port map( D => n6438, CK => CLK, Q => 
                           n20283, QN => n15029);
   REGISTERS_reg_15_40_inst : DFF_X1 port map( D => n6437, CK => CLK, Q => 
                           n20282, QN => n15030);
   REGISTERS_reg_15_39_inst : DFF_X1 port map( D => n6436, CK => CLK, Q => 
                           n20281, QN => n15031);
   REGISTERS_reg_15_38_inst : DFF_X1 port map( D => n6435, CK => CLK, Q => 
                           n20280, QN => n15032);
   REGISTERS_reg_15_37_inst : DFF_X1 port map( D => n6434, CK => CLK, Q => 
                           n20279, QN => n15033);
   REGISTERS_reg_15_36_inst : DFF_X1 port map( D => n6433, CK => CLK, Q => 
                           n20278, QN => n15034);
   REGISTERS_reg_15_35_inst : DFF_X1 port map( D => n6432, CK => CLK, Q => 
                           n20277, QN => n15035);
   REGISTERS_reg_15_34_inst : DFF_X1 port map( D => n6431, CK => CLK, Q => 
                           n20276, QN => n15036);
   REGISTERS_reg_15_33_inst : DFF_X1 port map( D => n6430, CK => CLK, Q => 
                           n20275, QN => n15037);
   REGISTERS_reg_15_32_inst : DFF_X1 port map( D => n6429, CK => CLK, Q => 
                           n20274, QN => n15038);
   REGISTERS_reg_15_31_inst : DFF_X1 port map( D => n6428, CK => CLK, Q => 
                           n20273, QN => n15039);
   REGISTERS_reg_15_30_inst : DFF_X1 port map( D => n6427, CK => CLK, Q => 
                           n20272, QN => n15040);
   REGISTERS_reg_15_29_inst : DFF_X1 port map( D => n6426, CK => CLK, Q => 
                           n20271, QN => n15041);
   REGISTERS_reg_15_28_inst : DFF_X1 port map( D => n6425, CK => CLK, Q => 
                           n20270, QN => n15042);
   REGISTERS_reg_15_27_inst : DFF_X1 port map( D => n6424, CK => CLK, Q => 
                           n20269, QN => n15043);
   REGISTERS_reg_15_26_inst : DFF_X1 port map( D => n6423, CK => CLK, Q => 
                           n20268, QN => n15044);
   REGISTERS_reg_15_25_inst : DFF_X1 port map( D => n6422, CK => CLK, Q => 
                           n20267, QN => n15045);
   REGISTERS_reg_15_24_inst : DFF_X1 port map( D => n6421, CK => CLK, Q => 
                           n20266, QN => n15046);
   REGISTERS_reg_15_23_inst : DFF_X1 port map( D => n6420, CK => CLK, Q => 
                           n20265, QN => n15047);
   REGISTERS_reg_15_22_inst : DFF_X1 port map( D => n6419, CK => CLK, Q => 
                           n20264, QN => n15048);
   REGISTERS_reg_15_21_inst : DFF_X1 port map( D => n6418, CK => CLK, Q => 
                           n20263, QN => n15049);
   REGISTERS_reg_15_20_inst : DFF_X1 port map( D => n6417, CK => CLK, Q => 
                           n20262, QN => n15050);
   REGISTERS_reg_15_19_inst : DFF_X1 port map( D => n6416, CK => CLK, Q => 
                           n20261, QN => n15051);
   REGISTERS_reg_15_18_inst : DFF_X1 port map( D => n6415, CK => CLK, Q => 
                           n20260, QN => n15052);
   REGISTERS_reg_15_17_inst : DFF_X1 port map( D => n6414, CK => CLK, Q => 
                           n20259, QN => n15053);
   REGISTERS_reg_15_16_inst : DFF_X1 port map( D => n6413, CK => CLK, Q => 
                           n20258, QN => n15054);
   REGISTERS_reg_15_15_inst : DFF_X1 port map( D => n6412, CK => CLK, Q => 
                           n20257, QN => n15055);
   REGISTERS_reg_15_14_inst : DFF_X1 port map( D => n6411, CK => CLK, Q => 
                           n20256, QN => n15056);
   REGISTERS_reg_15_13_inst : DFF_X1 port map( D => n6410, CK => CLK, Q => 
                           n20255, QN => n15057);
   REGISTERS_reg_15_12_inst : DFF_X1 port map( D => n6409, CK => CLK, Q => 
                           n20254, QN => n15058);
   REGISTERS_reg_15_11_inst : DFF_X1 port map( D => n6408, CK => CLK, Q => 
                           n20253, QN => n15059);
   REGISTERS_reg_15_10_inst : DFF_X1 port map( D => n6407, CK => CLK, Q => 
                           n20252, QN => n15060);
   REGISTERS_reg_15_9_inst : DFF_X1 port map( D => n6406, CK => CLK, Q => 
                           n20251, QN => n15061);
   REGISTERS_reg_15_8_inst : DFF_X1 port map( D => n6405, CK => CLK, Q => 
                           n20250, QN => n15062);
   REGISTERS_reg_15_7_inst : DFF_X1 port map( D => n6404, CK => CLK, Q => 
                           n20249, QN => n15063);
   REGISTERS_reg_15_6_inst : DFF_X1 port map( D => n6403, CK => CLK, Q => 
                           n20248, QN => n15064);
   REGISTERS_reg_15_5_inst : DFF_X1 port map( D => n6402, CK => CLK, Q => 
                           n20247, QN => n15065);
   REGISTERS_reg_15_4_inst : DFF_X1 port map( D => n6401, CK => CLK, Q => 
                           n20246, QN => n15066);
   REGISTERS_reg_15_3_inst : DFF_X1 port map( D => n6400, CK => CLK, Q => 
                           n20245, QN => n15067);
   REGISTERS_reg_15_2_inst : DFF_X1 port map( D => n6399, CK => CLK, Q => 
                           n20244, QN => n15068);
   REGISTERS_reg_15_1_inst : DFF_X1 port map( D => n6398, CK => CLK, Q => 
                           n20243, QN => n15069);
   REGISTERS_reg_15_0_inst : DFF_X1 port map( D => n6397, CK => CLK, Q => 
                           n20242, QN => n15070);
   REGISTERS_reg_13_59_inst : DFF_X1 port map( D => n6584, CK => CLK, Q => 
                           n8592, QN => n14879);
   REGISTERS_reg_13_58_inst : DFF_X1 port map( D => n6583, CK => CLK, Q => 
                           n8596, QN => n14880);
   REGISTERS_reg_13_57_inst : DFF_X1 port map( D => n6582, CK => CLK, Q => 
                           n8600, QN => n14881);
   REGISTERS_reg_13_56_inst : DFF_X1 port map( D => n6581, CK => CLK, Q => 
                           n8604, QN => n14882);
   REGISTERS_reg_13_55_inst : DFF_X1 port map( D => n6580, CK => CLK, Q => 
                           n8608, QN => n14883);
   REGISTERS_reg_13_54_inst : DFF_X1 port map( D => n6579, CK => CLK, Q => 
                           n8612, QN => n14884);
   REGISTERS_reg_13_53_inst : DFF_X1 port map( D => n6578, CK => CLK, Q => 
                           n8616, QN => n14885);
   REGISTERS_reg_13_52_inst : DFF_X1 port map( D => n6577, CK => CLK, Q => 
                           n8620, QN => n14886);
   REGISTERS_reg_13_51_inst : DFF_X1 port map( D => n6576, CK => CLK, Q => 
                           n8624, QN => n14887);
   REGISTERS_reg_13_50_inst : DFF_X1 port map( D => n6575, CK => CLK, Q => 
                           n8628, QN => n14888);
   REGISTERS_reg_13_49_inst : DFF_X1 port map( D => n6574, CK => CLK, Q => 
                           n8632, QN => n14889);
   REGISTERS_reg_13_48_inst : DFF_X1 port map( D => n6573, CK => CLK, Q => 
                           n8636, QN => n14890);
   REGISTERS_reg_13_47_inst : DFF_X1 port map( D => n6572, CK => CLK, Q => 
                           n8640, QN => n14891);
   REGISTERS_reg_13_46_inst : DFF_X1 port map( D => n6571, CK => CLK, Q => 
                           n8644, QN => n14892);
   REGISTERS_reg_13_45_inst : DFF_X1 port map( D => n6570, CK => CLK, Q => 
                           n8648, QN => n14893);
   REGISTERS_reg_13_44_inst : DFF_X1 port map( D => n6569, CK => CLK, Q => 
                           n8652, QN => n14894);
   REGISTERS_reg_13_43_inst : DFF_X1 port map( D => n6568, CK => CLK, Q => 
                           n8656, QN => n14895);
   REGISTERS_reg_13_42_inst : DFF_X1 port map( D => n6567, CK => CLK, Q => 
                           n8660, QN => n14896);
   REGISTERS_reg_13_41_inst : DFF_X1 port map( D => n6566, CK => CLK, Q => 
                           n8664, QN => n14897);
   REGISTERS_reg_13_40_inst : DFF_X1 port map( D => n6565, CK => CLK, Q => 
                           n8668, QN => n14898);
   REGISTERS_reg_13_39_inst : DFF_X1 port map( D => n6564, CK => CLK, Q => 
                           n8672, QN => n14899);
   REGISTERS_reg_13_38_inst : DFF_X1 port map( D => n6563, CK => CLK, Q => 
                           n8676, QN => n14900);
   REGISTERS_reg_13_37_inst : DFF_X1 port map( D => n6562, CK => CLK, Q => 
                           n8680, QN => n14901);
   REGISTERS_reg_13_36_inst : DFF_X1 port map( D => n6561, CK => CLK, Q => 
                           n8684, QN => n14902);
   REGISTERS_reg_13_35_inst : DFF_X1 port map( D => n6560, CK => CLK, Q => 
                           n8688, QN => n14903);
   REGISTERS_reg_13_34_inst : DFF_X1 port map( D => n6559, CK => CLK, Q => 
                           n8692, QN => n14904);
   REGISTERS_reg_13_33_inst : DFF_X1 port map( D => n6558, CK => CLK, Q => 
                           n8696, QN => n14905);
   REGISTERS_reg_13_32_inst : DFF_X1 port map( D => n6557, CK => CLK, Q => 
                           n8700, QN => n14906);
   REGISTERS_reg_13_31_inst : DFF_X1 port map( D => n6556, CK => CLK, Q => 
                           n8704, QN => n14907);
   REGISTERS_reg_13_30_inst : DFF_X1 port map( D => n6555, CK => CLK, Q => 
                           n8708, QN => n14908);
   REGISTERS_reg_13_29_inst : DFF_X1 port map( D => n6554, CK => CLK, Q => 
                           n8712, QN => n14909);
   REGISTERS_reg_13_28_inst : DFF_X1 port map( D => n6553, CK => CLK, Q => 
                           n8716, QN => n14910);
   REGISTERS_reg_13_27_inst : DFF_X1 port map( D => n6552, CK => CLK, Q => 
                           n8720, QN => n14911);
   REGISTERS_reg_13_26_inst : DFF_X1 port map( D => n6551, CK => CLK, Q => 
                           n8724, QN => n14912);
   REGISTERS_reg_13_25_inst : DFF_X1 port map( D => n6550, CK => CLK, Q => 
                           n8728, QN => n14913);
   REGISTERS_reg_13_24_inst : DFF_X1 port map( D => n6549, CK => CLK, Q => 
                           n8732, QN => n14914);
   REGISTERS_reg_13_23_inst : DFF_X1 port map( D => n6548, CK => CLK, Q => 
                           n8736, QN => n14915);
   REGISTERS_reg_13_22_inst : DFF_X1 port map( D => n6547, CK => CLK, Q => 
                           n8740, QN => n14916);
   REGISTERS_reg_13_21_inst : DFF_X1 port map( D => n6546, CK => CLK, Q => 
                           n8744, QN => n14917);
   REGISTERS_reg_13_20_inst : DFF_X1 port map( D => n6545, CK => CLK, Q => 
                           n8748, QN => n14918);
   REGISTERS_reg_13_19_inst : DFF_X1 port map( D => n6544, CK => CLK, Q => 
                           n8752, QN => n14919);
   REGISTERS_reg_13_18_inst : DFF_X1 port map( D => n6543, CK => CLK, Q => 
                           n8756, QN => n14920);
   REGISTERS_reg_13_17_inst : DFF_X1 port map( D => n6542, CK => CLK, Q => 
                           n8760, QN => n14921);
   REGISTERS_reg_13_16_inst : DFF_X1 port map( D => n6541, CK => CLK, Q => 
                           n8764, QN => n14922);
   REGISTERS_reg_13_15_inst : DFF_X1 port map( D => n6540, CK => CLK, Q => 
                           n8768, QN => n14923);
   REGISTERS_reg_13_14_inst : DFF_X1 port map( D => n6539, CK => CLK, Q => 
                           n8772, QN => n14924);
   REGISTERS_reg_13_13_inst : DFF_X1 port map( D => n6538, CK => CLK, Q => 
                           n8776, QN => n14925);
   REGISTERS_reg_13_12_inst : DFF_X1 port map( D => n6537, CK => CLK, Q => 
                           n8780, QN => n14926);
   REGISTERS_reg_13_11_inst : DFF_X1 port map( D => n6536, CK => CLK, Q => 
                           n8784, QN => n14927);
   REGISTERS_reg_13_10_inst : DFF_X1 port map( D => n6535, CK => CLK, Q => 
                           n8788, QN => n14928);
   REGISTERS_reg_13_9_inst : DFF_X1 port map( D => n6534, CK => CLK, Q => n8792
                           , QN => n14929);
   REGISTERS_reg_13_8_inst : DFF_X1 port map( D => n6533, CK => CLK, Q => n8796
                           , QN => n14930);
   REGISTERS_reg_13_7_inst : DFF_X1 port map( D => n6532, CK => CLK, Q => n8800
                           , QN => n14931);
   REGISTERS_reg_13_6_inst : DFF_X1 port map( D => n6531, CK => CLK, Q => n8804
                           , QN => n14932);
   REGISTERS_reg_13_5_inst : DFF_X1 port map( D => n6530, CK => CLK, Q => n8808
                           , QN => n14933);
   REGISTERS_reg_13_4_inst : DFF_X1 port map( D => n6529, CK => CLK, Q => n8812
                           , QN => n14934);
   REGISTERS_reg_13_3_inst : DFF_X1 port map( D => n6528, CK => CLK, Q => n8816
                           , QN => n14935);
   REGISTERS_reg_13_2_inst : DFF_X1 port map( D => n6527, CK => CLK, Q => n8820
                           , QN => n14936);
   REGISTERS_reg_13_1_inst : DFF_X1 port map( D => n6526, CK => CLK, Q => n8824
                           , QN => n14937);
   REGISTERS_reg_13_0_inst : DFF_X1 port map( D => n6525, CK => CLK, Q => n8828
                           , QN => n14938);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n7352, CK => CLK, Q => 
                           n20241, QN => n14078);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n7351, CK => CLK, Q => 
                           n20240, QN => n14079);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n7350, CK => CLK, Q => 
                           n20239, QN => n14080);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n7349, CK => CLK, Q => 
                           n20238, QN => n14081);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n7348, CK => CLK, Q => 
                           n20237, QN => n14082);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n7347, CK => CLK, Q => 
                           n20236, QN => n14083);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n7346, CK => CLK, Q => 
                           n20235, QN => n14084);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n7345, CK => CLK, Q => 
                           n20234, QN => n14085);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n7344, CK => CLK, Q => 
                           n20233, QN => n14086);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n7343, CK => CLK, Q => 
                           n20232, QN => n14087);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n7342, CK => CLK, Q => 
                           n20231, QN => n14088);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n7341, CK => CLK, Q => 
                           n20230, QN => n14089);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n7340, CK => CLK, Q => 
                           n20229, QN => n14090);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n7339, CK => CLK, Q => 
                           n20228, QN => n14091);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n7338, CK => CLK, Q => 
                           n20227, QN => n14092);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n7337, CK => CLK, Q => 
                           n20226, QN => n14093);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n7336, CK => CLK, Q => 
                           n20225, QN => n14094);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n7335, CK => CLK, Q => 
                           n20224, QN => n14095);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n7334, CK => CLK, Q => 
                           n20223, QN => n14096);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n7333, CK => CLK, Q => 
                           n20222, QN => n14097);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n7332, CK => CLK, Q => 
                           n20221, QN => n14098);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n7331, CK => CLK, Q => 
                           n20220, QN => n14099);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n7330, CK => CLK, Q => 
                           n20219, QN => n14100);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n7329, CK => CLK, Q => 
                           n20218, QN => n14101);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n7328, CK => CLK, Q => 
                           n20217, QN => n14102);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n7327, CK => CLK, Q => 
                           n20216, QN => n14103);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n7326, CK => CLK, Q => 
                           n20215, QN => n14104);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n7325, CK => CLK, Q => 
                           n20214, QN => n14105);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n7324, CK => CLK, Q => 
                           n20213, QN => n14106);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n7323, CK => CLK, Q => 
                           n20212, QN => n14107);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n7322, CK => CLK, Q => 
                           n20211, QN => n14108);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n7321, CK => CLK, Q => 
                           n20210, QN => n14109);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n7320, CK => CLK, Q => 
                           n20209, QN => n14110);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n7319, CK => CLK, Q => 
                           n20208, QN => n14111);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n7318, CK => CLK, Q => 
                           n20207, QN => n14112);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n7317, CK => CLK, Q => 
                           n20206, QN => n14113);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n7316, CK => CLK, Q => 
                           n20205, QN => n14114);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n7315, CK => CLK, Q => 
                           n20204, QN => n14115);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n7314, CK => CLK, Q => 
                           n20203, QN => n14116);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n7313, CK => CLK, Q => 
                           n20202, QN => n14117);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n7312, CK => CLK, Q => 
                           n20201, QN => n14118);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n7311, CK => CLK, Q => 
                           n20200, QN => n14119);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n7310, CK => CLK, Q => 
                           n20199, QN => n14120);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n7309, CK => CLK, Q => 
                           n20198, QN => n14121);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n7308, CK => CLK, Q => 
                           n20197, QN => n14122);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n7307, CK => CLK, Q => 
                           n20196, QN => n14123);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n7306, CK => CLK, Q => 
                           n20195, QN => n14124);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n7305, CK => CLK, Q => 
                           n20194, QN => n14125);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n7304, CK => CLK, Q => 
                           n20193, QN => n14126);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n7303, CK => CLK, Q => 
                           n20192, QN => n14127);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n7302, CK => CLK, Q => n20191
                           , QN => n14128);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n7301, CK => CLK, Q => n20190
                           , QN => n14129);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n7300, CK => CLK, Q => n20189
                           , QN => n14130);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n7299, CK => CLK, Q => n20188
                           , QN => n14131);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n7298, CK => CLK, Q => n20187
                           , QN => n14132);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n7297, CK => CLK, Q => n20186
                           , QN => n14133);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n7296, CK => CLK, Q => n20185
                           , QN => n14134);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n7295, CK => CLK, Q => n20184
                           , QN => n14135);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n7294, CK => CLK, Q => n20183
                           , QN => n14136);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n7293, CK => CLK, Q => n20182
                           , QN => n14137);
   REGISTERS_reg_30_59_inst : DFF_X1 port map( D => n5496, CK => CLK, Q => 
                           n20181, QN => n16009);
   REGISTERS_reg_30_58_inst : DFF_X1 port map( D => n5495, CK => CLK, Q => 
                           n20180, QN => n16010);
   REGISTERS_reg_30_57_inst : DFF_X1 port map( D => n5494, CK => CLK, Q => 
                           n20179, QN => n16011);
   REGISTERS_reg_30_56_inst : DFF_X1 port map( D => n5493, CK => CLK, Q => 
                           n20178, QN => n16012);
   REGISTERS_reg_30_55_inst : DFF_X1 port map( D => n5492, CK => CLK, Q => 
                           n20177, QN => n16013);
   REGISTERS_reg_30_54_inst : DFF_X1 port map( D => n5491, CK => CLK, Q => 
                           n20176, QN => n16014);
   REGISTERS_reg_30_53_inst : DFF_X1 port map( D => n5490, CK => CLK, Q => 
                           n20175, QN => n16015);
   REGISTERS_reg_30_52_inst : DFF_X1 port map( D => n5489, CK => CLK, Q => 
                           n20174, QN => n16016);
   REGISTERS_reg_30_51_inst : DFF_X1 port map( D => n5488, CK => CLK, Q => 
                           n20173, QN => n16017);
   REGISTERS_reg_30_50_inst : DFF_X1 port map( D => n5487, CK => CLK, Q => 
                           n20172, QN => n16018);
   REGISTERS_reg_30_49_inst : DFF_X1 port map( D => n5486, CK => CLK, Q => 
                           n20171, QN => n16019);
   REGISTERS_reg_30_48_inst : DFF_X1 port map( D => n5485, CK => CLK, Q => 
                           n20170, QN => n16020);
   REGISTERS_reg_30_47_inst : DFF_X1 port map( D => n5484, CK => CLK, Q => 
                           n20169, QN => n16021);
   REGISTERS_reg_30_46_inst : DFF_X1 port map( D => n5483, CK => CLK, Q => 
                           n20168, QN => n16022);
   REGISTERS_reg_30_45_inst : DFF_X1 port map( D => n5482, CK => CLK, Q => 
                           n20167, QN => n16023);
   REGISTERS_reg_30_44_inst : DFF_X1 port map( D => n5481, CK => CLK, Q => 
                           n20166, QN => n16024);
   REGISTERS_reg_30_43_inst : DFF_X1 port map( D => n5480, CK => CLK, Q => 
                           n20165, QN => n16025);
   REGISTERS_reg_30_42_inst : DFF_X1 port map( D => n5479, CK => CLK, Q => 
                           n20164, QN => n16026);
   REGISTERS_reg_30_41_inst : DFF_X1 port map( D => n5478, CK => CLK, Q => 
                           n20163, QN => n16027);
   REGISTERS_reg_30_40_inst : DFF_X1 port map( D => n5477, CK => CLK, Q => 
                           n20162, QN => n16028);
   REGISTERS_reg_30_39_inst : DFF_X1 port map( D => n5476, CK => CLK, Q => 
                           n20161, QN => n16029);
   REGISTERS_reg_30_38_inst : DFF_X1 port map( D => n5475, CK => CLK, Q => 
                           n20160, QN => n16030);
   REGISTERS_reg_30_37_inst : DFF_X1 port map( D => n5474, CK => CLK, Q => 
                           n20159, QN => n16031);
   REGISTERS_reg_30_36_inst : DFF_X1 port map( D => n5473, CK => CLK, Q => 
                           n20158, QN => n16032);
   REGISTERS_reg_30_35_inst : DFF_X1 port map( D => n5472, CK => CLK, Q => 
                           n20157, QN => n16033);
   REGISTERS_reg_30_34_inst : DFF_X1 port map( D => n5471, CK => CLK, Q => 
                           n20156, QN => n16034);
   REGISTERS_reg_30_33_inst : DFF_X1 port map( D => n5470, CK => CLK, Q => 
                           n20155, QN => n16035);
   REGISTERS_reg_30_32_inst : DFF_X1 port map( D => n5469, CK => CLK, Q => 
                           n20154, QN => n16036);
   REGISTERS_reg_30_31_inst : DFF_X1 port map( D => n5468, CK => CLK, Q => 
                           n20153, QN => n16037);
   REGISTERS_reg_30_30_inst : DFF_X1 port map( D => n5467, CK => CLK, Q => 
                           n20152, QN => n16038);
   REGISTERS_reg_30_29_inst : DFF_X1 port map( D => n5466, CK => CLK, Q => 
                           n20151, QN => n16039);
   REGISTERS_reg_30_28_inst : DFF_X1 port map( D => n5465, CK => CLK, Q => 
                           n20150, QN => n16040);
   REGISTERS_reg_30_27_inst : DFF_X1 port map( D => n5464, CK => CLK, Q => 
                           n20149, QN => n16041);
   REGISTERS_reg_30_26_inst : DFF_X1 port map( D => n5463, CK => CLK, Q => 
                           n20148, QN => n16042);
   REGISTERS_reg_30_25_inst : DFF_X1 port map( D => n5462, CK => CLK, Q => 
                           n20147, QN => n16043);
   REGISTERS_reg_30_24_inst : DFF_X1 port map( D => n5461, CK => CLK, Q => 
                           n20146, QN => n16044);
   REGISTERS_reg_30_23_inst : DFF_X1 port map( D => n5460, CK => CLK, Q => 
                           n20145, QN => n16045);
   REGISTERS_reg_30_22_inst : DFF_X1 port map( D => n5459, CK => CLK, Q => 
                           n20144, QN => n16046);
   REGISTERS_reg_30_21_inst : DFF_X1 port map( D => n5458, CK => CLK, Q => 
                           n20143, QN => n16047);
   REGISTERS_reg_30_20_inst : DFF_X1 port map( D => n5457, CK => CLK, Q => 
                           n20142, QN => n16048);
   REGISTERS_reg_30_19_inst : DFF_X1 port map( D => n5456, CK => CLK, Q => 
                           n20141, QN => n16049);
   REGISTERS_reg_30_18_inst : DFF_X1 port map( D => n5455, CK => CLK, Q => 
                           n20140, QN => n16050);
   REGISTERS_reg_30_17_inst : DFF_X1 port map( D => n5454, CK => CLK, Q => 
                           n20139, QN => n16051);
   REGISTERS_reg_30_16_inst : DFF_X1 port map( D => n5453, CK => CLK, Q => 
                           n20138, QN => n16052);
   REGISTERS_reg_30_15_inst : DFF_X1 port map( D => n5452, CK => CLK, Q => 
                           n20137, QN => n16053);
   REGISTERS_reg_30_14_inst : DFF_X1 port map( D => n5451, CK => CLK, Q => 
                           n20136, QN => n16054);
   REGISTERS_reg_30_13_inst : DFF_X1 port map( D => n5450, CK => CLK, Q => 
                           n20135, QN => n16055);
   REGISTERS_reg_30_12_inst : DFF_X1 port map( D => n5449, CK => CLK, Q => 
                           n20134, QN => n16056);
   REGISTERS_reg_30_11_inst : DFF_X1 port map( D => n5448, CK => CLK, Q => 
                           n20133, QN => n16057);
   REGISTERS_reg_30_10_inst : DFF_X1 port map( D => n5447, CK => CLK, Q => 
                           n20132, QN => n16058);
   REGISTERS_reg_30_9_inst : DFF_X1 port map( D => n5446, CK => CLK, Q => 
                           n20131, QN => n16059);
   REGISTERS_reg_30_8_inst : DFF_X1 port map( D => n5445, CK => CLK, Q => 
                           n20130, QN => n16060);
   REGISTERS_reg_30_7_inst : DFF_X1 port map( D => n5444, CK => CLK, Q => 
                           n20129, QN => n16061);
   REGISTERS_reg_30_6_inst : DFF_X1 port map( D => n5443, CK => CLK, Q => 
                           n20128, QN => n16062);
   REGISTERS_reg_30_5_inst : DFF_X1 port map( D => n5442, CK => CLK, Q => 
                           n20127, QN => n16063);
   REGISTERS_reg_30_4_inst : DFF_X1 port map( D => n5441, CK => CLK, Q => 
                           n20126, QN => n16064);
   REGISTERS_reg_30_3_inst : DFF_X1 port map( D => n5440, CK => CLK, Q => 
                           n20125, QN => n16065);
   REGISTERS_reg_30_2_inst : DFF_X1 port map( D => n5439, CK => CLK, Q => 
                           n20124, QN => n16066);
   REGISTERS_reg_30_1_inst : DFF_X1 port map( D => n5438, CK => CLK, Q => 
                           n20123, QN => n16067);
   REGISTERS_reg_30_0_inst : DFF_X1 port map( D => n5437, CK => CLK, Q => 
                           n20122, QN => n16068);
   REGISTERS_reg_29_59_inst : DFF_X1 port map( D => n5560, CK => CLK, Q => 
                           n18628, QN => n15943);
   REGISTERS_reg_29_58_inst : DFF_X1 port map( D => n5559, CK => CLK, Q => 
                           n18648, QN => n15944);
   REGISTERS_reg_29_57_inst : DFF_X1 port map( D => n5558, CK => CLK, Q => 
                           n18668, QN => n15945);
   REGISTERS_reg_29_56_inst : DFF_X1 port map( D => n5557, CK => CLK, Q => 
                           n18688, QN => n15946);
   REGISTERS_reg_29_55_inst : DFF_X1 port map( D => n5556, CK => CLK, Q => 
                           n18708, QN => n15947);
   REGISTERS_reg_29_54_inst : DFF_X1 port map( D => n5555, CK => CLK, Q => 
                           n18728, QN => n15948);
   REGISTERS_reg_29_53_inst : DFF_X1 port map( D => n5554, CK => CLK, Q => 
                           n18748, QN => n15949);
   REGISTERS_reg_29_52_inst : DFF_X1 port map( D => n5553, CK => CLK, Q => 
                           n18768, QN => n15950);
   REGISTERS_reg_29_51_inst : DFF_X1 port map( D => n5552, CK => CLK, Q => 
                           n18788, QN => n15951);
   REGISTERS_reg_29_50_inst : DFF_X1 port map( D => n5551, CK => CLK, Q => 
                           n18808, QN => n15952);
   REGISTERS_reg_29_49_inst : DFF_X1 port map( D => n5550, CK => CLK, Q => 
                           n18828, QN => n15953);
   REGISTERS_reg_29_48_inst : DFF_X1 port map( D => n5549, CK => CLK, Q => 
                           n18848, QN => n15954);
   REGISTERS_reg_29_47_inst : DFF_X1 port map( D => n5548, CK => CLK, Q => 
                           n18868, QN => n15955);
   REGISTERS_reg_29_46_inst : DFF_X1 port map( D => n5547, CK => CLK, Q => 
                           n18888, QN => n15956);
   REGISTERS_reg_29_45_inst : DFF_X1 port map( D => n5546, CK => CLK, Q => 
                           n18908, QN => n15957);
   REGISTERS_reg_29_44_inst : DFF_X1 port map( D => n5545, CK => CLK, Q => 
                           n18928, QN => n15958);
   REGISTERS_reg_29_43_inst : DFF_X1 port map( D => n5544, CK => CLK, Q => 
                           n18948, QN => n15959);
   REGISTERS_reg_29_42_inst : DFF_X1 port map( D => n5543, CK => CLK, Q => 
                           n18968, QN => n15960);
   REGISTERS_reg_29_41_inst : DFF_X1 port map( D => n5542, CK => CLK, Q => 
                           n18988, QN => n15961);
   REGISTERS_reg_29_40_inst : DFF_X1 port map( D => n5541, CK => CLK, Q => 
                           n19008, QN => n15962);
   REGISTERS_reg_29_39_inst : DFF_X1 port map( D => n5540, CK => CLK, Q => 
                           n19028, QN => n15963);
   REGISTERS_reg_29_38_inst : DFF_X1 port map( D => n5539, CK => CLK, Q => 
                           n19048, QN => n15964);
   REGISTERS_reg_29_37_inst : DFF_X1 port map( D => n5538, CK => CLK, Q => 
                           n19068, QN => n15965);
   REGISTERS_reg_29_36_inst : DFF_X1 port map( D => n5537, CK => CLK, Q => 
                           n19088, QN => n15966);
   REGISTERS_reg_29_35_inst : DFF_X1 port map( D => n5536, CK => CLK, Q => 
                           n19108, QN => n15967);
   REGISTERS_reg_29_34_inst : DFF_X1 port map( D => n5535, CK => CLK, Q => 
                           n19128, QN => n15968);
   REGISTERS_reg_29_33_inst : DFF_X1 port map( D => n5534, CK => CLK, Q => 
                           n19148, QN => n15969);
   REGISTERS_reg_29_32_inst : DFF_X1 port map( D => n5533, CK => CLK, Q => 
                           n19168, QN => n15970);
   REGISTERS_reg_29_31_inst : DFF_X1 port map( D => n5532, CK => CLK, Q => 
                           n19188, QN => n15971);
   REGISTERS_reg_29_30_inst : DFF_X1 port map( D => n5531, CK => CLK, Q => 
                           n19208, QN => n15972);
   REGISTERS_reg_29_29_inst : DFF_X1 port map( D => n5530, CK => CLK, Q => 
                           n19228, QN => n15973);
   REGISTERS_reg_29_28_inst : DFF_X1 port map( D => n5529, CK => CLK, Q => 
                           n19248, QN => n15974);
   REGISTERS_reg_29_27_inst : DFF_X1 port map( D => n5528, CK => CLK, Q => 
                           n19268, QN => n15975);
   REGISTERS_reg_29_26_inst : DFF_X1 port map( D => n5527, CK => CLK, Q => 
                           n19288, QN => n15976);
   REGISTERS_reg_29_25_inst : DFF_X1 port map( D => n5526, CK => CLK, Q => 
                           n19308, QN => n15977);
   REGISTERS_reg_29_24_inst : DFF_X1 port map( D => n5525, CK => CLK, Q => 
                           n19328, QN => n15978);
   REGISTERS_reg_29_23_inst : DFF_X1 port map( D => n5524, CK => CLK, Q => 
                           n19348, QN => n15979);
   REGISTERS_reg_29_22_inst : DFF_X1 port map( D => n5523, CK => CLK, Q => 
                           n19368, QN => n15980);
   REGISTERS_reg_29_21_inst : DFF_X1 port map( D => n5522, CK => CLK, Q => 
                           n19388, QN => n15981);
   REGISTERS_reg_29_20_inst : DFF_X1 port map( D => n5521, CK => CLK, Q => 
                           n19408, QN => n15982);
   REGISTERS_reg_29_19_inst : DFF_X1 port map( D => n5520, CK => CLK, Q => 
                           n19428, QN => n15983);
   REGISTERS_reg_29_18_inst : DFF_X1 port map( D => n5519, CK => CLK, Q => 
                           n19448, QN => n15984);
   REGISTERS_reg_29_17_inst : DFF_X1 port map( D => n5518, CK => CLK, Q => 
                           n19468, QN => n15985);
   REGISTERS_reg_29_16_inst : DFF_X1 port map( D => n5517, CK => CLK, Q => 
                           n19488, QN => n15986);
   REGISTERS_reg_29_15_inst : DFF_X1 port map( D => n5516, CK => CLK, Q => 
                           n19508, QN => n15987);
   REGISTERS_reg_29_14_inst : DFF_X1 port map( D => n5515, CK => CLK, Q => 
                           n19528, QN => n15988);
   REGISTERS_reg_29_13_inst : DFF_X1 port map( D => n5514, CK => CLK, Q => 
                           n19548, QN => n15989);
   REGISTERS_reg_29_12_inst : DFF_X1 port map( D => n5513, CK => CLK, Q => 
                           n19568, QN => n15990);
   REGISTERS_reg_29_11_inst : DFF_X1 port map( D => n5512, CK => CLK, Q => 
                           n19588, QN => n15991);
   REGISTERS_reg_29_10_inst : DFF_X1 port map( D => n5511, CK => CLK, Q => 
                           n19608, QN => n15992);
   REGISTERS_reg_29_9_inst : DFF_X1 port map( D => n5510, CK => CLK, Q => 
                           n19628, QN => n15993);
   REGISTERS_reg_29_8_inst : DFF_X1 port map( D => n5509, CK => CLK, Q => 
                           n19648, QN => n15994);
   REGISTERS_reg_29_7_inst : DFF_X1 port map( D => n5508, CK => CLK, Q => 
                           n19668, QN => n15995);
   REGISTERS_reg_29_6_inst : DFF_X1 port map( D => n5507, CK => CLK, Q => 
                           n19688, QN => n15996);
   REGISTERS_reg_29_5_inst : DFF_X1 port map( D => n5506, CK => CLK, Q => 
                           n19708, QN => n15997);
   REGISTERS_reg_29_4_inst : DFF_X1 port map( D => n5505, CK => CLK, Q => 
                           n19728, QN => n15998);
   REGISTERS_reg_29_3_inst : DFF_X1 port map( D => n5504, CK => CLK, Q => 
                           n19748, QN => n15999);
   REGISTERS_reg_29_2_inst : DFF_X1 port map( D => n5503, CK => CLK, Q => 
                           n19768, QN => n16000);
   REGISTERS_reg_29_1_inst : DFF_X1 port map( D => n5502, CK => CLK, Q => 
                           n19788, QN => n16001);
   REGISTERS_reg_29_0_inst : DFF_X1 port map( D => n5501, CK => CLK, Q => 
                           n19808, QN => n16002);
   REGISTERS_reg_28_59_inst : DFF_X1 port map( D => n5624, CK => CLK, Q => 
                           n20121, QN => n15877);
   REGISTERS_reg_28_58_inst : DFF_X1 port map( D => n5623, CK => CLK, Q => 
                           n20120, QN => n15878);
   REGISTERS_reg_28_57_inst : DFF_X1 port map( D => n5622, CK => CLK, Q => 
                           n20119, QN => n15879);
   REGISTERS_reg_28_56_inst : DFF_X1 port map( D => n5621, CK => CLK, Q => 
                           n20118, QN => n15880);
   REGISTERS_reg_28_55_inst : DFF_X1 port map( D => n5620, CK => CLK, Q => 
                           n20117, QN => n15881);
   REGISTERS_reg_28_54_inst : DFF_X1 port map( D => n5619, CK => CLK, Q => 
                           n20116, QN => n15882);
   REGISTERS_reg_28_53_inst : DFF_X1 port map( D => n5618, CK => CLK, Q => 
                           n20115, QN => n15883);
   REGISTERS_reg_28_52_inst : DFF_X1 port map( D => n5617, CK => CLK, Q => 
                           n20114, QN => n15884);
   REGISTERS_reg_28_51_inst : DFF_X1 port map( D => n5616, CK => CLK, Q => 
                           n20113, QN => n15885);
   REGISTERS_reg_28_50_inst : DFF_X1 port map( D => n5615, CK => CLK, Q => 
                           n20112, QN => n15886);
   REGISTERS_reg_28_49_inst : DFF_X1 port map( D => n5614, CK => CLK, Q => 
                           n20111, QN => n15887);
   REGISTERS_reg_28_48_inst : DFF_X1 port map( D => n5613, CK => CLK, Q => 
                           n20110, QN => n15888);
   REGISTERS_reg_28_47_inst : DFF_X1 port map( D => n5612, CK => CLK, Q => 
                           n20109, QN => n15889);
   REGISTERS_reg_28_46_inst : DFF_X1 port map( D => n5611, CK => CLK, Q => 
                           n20108, QN => n15890);
   REGISTERS_reg_28_45_inst : DFF_X1 port map( D => n5610, CK => CLK, Q => 
                           n20107, QN => n15891);
   REGISTERS_reg_28_44_inst : DFF_X1 port map( D => n5609, CK => CLK, Q => 
                           n20106, QN => n15892);
   REGISTERS_reg_28_43_inst : DFF_X1 port map( D => n5608, CK => CLK, Q => 
                           n20105, QN => n15893);
   REGISTERS_reg_28_42_inst : DFF_X1 port map( D => n5607, CK => CLK, Q => 
                           n20104, QN => n15894);
   REGISTERS_reg_28_41_inst : DFF_X1 port map( D => n5606, CK => CLK, Q => 
                           n20103, QN => n15895);
   REGISTERS_reg_28_40_inst : DFF_X1 port map( D => n5605, CK => CLK, Q => 
                           n20102, QN => n15896);
   REGISTERS_reg_28_39_inst : DFF_X1 port map( D => n5604, CK => CLK, Q => 
                           n20101, QN => n15897);
   REGISTERS_reg_28_38_inst : DFF_X1 port map( D => n5603, CK => CLK, Q => 
                           n20100, QN => n15898);
   REGISTERS_reg_28_37_inst : DFF_X1 port map( D => n5602, CK => CLK, Q => 
                           n20099, QN => n15899);
   REGISTERS_reg_28_36_inst : DFF_X1 port map( D => n5601, CK => CLK, Q => 
                           n20098, QN => n15900);
   REGISTERS_reg_28_35_inst : DFF_X1 port map( D => n5600, CK => CLK, Q => 
                           n20097, QN => n15901);
   REGISTERS_reg_28_34_inst : DFF_X1 port map( D => n5599, CK => CLK, Q => 
                           n20096, QN => n15902);
   REGISTERS_reg_28_33_inst : DFF_X1 port map( D => n5598, CK => CLK, Q => 
                           n20095, QN => n15903);
   REGISTERS_reg_28_32_inst : DFF_X1 port map( D => n5597, CK => CLK, Q => 
                           n20094, QN => n15904);
   REGISTERS_reg_28_31_inst : DFF_X1 port map( D => n5596, CK => CLK, Q => 
                           n20093, QN => n15905);
   REGISTERS_reg_28_30_inst : DFF_X1 port map( D => n5595, CK => CLK, Q => 
                           n20092, QN => n15906);
   REGISTERS_reg_28_29_inst : DFF_X1 port map( D => n5594, CK => CLK, Q => 
                           n20091, QN => n15907);
   REGISTERS_reg_28_28_inst : DFF_X1 port map( D => n5593, CK => CLK, Q => 
                           n20090, QN => n15908);
   REGISTERS_reg_28_27_inst : DFF_X1 port map( D => n5592, CK => CLK, Q => 
                           n20089, QN => n15909);
   REGISTERS_reg_28_26_inst : DFF_X1 port map( D => n5591, CK => CLK, Q => 
                           n20088, QN => n15910);
   REGISTERS_reg_28_25_inst : DFF_X1 port map( D => n5590, CK => CLK, Q => 
                           n20087, QN => n15911);
   REGISTERS_reg_28_24_inst : DFF_X1 port map( D => n5589, CK => CLK, Q => 
                           n20086, QN => n15912);
   REGISTERS_reg_28_23_inst : DFF_X1 port map( D => n5588, CK => CLK, Q => 
                           n20085, QN => n15913);
   REGISTERS_reg_28_22_inst : DFF_X1 port map( D => n5587, CK => CLK, Q => 
                           n20084, QN => n15914);
   REGISTERS_reg_28_21_inst : DFF_X1 port map( D => n5586, CK => CLK, Q => 
                           n20083, QN => n15915);
   REGISTERS_reg_28_20_inst : DFF_X1 port map( D => n5585, CK => CLK, Q => 
                           n20082, QN => n15916);
   REGISTERS_reg_28_19_inst : DFF_X1 port map( D => n5584, CK => CLK, Q => 
                           n20081, QN => n15917);
   REGISTERS_reg_28_18_inst : DFF_X1 port map( D => n5583, CK => CLK, Q => 
                           n20080, QN => n15918);
   REGISTERS_reg_28_17_inst : DFF_X1 port map( D => n5582, CK => CLK, Q => 
                           n20079, QN => n15919);
   REGISTERS_reg_28_16_inst : DFF_X1 port map( D => n5581, CK => CLK, Q => 
                           n20078, QN => n15920);
   REGISTERS_reg_28_15_inst : DFF_X1 port map( D => n5580, CK => CLK, Q => 
                           n20077, QN => n15921);
   REGISTERS_reg_28_14_inst : DFF_X1 port map( D => n5579, CK => CLK, Q => 
                           n20076, QN => n15922);
   REGISTERS_reg_28_13_inst : DFF_X1 port map( D => n5578, CK => CLK, Q => 
                           n20075, QN => n15923);
   REGISTERS_reg_28_12_inst : DFF_X1 port map( D => n5577, CK => CLK, Q => 
                           n20074, QN => n15924);
   REGISTERS_reg_28_11_inst : DFF_X1 port map( D => n5576, CK => CLK, Q => 
                           n20073, QN => n15925);
   REGISTERS_reg_28_10_inst : DFF_X1 port map( D => n5575, CK => CLK, Q => 
                           n20072, QN => n15926);
   REGISTERS_reg_28_9_inst : DFF_X1 port map( D => n5574, CK => CLK, Q => 
                           n20071, QN => n15927);
   REGISTERS_reg_28_8_inst : DFF_X1 port map( D => n5573, CK => CLK, Q => 
                           n20070, QN => n15928);
   REGISTERS_reg_28_7_inst : DFF_X1 port map( D => n5572, CK => CLK, Q => 
                           n20069, QN => n15929);
   REGISTERS_reg_28_6_inst : DFF_X1 port map( D => n5571, CK => CLK, Q => 
                           n20068, QN => n15930);
   REGISTERS_reg_28_5_inst : DFF_X1 port map( D => n5570, CK => CLK, Q => 
                           n20067, QN => n15931);
   REGISTERS_reg_28_4_inst : DFF_X1 port map( D => n5569, CK => CLK, Q => 
                           n20066, QN => n15932);
   REGISTERS_reg_28_3_inst : DFF_X1 port map( D => n5568, CK => CLK, Q => 
                           n20065, QN => n15933);
   REGISTERS_reg_28_2_inst : DFF_X1 port map( D => n5567, CK => CLK, Q => 
                           n20064, QN => n15934);
   REGISTERS_reg_28_1_inst : DFF_X1 port map( D => n5566, CK => CLK, Q => 
                           n20063, QN => n15935);
   REGISTERS_reg_28_0_inst : DFF_X1 port map( D => n5565, CK => CLK, Q => 
                           n20062, QN => n15936);
   REGISTERS_reg_27_59_inst : DFF_X1 port map( D => n5688, CK => CLK, Q => 
                           n18630, QN => n15811);
   REGISTERS_reg_27_58_inst : DFF_X1 port map( D => n5687, CK => CLK, Q => 
                           n18650, QN => n15812);
   REGISTERS_reg_27_57_inst : DFF_X1 port map( D => n5686, CK => CLK, Q => 
                           n18670, QN => n15813);
   REGISTERS_reg_27_56_inst : DFF_X1 port map( D => n5685, CK => CLK, Q => 
                           n18690, QN => n15814);
   REGISTERS_reg_27_55_inst : DFF_X1 port map( D => n5684, CK => CLK, Q => 
                           n18710, QN => n15815);
   REGISTERS_reg_27_54_inst : DFF_X1 port map( D => n5683, CK => CLK, Q => 
                           n18730, QN => n15816);
   REGISTERS_reg_27_53_inst : DFF_X1 port map( D => n5682, CK => CLK, Q => 
                           n18750, QN => n15817);
   REGISTERS_reg_27_52_inst : DFF_X1 port map( D => n5681, CK => CLK, Q => 
                           n18770, QN => n15818);
   REGISTERS_reg_27_51_inst : DFF_X1 port map( D => n5680, CK => CLK, Q => 
                           n18790, QN => n15819);
   REGISTERS_reg_27_50_inst : DFF_X1 port map( D => n5679, CK => CLK, Q => 
                           n18810, QN => n15820);
   REGISTERS_reg_27_49_inst : DFF_X1 port map( D => n5678, CK => CLK, Q => 
                           n18830, QN => n15821);
   REGISTERS_reg_27_48_inst : DFF_X1 port map( D => n5677, CK => CLK, Q => 
                           n18850, QN => n15822);
   REGISTERS_reg_27_47_inst : DFF_X1 port map( D => n5676, CK => CLK, Q => 
                           n18870, QN => n15823);
   REGISTERS_reg_27_46_inst : DFF_X1 port map( D => n5675, CK => CLK, Q => 
                           n18890, QN => n15824);
   REGISTERS_reg_27_45_inst : DFF_X1 port map( D => n5674, CK => CLK, Q => 
                           n18910, QN => n15825);
   REGISTERS_reg_27_44_inst : DFF_X1 port map( D => n5673, CK => CLK, Q => 
                           n18930, QN => n15826);
   REGISTERS_reg_27_43_inst : DFF_X1 port map( D => n5672, CK => CLK, Q => 
                           n18950, QN => n15827);
   REGISTERS_reg_27_42_inst : DFF_X1 port map( D => n5671, CK => CLK, Q => 
                           n18970, QN => n15828);
   REGISTERS_reg_27_41_inst : DFF_X1 port map( D => n5670, CK => CLK, Q => 
                           n18990, QN => n15829);
   REGISTERS_reg_27_40_inst : DFF_X1 port map( D => n5669, CK => CLK, Q => 
                           n19010, QN => n15830);
   REGISTERS_reg_27_39_inst : DFF_X1 port map( D => n5668, CK => CLK, Q => 
                           n19030, QN => n15831);
   REGISTERS_reg_27_38_inst : DFF_X1 port map( D => n5667, CK => CLK, Q => 
                           n19050, QN => n15832);
   REGISTERS_reg_27_37_inst : DFF_X1 port map( D => n5666, CK => CLK, Q => 
                           n19070, QN => n15833);
   REGISTERS_reg_27_36_inst : DFF_X1 port map( D => n5665, CK => CLK, Q => 
                           n19090, QN => n15834);
   REGISTERS_reg_27_35_inst : DFF_X1 port map( D => n5664, CK => CLK, Q => 
                           n19110, QN => n15835);
   REGISTERS_reg_27_34_inst : DFF_X1 port map( D => n5663, CK => CLK, Q => 
                           n19130, QN => n15836);
   REGISTERS_reg_27_33_inst : DFF_X1 port map( D => n5662, CK => CLK, Q => 
                           n19150, QN => n15837);
   REGISTERS_reg_27_32_inst : DFF_X1 port map( D => n5661, CK => CLK, Q => 
                           n19170, QN => n15838);
   REGISTERS_reg_27_31_inst : DFF_X1 port map( D => n5660, CK => CLK, Q => 
                           n19190, QN => n15839);
   REGISTERS_reg_27_30_inst : DFF_X1 port map( D => n5659, CK => CLK, Q => 
                           n19210, QN => n15840);
   REGISTERS_reg_27_29_inst : DFF_X1 port map( D => n5658, CK => CLK, Q => 
                           n19230, QN => n15841);
   REGISTERS_reg_27_28_inst : DFF_X1 port map( D => n5657, CK => CLK, Q => 
                           n19250, QN => n15842);
   REGISTERS_reg_27_27_inst : DFF_X1 port map( D => n5656, CK => CLK, Q => 
                           n19270, QN => n15843);
   REGISTERS_reg_27_26_inst : DFF_X1 port map( D => n5655, CK => CLK, Q => 
                           n19290, QN => n15844);
   REGISTERS_reg_27_25_inst : DFF_X1 port map( D => n5654, CK => CLK, Q => 
                           n19310, QN => n15845);
   REGISTERS_reg_27_24_inst : DFF_X1 port map( D => n5653, CK => CLK, Q => 
                           n19330, QN => n15846);
   REGISTERS_reg_27_23_inst : DFF_X1 port map( D => n5652, CK => CLK, Q => 
                           n19350, QN => n15847);
   REGISTERS_reg_27_22_inst : DFF_X1 port map( D => n5651, CK => CLK, Q => 
                           n19370, QN => n15848);
   REGISTERS_reg_27_21_inst : DFF_X1 port map( D => n5650, CK => CLK, Q => 
                           n19390, QN => n15849);
   REGISTERS_reg_27_20_inst : DFF_X1 port map( D => n5649, CK => CLK, Q => 
                           n19410, QN => n15850);
   REGISTERS_reg_27_19_inst : DFF_X1 port map( D => n5648, CK => CLK, Q => 
                           n19430, QN => n15851);
   REGISTERS_reg_27_18_inst : DFF_X1 port map( D => n5647, CK => CLK, Q => 
                           n19450, QN => n15852);
   REGISTERS_reg_27_17_inst : DFF_X1 port map( D => n5646, CK => CLK, Q => 
                           n19470, QN => n15853);
   REGISTERS_reg_27_16_inst : DFF_X1 port map( D => n5645, CK => CLK, Q => 
                           n19490, QN => n15854);
   REGISTERS_reg_27_15_inst : DFF_X1 port map( D => n5644, CK => CLK, Q => 
                           n19510, QN => n15855);
   REGISTERS_reg_27_14_inst : DFF_X1 port map( D => n5643, CK => CLK, Q => 
                           n19530, QN => n15856);
   REGISTERS_reg_27_13_inst : DFF_X1 port map( D => n5642, CK => CLK, Q => 
                           n19550, QN => n15857);
   REGISTERS_reg_27_12_inst : DFF_X1 port map( D => n5641, CK => CLK, Q => 
                           n19570, QN => n15858);
   REGISTERS_reg_27_11_inst : DFF_X1 port map( D => n5640, CK => CLK, Q => 
                           n19590, QN => n15859);
   REGISTERS_reg_27_10_inst : DFF_X1 port map( D => n5639, CK => CLK, Q => 
                           n19610, QN => n15860);
   REGISTERS_reg_27_9_inst : DFF_X1 port map( D => n5638, CK => CLK, Q => 
                           n19630, QN => n15861);
   REGISTERS_reg_27_8_inst : DFF_X1 port map( D => n5637, CK => CLK, Q => 
                           n19650, QN => n15862);
   REGISTERS_reg_27_7_inst : DFF_X1 port map( D => n5636, CK => CLK, Q => 
                           n19670, QN => n15863);
   REGISTERS_reg_27_6_inst : DFF_X1 port map( D => n5635, CK => CLK, Q => 
                           n19690, QN => n15864);
   REGISTERS_reg_27_5_inst : DFF_X1 port map( D => n5634, CK => CLK, Q => 
                           n19710, QN => n15865);
   REGISTERS_reg_27_4_inst : DFF_X1 port map( D => n5633, CK => CLK, Q => 
                           n19730, QN => n15866);
   REGISTERS_reg_27_3_inst : DFF_X1 port map( D => n5632, CK => CLK, Q => 
                           n19750, QN => n15867);
   REGISTERS_reg_27_2_inst : DFF_X1 port map( D => n5631, CK => CLK, Q => 
                           n19770, QN => n15868);
   REGISTERS_reg_27_1_inst : DFF_X1 port map( D => n5630, CK => CLK, Q => 
                           n19790, QN => n15869);
   REGISTERS_reg_27_0_inst : DFF_X1 port map( D => n5629, CK => CLK, Q => 
                           n19810, QN => n15870);
   REGISTERS_reg_26_59_inst : DFF_X1 port map( D => n5752, CK => CLK, Q => 
                           n20061, QN => n15745);
   REGISTERS_reg_26_58_inst : DFF_X1 port map( D => n5751, CK => CLK, Q => 
                           n20060, QN => n15746);
   REGISTERS_reg_26_57_inst : DFF_X1 port map( D => n5750, CK => CLK, Q => 
                           n20059, QN => n15747);
   REGISTERS_reg_26_56_inst : DFF_X1 port map( D => n5749, CK => CLK, Q => 
                           n20058, QN => n15748);
   REGISTERS_reg_26_55_inst : DFF_X1 port map( D => n5748, CK => CLK, Q => 
                           n20057, QN => n15749);
   REGISTERS_reg_26_54_inst : DFF_X1 port map( D => n5747, CK => CLK, Q => 
                           n20056, QN => n15750);
   REGISTERS_reg_26_53_inst : DFF_X1 port map( D => n5746, CK => CLK, Q => 
                           n20055, QN => n15751);
   REGISTERS_reg_26_52_inst : DFF_X1 port map( D => n5745, CK => CLK, Q => 
                           n20054, QN => n15752);
   REGISTERS_reg_26_51_inst : DFF_X1 port map( D => n5744, CK => CLK, Q => 
                           n20053, QN => n15753);
   REGISTERS_reg_26_50_inst : DFF_X1 port map( D => n5743, CK => CLK, Q => 
                           n20052, QN => n15754);
   REGISTERS_reg_26_49_inst : DFF_X1 port map( D => n5742, CK => CLK, Q => 
                           n20051, QN => n15755);
   REGISTERS_reg_26_48_inst : DFF_X1 port map( D => n5741, CK => CLK, Q => 
                           n20050, QN => n15756);
   REGISTERS_reg_26_47_inst : DFF_X1 port map( D => n5740, CK => CLK, Q => 
                           n20049, QN => n15757);
   REGISTERS_reg_26_46_inst : DFF_X1 port map( D => n5739, CK => CLK, Q => 
                           n20048, QN => n15758);
   REGISTERS_reg_26_45_inst : DFF_X1 port map( D => n5738, CK => CLK, Q => 
                           n20047, QN => n15759);
   REGISTERS_reg_26_44_inst : DFF_X1 port map( D => n5737, CK => CLK, Q => 
                           n20046, QN => n15760);
   REGISTERS_reg_26_43_inst : DFF_X1 port map( D => n5736, CK => CLK, Q => 
                           n20045, QN => n15761);
   REGISTERS_reg_26_42_inst : DFF_X1 port map( D => n5735, CK => CLK, Q => 
                           n20044, QN => n15762);
   REGISTERS_reg_26_41_inst : DFF_X1 port map( D => n5734, CK => CLK, Q => 
                           n20043, QN => n15763);
   REGISTERS_reg_26_40_inst : DFF_X1 port map( D => n5733, CK => CLK, Q => 
                           n20042, QN => n15764);
   REGISTERS_reg_26_39_inst : DFF_X1 port map( D => n5732, CK => CLK, Q => 
                           n20041, QN => n15765);
   REGISTERS_reg_26_38_inst : DFF_X1 port map( D => n5731, CK => CLK, Q => 
                           n20040, QN => n15766);
   REGISTERS_reg_26_37_inst : DFF_X1 port map( D => n5730, CK => CLK, Q => 
                           n20039, QN => n15767);
   REGISTERS_reg_26_36_inst : DFF_X1 port map( D => n5729, CK => CLK, Q => 
                           n20038, QN => n15768);
   REGISTERS_reg_26_35_inst : DFF_X1 port map( D => n5728, CK => CLK, Q => 
                           n20037, QN => n15769);
   REGISTERS_reg_26_34_inst : DFF_X1 port map( D => n5727, CK => CLK, Q => 
                           n20036, QN => n15770);
   REGISTERS_reg_26_33_inst : DFF_X1 port map( D => n5726, CK => CLK, Q => 
                           n20035, QN => n15771);
   REGISTERS_reg_26_32_inst : DFF_X1 port map( D => n5725, CK => CLK, Q => 
                           n20034, QN => n15772);
   REGISTERS_reg_26_31_inst : DFF_X1 port map( D => n5724, CK => CLK, Q => 
                           n20033, QN => n15773);
   REGISTERS_reg_26_30_inst : DFF_X1 port map( D => n5723, CK => CLK, Q => 
                           n20032, QN => n15774);
   REGISTERS_reg_26_29_inst : DFF_X1 port map( D => n5722, CK => CLK, Q => 
                           n20031, QN => n15775);
   REGISTERS_reg_26_28_inst : DFF_X1 port map( D => n5721, CK => CLK, Q => 
                           n20030, QN => n15776);
   REGISTERS_reg_26_27_inst : DFF_X1 port map( D => n5720, CK => CLK, Q => 
                           n20029, QN => n15777);
   REGISTERS_reg_26_26_inst : DFF_X1 port map( D => n5719, CK => CLK, Q => 
                           n20028, QN => n15778);
   REGISTERS_reg_26_25_inst : DFF_X1 port map( D => n5718, CK => CLK, Q => 
                           n20027, QN => n15779);
   REGISTERS_reg_26_24_inst : DFF_X1 port map( D => n5717, CK => CLK, Q => 
                           n20026, QN => n15780);
   REGISTERS_reg_26_23_inst : DFF_X1 port map( D => n5716, CK => CLK, Q => 
                           n20025, QN => n15781);
   REGISTERS_reg_26_22_inst : DFF_X1 port map( D => n5715, CK => CLK, Q => 
                           n20024, QN => n15782);
   REGISTERS_reg_26_21_inst : DFF_X1 port map( D => n5714, CK => CLK, Q => 
                           n20023, QN => n15783);
   REGISTERS_reg_26_20_inst : DFF_X1 port map( D => n5713, CK => CLK, Q => 
                           n20022, QN => n15784);
   REGISTERS_reg_26_19_inst : DFF_X1 port map( D => n5712, CK => CLK, Q => 
                           n20021, QN => n15785);
   REGISTERS_reg_26_18_inst : DFF_X1 port map( D => n5711, CK => CLK, Q => 
                           n20020, QN => n15786);
   REGISTERS_reg_26_17_inst : DFF_X1 port map( D => n5710, CK => CLK, Q => 
                           n20019, QN => n15787);
   REGISTERS_reg_26_16_inst : DFF_X1 port map( D => n5709, CK => CLK, Q => 
                           n20018, QN => n15788);
   REGISTERS_reg_26_15_inst : DFF_X1 port map( D => n5708, CK => CLK, Q => 
                           n20017, QN => n15789);
   REGISTERS_reg_26_14_inst : DFF_X1 port map( D => n5707, CK => CLK, Q => 
                           n20016, QN => n15790);
   REGISTERS_reg_26_13_inst : DFF_X1 port map( D => n5706, CK => CLK, Q => 
                           n20015, QN => n15791);
   REGISTERS_reg_26_12_inst : DFF_X1 port map( D => n5705, CK => CLK, Q => 
                           n20014, QN => n15792);
   REGISTERS_reg_26_11_inst : DFF_X1 port map( D => n5704, CK => CLK, Q => 
                           n20013, QN => n15793);
   REGISTERS_reg_26_10_inst : DFF_X1 port map( D => n5703, CK => CLK, Q => 
                           n20012, QN => n15794);
   REGISTERS_reg_26_9_inst : DFF_X1 port map( D => n5702, CK => CLK, Q => 
                           n20011, QN => n15795);
   REGISTERS_reg_26_8_inst : DFF_X1 port map( D => n5701, CK => CLK, Q => 
                           n20010, QN => n15796);
   REGISTERS_reg_26_7_inst : DFF_X1 port map( D => n5700, CK => CLK, Q => 
                           n20009, QN => n15797);
   REGISTERS_reg_26_6_inst : DFF_X1 port map( D => n5699, CK => CLK, Q => 
                           n20008, QN => n15798);
   REGISTERS_reg_26_5_inst : DFF_X1 port map( D => n5698, CK => CLK, Q => 
                           n20007, QN => n15799);
   REGISTERS_reg_26_4_inst : DFF_X1 port map( D => n5697, CK => CLK, Q => 
                           n20006, QN => n15800);
   REGISTERS_reg_26_3_inst : DFF_X1 port map( D => n5696, CK => CLK, Q => 
                           n20005, QN => n15801);
   REGISTERS_reg_26_2_inst : DFF_X1 port map( D => n5695, CK => CLK, Q => 
                           n20004, QN => n15802);
   REGISTERS_reg_26_1_inst : DFF_X1 port map( D => n5694, CK => CLK, Q => 
                           n20003, QN => n15803);
   REGISTERS_reg_26_0_inst : DFF_X1 port map( D => n5693, CK => CLK, Q => 
                           n20002, QN => n15804);
   REGISTERS_reg_25_59_inst : DFF_X1 port map( D => n5816, CK => CLK, Q => 
                           n8973, QN => n15676);
   REGISTERS_reg_25_58_inst : DFF_X1 port map( D => n5815, CK => CLK, Q => 
                           n8977, QN => n15677);
   REGISTERS_reg_25_57_inst : DFF_X1 port map( D => n5814, CK => CLK, Q => 
                           n8981, QN => n15678);
   REGISTERS_reg_25_56_inst : DFF_X1 port map( D => n5813, CK => CLK, Q => 
                           n8985, QN => n15679);
   REGISTERS_reg_25_55_inst : DFF_X1 port map( D => n5812, CK => CLK, Q => 
                           n8989, QN => n15680);
   REGISTERS_reg_25_54_inst : DFF_X1 port map( D => n5811, CK => CLK, Q => 
                           n8993, QN => n15681);
   REGISTERS_reg_25_53_inst : DFF_X1 port map( D => n5810, CK => CLK, Q => 
                           n8997, QN => n15682);
   REGISTERS_reg_25_52_inst : DFF_X1 port map( D => n5809, CK => CLK, Q => 
                           n9001, QN => n15683);
   REGISTERS_reg_25_51_inst : DFF_X1 port map( D => n5808, CK => CLK, Q => 
                           n9005, QN => n15684);
   REGISTERS_reg_25_50_inst : DFF_X1 port map( D => n5807, CK => CLK, Q => 
                           n9009, QN => n15685);
   REGISTERS_reg_25_49_inst : DFF_X1 port map( D => n5806, CK => CLK, Q => 
                           n9013, QN => n15686);
   REGISTERS_reg_25_48_inst : DFF_X1 port map( D => n5805, CK => CLK, Q => 
                           n9017, QN => n15687);
   REGISTERS_reg_25_47_inst : DFF_X1 port map( D => n5804, CK => CLK, Q => 
                           n9021, QN => n15688);
   REGISTERS_reg_25_46_inst : DFF_X1 port map( D => n5803, CK => CLK, Q => 
                           n9025, QN => n15689);
   REGISTERS_reg_25_45_inst : DFF_X1 port map( D => n5802, CK => CLK, Q => 
                           n9029, QN => n15690);
   REGISTERS_reg_25_44_inst : DFF_X1 port map( D => n5801, CK => CLK, Q => 
                           n9033, QN => n15691);
   REGISTERS_reg_25_43_inst : DFF_X1 port map( D => n5800, CK => CLK, Q => 
                           n9037, QN => n15692);
   REGISTERS_reg_25_42_inst : DFF_X1 port map( D => n5799, CK => CLK, Q => 
                           n9041, QN => n15693);
   REGISTERS_reg_25_41_inst : DFF_X1 port map( D => n5798, CK => CLK, Q => 
                           n9045, QN => n15694);
   REGISTERS_reg_25_40_inst : DFF_X1 port map( D => n5797, CK => CLK, Q => 
                           n9049, QN => n15695);
   REGISTERS_reg_25_39_inst : DFF_X1 port map( D => n5796, CK => CLK, Q => 
                           n9053, QN => n15696);
   REGISTERS_reg_25_38_inst : DFF_X1 port map( D => n5795, CK => CLK, Q => 
                           n9057, QN => n15697);
   REGISTERS_reg_25_37_inst : DFF_X1 port map( D => n5794, CK => CLK, Q => 
                           n9061, QN => n15698);
   REGISTERS_reg_25_36_inst : DFF_X1 port map( D => n5793, CK => CLK, Q => 
                           n9065, QN => n15699);
   REGISTERS_reg_25_35_inst : DFF_X1 port map( D => n5792, CK => CLK, Q => 
                           n9069, QN => n15700);
   REGISTERS_reg_25_34_inst : DFF_X1 port map( D => n5791, CK => CLK, Q => 
                           n9073, QN => n15701);
   REGISTERS_reg_25_33_inst : DFF_X1 port map( D => n5790, CK => CLK, Q => 
                           n9077, QN => n15702);
   REGISTERS_reg_25_32_inst : DFF_X1 port map( D => n5789, CK => CLK, Q => 
                           n9081, QN => n15703);
   REGISTERS_reg_25_31_inst : DFF_X1 port map( D => n5788, CK => CLK, Q => 
                           n9085, QN => n15704);
   REGISTERS_reg_25_30_inst : DFF_X1 port map( D => n5787, CK => CLK, Q => 
                           n9089, QN => n15705);
   REGISTERS_reg_25_29_inst : DFF_X1 port map( D => n5786, CK => CLK, Q => 
                           n9093, QN => n15706);
   REGISTERS_reg_25_28_inst : DFF_X1 port map( D => n5785, CK => CLK, Q => 
                           n9097, QN => n15707);
   REGISTERS_reg_25_27_inst : DFF_X1 port map( D => n5784, CK => CLK, Q => 
                           n9101, QN => n15708);
   REGISTERS_reg_25_26_inst : DFF_X1 port map( D => n5783, CK => CLK, Q => 
                           n9105, QN => n15709);
   REGISTERS_reg_25_25_inst : DFF_X1 port map( D => n5782, CK => CLK, Q => 
                           n9109, QN => n15710);
   REGISTERS_reg_25_24_inst : DFF_X1 port map( D => n5781, CK => CLK, Q => 
                           n9113, QN => n15711);
   REGISTERS_reg_25_23_inst : DFF_X1 port map( D => n5780, CK => CLK, Q => 
                           n9117, QN => n15712);
   REGISTERS_reg_25_22_inst : DFF_X1 port map( D => n5779, CK => CLK, Q => 
                           n9121, QN => n15713);
   REGISTERS_reg_25_21_inst : DFF_X1 port map( D => n5778, CK => CLK, Q => 
                           n9125, QN => n15714);
   REGISTERS_reg_25_20_inst : DFF_X1 port map( D => n5777, CK => CLK, Q => 
                           n9129, QN => n15715);
   REGISTERS_reg_25_19_inst : DFF_X1 port map( D => n5776, CK => CLK, Q => 
                           n9133, QN => n15716);
   REGISTERS_reg_25_18_inst : DFF_X1 port map( D => n5775, CK => CLK, Q => 
                           n9137, QN => n15717);
   REGISTERS_reg_25_17_inst : DFF_X1 port map( D => n5774, CK => CLK, Q => 
                           n9141, QN => n15718);
   REGISTERS_reg_25_16_inst : DFF_X1 port map( D => n5773, CK => CLK, Q => 
                           n9145, QN => n15719);
   REGISTERS_reg_25_15_inst : DFF_X1 port map( D => n5772, CK => CLK, Q => 
                           n9149, QN => n15720);
   REGISTERS_reg_25_14_inst : DFF_X1 port map( D => n5771, CK => CLK, Q => 
                           n9153, QN => n15721);
   REGISTERS_reg_25_13_inst : DFF_X1 port map( D => n5770, CK => CLK, Q => 
                           n9157, QN => n15722);
   REGISTERS_reg_25_12_inst : DFF_X1 port map( D => n5769, CK => CLK, Q => 
                           n9161, QN => n15723);
   REGISTERS_reg_25_11_inst : DFF_X1 port map( D => n5768, CK => CLK, Q => 
                           n9165, QN => n15724);
   REGISTERS_reg_25_10_inst : DFF_X1 port map( D => n5767, CK => CLK, Q => 
                           n9169, QN => n15725);
   REGISTERS_reg_25_9_inst : DFF_X1 port map( D => n5766, CK => CLK, Q => n9173
                           , QN => n15726);
   REGISTERS_reg_25_8_inst : DFF_X1 port map( D => n5765, CK => CLK, Q => n9177
                           , QN => n15727);
   REGISTERS_reg_25_7_inst : DFF_X1 port map( D => n5764, CK => CLK, Q => n9181
                           , QN => n15728);
   REGISTERS_reg_25_6_inst : DFF_X1 port map( D => n5763, CK => CLK, Q => n9185
                           , QN => n15729);
   REGISTERS_reg_25_5_inst : DFF_X1 port map( D => n5762, CK => CLK, Q => n9189
                           , QN => n15730);
   REGISTERS_reg_25_4_inst : DFF_X1 port map( D => n5761, CK => CLK, Q => n9193
                           , QN => n15731);
   REGISTERS_reg_25_3_inst : DFF_X1 port map( D => n5760, CK => CLK, Q => n9197
                           , QN => n15732);
   REGISTERS_reg_25_2_inst : DFF_X1 port map( D => n5759, CK => CLK, Q => n9201
                           , QN => n15733);
   REGISTERS_reg_25_1_inst : DFF_X1 port map( D => n5758, CK => CLK, Q => n9205
                           , QN => n15734);
   REGISTERS_reg_25_0_inst : DFF_X1 port map( D => n5757, CK => CLK, Q => n9209
                           , QN => n15735);
   REGISTERS_reg_31_59_inst : DFF_X1 port map( D => n5428, CK => CLK, Q => 
                           n18624, QN => n16181);
   REGISTERS_reg_31_58_inst : DFF_X1 port map( D => n5426, CK => CLK, Q => 
                           n18644, QN => n16200);
   REGISTERS_reg_31_57_inst : DFF_X1 port map( D => n5424, CK => CLK, Q => 
                           n18664, QN => n16219);
   REGISTERS_reg_31_56_inst : DFF_X1 port map( D => n5422, CK => CLK, Q => 
                           n18684, QN => n16238);
   REGISTERS_reg_31_55_inst : DFF_X1 port map( D => n5420, CK => CLK, Q => 
                           n18704, QN => n16257);
   REGISTERS_reg_31_54_inst : DFF_X1 port map( D => n5418, CK => CLK, Q => 
                           n18724, QN => n16276);
   REGISTERS_reg_31_53_inst : DFF_X1 port map( D => n5416, CK => CLK, Q => 
                           n18744, QN => n16295);
   REGISTERS_reg_31_52_inst : DFF_X1 port map( D => n5414, CK => CLK, Q => 
                           n18764, QN => n16314);
   REGISTERS_reg_31_51_inst : DFF_X1 port map( D => n5412, CK => CLK, Q => 
                           n18784, QN => n16333);
   REGISTERS_reg_31_50_inst : DFF_X1 port map( D => n5410, CK => CLK, Q => 
                           n18804, QN => n16352);
   REGISTERS_reg_31_49_inst : DFF_X1 port map( D => n5408, CK => CLK, Q => 
                           n18824, QN => n16371);
   REGISTERS_reg_31_48_inst : DFF_X1 port map( D => n5406, CK => CLK, Q => 
                           n18844, QN => n16390);
   REGISTERS_reg_31_47_inst : DFF_X1 port map( D => n5404, CK => CLK, Q => 
                           n18864, QN => n16409);
   REGISTERS_reg_31_46_inst : DFF_X1 port map( D => n5402, CK => CLK, Q => 
                           n18884, QN => n16428);
   REGISTERS_reg_31_45_inst : DFF_X1 port map( D => n5400, CK => CLK, Q => 
                           n18904, QN => n16447);
   REGISTERS_reg_31_44_inst : DFF_X1 port map( D => n5398, CK => CLK, Q => 
                           n18924, QN => n16466);
   REGISTERS_reg_31_43_inst : DFF_X1 port map( D => n5396, CK => CLK, Q => 
                           n18944, QN => n16485);
   REGISTERS_reg_31_42_inst : DFF_X1 port map( D => n5394, CK => CLK, Q => 
                           n18964, QN => n16504);
   REGISTERS_reg_31_41_inst : DFF_X1 port map( D => n5392, CK => CLK, Q => 
                           n18984, QN => n16523);
   REGISTERS_reg_31_40_inst : DFF_X1 port map( D => n5390, CK => CLK, Q => 
                           n19004, QN => n16542);
   REGISTERS_reg_31_39_inst : DFF_X1 port map( D => n5388, CK => CLK, Q => 
                           n19024, QN => n16561);
   REGISTERS_reg_31_38_inst : DFF_X1 port map( D => n5386, CK => CLK, Q => 
                           n19044, QN => n16580);
   REGISTERS_reg_31_37_inst : DFF_X1 port map( D => n5384, CK => CLK, Q => 
                           n19064, QN => n16599);
   REGISTERS_reg_31_36_inst : DFF_X1 port map( D => n5382, CK => CLK, Q => 
                           n19084, QN => n16618);
   REGISTERS_reg_31_35_inst : DFF_X1 port map( D => n5380, CK => CLK, Q => 
                           n19104, QN => n16637);
   REGISTERS_reg_31_34_inst : DFF_X1 port map( D => n5378, CK => CLK, Q => 
                           n19124, QN => n16656);
   REGISTERS_reg_31_33_inst : DFF_X1 port map( D => n5376, CK => CLK, Q => 
                           n19144, QN => n16675);
   REGISTERS_reg_31_32_inst : DFF_X1 port map( D => n5374, CK => CLK, Q => 
                           n19164, QN => n16694);
   REGISTERS_reg_31_31_inst : DFF_X1 port map( D => n5372, CK => CLK, Q => 
                           n19184, QN => n16713);
   REGISTERS_reg_31_30_inst : DFF_X1 port map( D => n5370, CK => CLK, Q => 
                           n19204, QN => n16732);
   REGISTERS_reg_31_29_inst : DFF_X1 port map( D => n5368, CK => CLK, Q => 
                           n19224, QN => n16751);
   REGISTERS_reg_31_28_inst : DFF_X1 port map( D => n5366, CK => CLK, Q => 
                           n19244, QN => n16770);
   REGISTERS_reg_31_27_inst : DFF_X1 port map( D => n5364, CK => CLK, Q => 
                           n19264, QN => n16789);
   REGISTERS_reg_31_26_inst : DFF_X1 port map( D => n5362, CK => CLK, Q => 
                           n19284, QN => n16808);
   REGISTERS_reg_31_25_inst : DFF_X1 port map( D => n5360, CK => CLK, Q => 
                           n19304, QN => n16827);
   REGISTERS_reg_31_24_inst : DFF_X1 port map( D => n5358, CK => CLK, Q => 
                           n19324, QN => n16846);
   REGISTERS_reg_31_23_inst : DFF_X1 port map( D => n5356, CK => CLK, Q => 
                           n19344, QN => n16865);
   REGISTERS_reg_31_22_inst : DFF_X1 port map( D => n5354, CK => CLK, Q => 
                           n19364, QN => n16884);
   REGISTERS_reg_31_21_inst : DFF_X1 port map( D => n5352, CK => CLK, Q => 
                           n19384, QN => n16903);
   REGISTERS_reg_31_20_inst : DFF_X1 port map( D => n5350, CK => CLK, Q => 
                           n19404, QN => n16922);
   REGISTERS_reg_31_19_inst : DFF_X1 port map( D => n5348, CK => CLK, Q => 
                           n19424, QN => n16941);
   REGISTERS_reg_31_18_inst : DFF_X1 port map( D => n5346, CK => CLK, Q => 
                           n19444, QN => n16960);
   REGISTERS_reg_31_17_inst : DFF_X1 port map( D => n5344, CK => CLK, Q => 
                           n19464, QN => n16979);
   REGISTERS_reg_31_16_inst : DFF_X1 port map( D => n5342, CK => CLK, Q => 
                           n19484, QN => n16998);
   REGISTERS_reg_31_15_inst : DFF_X1 port map( D => n5340, CK => CLK, Q => 
                           n19504, QN => n17017);
   REGISTERS_reg_31_14_inst : DFF_X1 port map( D => n5338, CK => CLK, Q => 
                           n19524, QN => n17036);
   REGISTERS_reg_31_13_inst : DFF_X1 port map( D => n5336, CK => CLK, Q => 
                           n19544, QN => n17055);
   REGISTERS_reg_31_12_inst : DFF_X1 port map( D => n5334, CK => CLK, Q => 
                           n19564, QN => n17074);
   REGISTERS_reg_31_11_inst : DFF_X1 port map( D => n5332, CK => CLK, Q => 
                           n19584, QN => n17093);
   REGISTERS_reg_31_10_inst : DFF_X1 port map( D => n5330, CK => CLK, Q => 
                           n19604, QN => n17112);
   REGISTERS_reg_31_9_inst : DFF_X1 port map( D => n5328, CK => CLK, Q => 
                           n19624, QN => n17131);
   REGISTERS_reg_31_8_inst : DFF_X1 port map( D => n5326, CK => CLK, Q => 
                           n19644, QN => n17150);
   REGISTERS_reg_31_7_inst : DFF_X1 port map( D => n5324, CK => CLK, Q => 
                           n19664, QN => n17169);
   REGISTERS_reg_31_6_inst : DFF_X1 port map( D => n5322, CK => CLK, Q => 
                           n19684, QN => n17188);
   REGISTERS_reg_31_5_inst : DFF_X1 port map( D => n5320, CK => CLK, Q => 
                           n19704, QN => n17207);
   REGISTERS_reg_31_4_inst : DFF_X1 port map( D => n5318, CK => CLK, Q => 
                           n19724, QN => n17226);
   REGISTERS_reg_31_3_inst : DFF_X1 port map( D => n5316, CK => CLK, Q => 
                           n19744, QN => n17245);
   REGISTERS_reg_31_2_inst : DFF_X1 port map( D => n5314, CK => CLK, Q => 
                           n19764, QN => n17264);
   REGISTERS_reg_31_1_inst : DFF_X1 port map( D => n5312, CK => CLK, Q => 
                           n19784, QN => n17283);
   REGISTERS_reg_31_0_inst : DFF_X1 port map( D => n5310, CK => CLK, Q => 
                           n19804, QN => n17302);
   REGISTERS_reg_23_59_inst : DFF_X1 port map( D => n5944, CK => CLK, Q => 
                           n8837, QN => n15543);
   REGISTERS_reg_23_58_inst : DFF_X1 port map( D => n5943, CK => CLK, Q => 
                           n8839, QN => n15544);
   REGISTERS_reg_23_57_inst : DFF_X1 port map( D => n5942, CK => CLK, Q => 
                           n8841, QN => n15545);
   REGISTERS_reg_23_56_inst : DFF_X1 port map( D => n5941, CK => CLK, Q => 
                           n8843, QN => n15546);
   REGISTERS_reg_23_55_inst : DFF_X1 port map( D => n5940, CK => CLK, Q => 
                           n8845, QN => n15547);
   REGISTERS_reg_23_54_inst : DFF_X1 port map( D => n5939, CK => CLK, Q => 
                           n8847, QN => n15548);
   REGISTERS_reg_23_53_inst : DFF_X1 port map( D => n5938, CK => CLK, Q => 
                           n8849, QN => n15549);
   REGISTERS_reg_23_52_inst : DFF_X1 port map( D => n5937, CK => CLK, Q => 
                           n8851, QN => n15550);
   REGISTERS_reg_23_51_inst : DFF_X1 port map( D => n5936, CK => CLK, Q => 
                           n8853, QN => n15551);
   REGISTERS_reg_23_50_inst : DFF_X1 port map( D => n5935, CK => CLK, Q => 
                           n8855, QN => n15552);
   REGISTERS_reg_23_49_inst : DFF_X1 port map( D => n5934, CK => CLK, Q => 
                           n8857, QN => n15553);
   REGISTERS_reg_23_48_inst : DFF_X1 port map( D => n5933, CK => CLK, Q => 
                           n8859, QN => n15554);
   REGISTERS_reg_23_47_inst : DFF_X1 port map( D => n5932, CK => CLK, Q => 
                           n8861, QN => n15555);
   REGISTERS_reg_23_46_inst : DFF_X1 port map( D => n5931, CK => CLK, Q => 
                           n8863, QN => n15556);
   REGISTERS_reg_23_45_inst : DFF_X1 port map( D => n5930, CK => CLK, Q => 
                           n8865, QN => n15557);
   REGISTERS_reg_23_44_inst : DFF_X1 port map( D => n5929, CK => CLK, Q => 
                           n8867, QN => n15558);
   REGISTERS_reg_23_43_inst : DFF_X1 port map( D => n5928, CK => CLK, Q => 
                           n8869, QN => n15559);
   REGISTERS_reg_23_42_inst : DFF_X1 port map( D => n5927, CK => CLK, Q => 
                           n8871, QN => n15560);
   REGISTERS_reg_23_41_inst : DFF_X1 port map( D => n5926, CK => CLK, Q => 
                           n8873, QN => n15561);
   REGISTERS_reg_23_40_inst : DFF_X1 port map( D => n5925, CK => CLK, Q => 
                           n8875, QN => n15562);
   REGISTERS_reg_23_39_inst : DFF_X1 port map( D => n5924, CK => CLK, Q => 
                           n8877, QN => n15563);
   REGISTERS_reg_23_38_inst : DFF_X1 port map( D => n5923, CK => CLK, Q => 
                           n8879, QN => n15564);
   REGISTERS_reg_23_37_inst : DFF_X1 port map( D => n5922, CK => CLK, Q => 
                           n8881, QN => n15565);
   REGISTERS_reg_23_36_inst : DFF_X1 port map( D => n5921, CK => CLK, Q => 
                           n8883, QN => n15566);
   REGISTERS_reg_23_35_inst : DFF_X1 port map( D => n5920, CK => CLK, Q => 
                           n8885, QN => n15567);
   REGISTERS_reg_23_34_inst : DFF_X1 port map( D => n5919, CK => CLK, Q => 
                           n8887, QN => n15568);
   REGISTERS_reg_23_33_inst : DFF_X1 port map( D => n5918, CK => CLK, Q => 
                           n8889, QN => n15569);
   REGISTERS_reg_23_32_inst : DFF_X1 port map( D => n5917, CK => CLK, Q => 
                           n8891, QN => n15570);
   REGISTERS_reg_23_31_inst : DFF_X1 port map( D => n5916, CK => CLK, Q => 
                           n8893, QN => n15571);
   REGISTERS_reg_23_30_inst : DFF_X1 port map( D => n5915, CK => CLK, Q => 
                           n8895, QN => n15572);
   REGISTERS_reg_23_29_inst : DFF_X1 port map( D => n5914, CK => CLK, Q => 
                           n8897, QN => n15573);
   REGISTERS_reg_23_28_inst : DFF_X1 port map( D => n5913, CK => CLK, Q => 
                           n8899, QN => n15574);
   REGISTERS_reg_23_27_inst : DFF_X1 port map( D => n5912, CK => CLK, Q => 
                           n8901, QN => n15575);
   REGISTERS_reg_23_26_inst : DFF_X1 port map( D => n5911, CK => CLK, Q => 
                           n8903, QN => n15576);
   REGISTERS_reg_23_25_inst : DFF_X1 port map( D => n5910, CK => CLK, Q => 
                           n8905, QN => n15577);
   REGISTERS_reg_23_24_inst : DFF_X1 port map( D => n5909, CK => CLK, Q => 
                           n8907, QN => n15578);
   REGISTERS_reg_23_23_inst : DFF_X1 port map( D => n5908, CK => CLK, Q => 
                           n8909, QN => n15579);
   REGISTERS_reg_23_22_inst : DFF_X1 port map( D => n5907, CK => CLK, Q => 
                           n8911, QN => n15580);
   REGISTERS_reg_23_21_inst : DFF_X1 port map( D => n5906, CK => CLK, Q => 
                           n8913, QN => n15581);
   REGISTERS_reg_23_20_inst : DFF_X1 port map( D => n5905, CK => CLK, Q => 
                           n8915, QN => n15582);
   REGISTERS_reg_23_19_inst : DFF_X1 port map( D => n5904, CK => CLK, Q => 
                           n8917, QN => n15583);
   REGISTERS_reg_23_18_inst : DFF_X1 port map( D => n5903, CK => CLK, Q => 
                           n8919, QN => n15584);
   REGISTERS_reg_23_17_inst : DFF_X1 port map( D => n5902, CK => CLK, Q => 
                           n8921, QN => n15585);
   REGISTERS_reg_23_16_inst : DFF_X1 port map( D => n5901, CK => CLK, Q => 
                           n8923, QN => n15586);
   REGISTERS_reg_23_15_inst : DFF_X1 port map( D => n5900, CK => CLK, Q => 
                           n8925, QN => n15587);
   REGISTERS_reg_23_14_inst : DFF_X1 port map( D => n5899, CK => CLK, Q => 
                           n8927, QN => n15588);
   REGISTERS_reg_23_13_inst : DFF_X1 port map( D => n5898, CK => CLK, Q => 
                           n8929, QN => n15589);
   REGISTERS_reg_23_12_inst : DFF_X1 port map( D => n5897, CK => CLK, Q => 
                           n8931, QN => n15590);
   REGISTERS_reg_23_11_inst : DFF_X1 port map( D => n5896, CK => CLK, Q => 
                           n8933, QN => n15591);
   REGISTERS_reg_23_10_inst : DFF_X1 port map( D => n5895, CK => CLK, Q => 
                           n8935, QN => n15592);
   REGISTERS_reg_23_9_inst : DFF_X1 port map( D => n5894, CK => CLK, Q => n8937
                           , QN => n15593);
   REGISTERS_reg_23_8_inst : DFF_X1 port map( D => n5893, CK => CLK, Q => n8939
                           , QN => n15594);
   REGISTERS_reg_23_7_inst : DFF_X1 port map( D => n5892, CK => CLK, Q => n8941
                           , QN => n15595);
   REGISTERS_reg_23_6_inst : DFF_X1 port map( D => n5891, CK => CLK, Q => n8943
                           , QN => n15596);
   REGISTERS_reg_23_5_inst : DFF_X1 port map( D => n5890, CK => CLK, Q => n8945
                           , QN => n15597);
   REGISTERS_reg_23_4_inst : DFF_X1 port map( D => n5889, CK => CLK, Q => n8947
                           , QN => n15598);
   REGISTERS_reg_23_3_inst : DFF_X1 port map( D => n5888, CK => CLK, Q => n8949
                           , QN => n15599);
   REGISTERS_reg_23_2_inst : DFF_X1 port map( D => n5887, CK => CLK, Q => n8951
                           , QN => n15600);
   REGISTERS_reg_23_1_inst : DFF_X1 port map( D => n5886, CK => CLK, Q => n8953
                           , QN => n15601);
   REGISTERS_reg_23_0_inst : DFF_X1 port map( D => n5885, CK => CLK, Q => n8955
                           , QN => n15602);
   REGISTERS_reg_22_59_inst : DFF_X1 port map( D => n6008, CK => CLK, Q => 
                           n18629, QN => n15476);
   REGISTERS_reg_22_58_inst : DFF_X1 port map( D => n6007, CK => CLK, Q => 
                           n18649, QN => n15477);
   REGISTERS_reg_22_57_inst : DFF_X1 port map( D => n6006, CK => CLK, Q => 
                           n18669, QN => n15478);
   REGISTERS_reg_22_56_inst : DFF_X1 port map( D => n6005, CK => CLK, Q => 
                           n18689, QN => n15479);
   REGISTERS_reg_22_55_inst : DFF_X1 port map( D => n6004, CK => CLK, Q => 
                           n18709, QN => n15480);
   REGISTERS_reg_22_54_inst : DFF_X1 port map( D => n6003, CK => CLK, Q => 
                           n18729, QN => n15481);
   REGISTERS_reg_22_53_inst : DFF_X1 port map( D => n6002, CK => CLK, Q => 
                           n18749, QN => n15482);
   REGISTERS_reg_22_52_inst : DFF_X1 port map( D => n6001, CK => CLK, Q => 
                           n18769, QN => n15483);
   REGISTERS_reg_22_51_inst : DFF_X1 port map( D => n6000, CK => CLK, Q => 
                           n18789, QN => n15484);
   REGISTERS_reg_22_50_inst : DFF_X1 port map( D => n5999, CK => CLK, Q => 
                           n18809, QN => n15485);
   REGISTERS_reg_22_49_inst : DFF_X1 port map( D => n5998, CK => CLK, Q => 
                           n18829, QN => n15486);
   REGISTERS_reg_22_48_inst : DFF_X1 port map( D => n5997, CK => CLK, Q => 
                           n18849, QN => n15487);
   REGISTERS_reg_22_47_inst : DFF_X1 port map( D => n5996, CK => CLK, Q => 
                           n18869, QN => n15488);
   REGISTERS_reg_22_46_inst : DFF_X1 port map( D => n5995, CK => CLK, Q => 
                           n18889, QN => n15489);
   REGISTERS_reg_22_45_inst : DFF_X1 port map( D => n5994, CK => CLK, Q => 
                           n18909, QN => n15490);
   REGISTERS_reg_22_44_inst : DFF_X1 port map( D => n5993, CK => CLK, Q => 
                           n18929, QN => n15491);
   REGISTERS_reg_22_43_inst : DFF_X1 port map( D => n5992, CK => CLK, Q => 
                           n18949, QN => n15492);
   REGISTERS_reg_22_42_inst : DFF_X1 port map( D => n5991, CK => CLK, Q => 
                           n18969, QN => n15493);
   REGISTERS_reg_22_41_inst : DFF_X1 port map( D => n5990, CK => CLK, Q => 
                           n18989, QN => n15494);
   REGISTERS_reg_22_40_inst : DFF_X1 port map( D => n5989, CK => CLK, Q => 
                           n19009, QN => n15495);
   REGISTERS_reg_22_39_inst : DFF_X1 port map( D => n5988, CK => CLK, Q => 
                           n19029, QN => n15496);
   REGISTERS_reg_22_38_inst : DFF_X1 port map( D => n5987, CK => CLK, Q => 
                           n19049, QN => n15497);
   REGISTERS_reg_22_37_inst : DFF_X1 port map( D => n5986, CK => CLK, Q => 
                           n19069, QN => n15498);
   REGISTERS_reg_22_36_inst : DFF_X1 port map( D => n5985, CK => CLK, Q => 
                           n19089, QN => n15499);
   REGISTERS_reg_22_35_inst : DFF_X1 port map( D => n5984, CK => CLK, Q => 
                           n19109, QN => n15500);
   REGISTERS_reg_22_34_inst : DFF_X1 port map( D => n5983, CK => CLK, Q => 
                           n19129, QN => n15501);
   REGISTERS_reg_22_33_inst : DFF_X1 port map( D => n5982, CK => CLK, Q => 
                           n19149, QN => n15502);
   REGISTERS_reg_22_32_inst : DFF_X1 port map( D => n5981, CK => CLK, Q => 
                           n19169, QN => n15503);
   REGISTERS_reg_22_31_inst : DFF_X1 port map( D => n5980, CK => CLK, Q => 
                           n19189, QN => n15504);
   REGISTERS_reg_22_30_inst : DFF_X1 port map( D => n5979, CK => CLK, Q => 
                           n19209, QN => n15505);
   REGISTERS_reg_22_29_inst : DFF_X1 port map( D => n5978, CK => CLK, Q => 
                           n19229, QN => n15506);
   REGISTERS_reg_22_28_inst : DFF_X1 port map( D => n5977, CK => CLK, Q => 
                           n19249, QN => n15507);
   REGISTERS_reg_22_27_inst : DFF_X1 port map( D => n5976, CK => CLK, Q => 
                           n19269, QN => n15508);
   REGISTERS_reg_22_26_inst : DFF_X1 port map( D => n5975, CK => CLK, Q => 
                           n19289, QN => n15509);
   REGISTERS_reg_22_25_inst : DFF_X1 port map( D => n5974, CK => CLK, Q => 
                           n19309, QN => n15510);
   REGISTERS_reg_22_24_inst : DFF_X1 port map( D => n5973, CK => CLK, Q => 
                           n19329, QN => n15511);
   REGISTERS_reg_22_23_inst : DFF_X1 port map( D => n5972, CK => CLK, Q => 
                           n19349, QN => n15512);
   REGISTERS_reg_22_22_inst : DFF_X1 port map( D => n5971, CK => CLK, Q => 
                           n19369, QN => n15513);
   REGISTERS_reg_22_21_inst : DFF_X1 port map( D => n5970, CK => CLK, Q => 
                           n19389, QN => n15514);
   REGISTERS_reg_22_20_inst : DFF_X1 port map( D => n5969, CK => CLK, Q => 
                           n19409, QN => n15515);
   REGISTERS_reg_22_19_inst : DFF_X1 port map( D => n5968, CK => CLK, Q => 
                           n19429, QN => n15516);
   REGISTERS_reg_22_18_inst : DFF_X1 port map( D => n5967, CK => CLK, Q => 
                           n19449, QN => n15517);
   REGISTERS_reg_22_17_inst : DFF_X1 port map( D => n5966, CK => CLK, Q => 
                           n19469, QN => n15518);
   REGISTERS_reg_22_16_inst : DFF_X1 port map( D => n5965, CK => CLK, Q => 
                           n19489, QN => n15519);
   REGISTERS_reg_22_15_inst : DFF_X1 port map( D => n5964, CK => CLK, Q => 
                           n19509, QN => n15520);
   REGISTERS_reg_22_14_inst : DFF_X1 port map( D => n5963, CK => CLK, Q => 
                           n19529, QN => n15521);
   REGISTERS_reg_22_13_inst : DFF_X1 port map( D => n5962, CK => CLK, Q => 
                           n19549, QN => n15522);
   REGISTERS_reg_22_12_inst : DFF_X1 port map( D => n5961, CK => CLK, Q => 
                           n19569, QN => n15523);
   REGISTERS_reg_22_11_inst : DFF_X1 port map( D => n5960, CK => CLK, Q => 
                           n19589, QN => n15524);
   REGISTERS_reg_22_10_inst : DFF_X1 port map( D => n5959, CK => CLK, Q => 
                           n19609, QN => n15525);
   REGISTERS_reg_22_9_inst : DFF_X1 port map( D => n5958, CK => CLK, Q => 
                           n19629, QN => n15526);
   REGISTERS_reg_22_8_inst : DFF_X1 port map( D => n5957, CK => CLK, Q => 
                           n19649, QN => n15527);
   REGISTERS_reg_22_7_inst : DFF_X1 port map( D => n5956, CK => CLK, Q => 
                           n19669, QN => n15528);
   REGISTERS_reg_22_6_inst : DFF_X1 port map( D => n5955, CK => CLK, Q => 
                           n19689, QN => n15529);
   REGISTERS_reg_22_5_inst : DFF_X1 port map( D => n5954, CK => CLK, Q => 
                           n19709, QN => n15530);
   REGISTERS_reg_22_4_inst : DFF_X1 port map( D => n5953, CK => CLK, Q => 
                           n19729, QN => n15531);
   REGISTERS_reg_22_3_inst : DFF_X1 port map( D => n5952, CK => CLK, Q => 
                           n19749, QN => n15532);
   REGISTERS_reg_22_2_inst : DFF_X1 port map( D => n5951, CK => CLK, Q => 
                           n19769, QN => n15533);
   REGISTERS_reg_22_1_inst : DFF_X1 port map( D => n5950, CK => CLK, Q => 
                           n19789, QN => n15534);
   REGISTERS_reg_22_0_inst : DFF_X1 port map( D => n5949, CK => CLK, Q => 
                           n19809, QN => n15535);
   REGISTERS_reg_21_59_inst : DFF_X1 port map( D => n6072, CK => CLK, Q => 
                           n20001, QN => n15410);
   REGISTERS_reg_21_58_inst : DFF_X1 port map( D => n6071, CK => CLK, Q => 
                           n20000, QN => n15411);
   REGISTERS_reg_21_57_inst : DFF_X1 port map( D => n6070, CK => CLK, Q => 
                           n19999, QN => n15412);
   REGISTERS_reg_21_56_inst : DFF_X1 port map( D => n6069, CK => CLK, Q => 
                           n19998, QN => n15413);
   REGISTERS_reg_21_55_inst : DFF_X1 port map( D => n6068, CK => CLK, Q => 
                           n19997, QN => n15414);
   REGISTERS_reg_21_54_inst : DFF_X1 port map( D => n6067, CK => CLK, Q => 
                           n19996, QN => n15415);
   REGISTERS_reg_21_53_inst : DFF_X1 port map( D => n6066, CK => CLK, Q => 
                           n19995, QN => n15416);
   REGISTERS_reg_21_52_inst : DFF_X1 port map( D => n6065, CK => CLK, Q => 
                           n19994, QN => n15417);
   REGISTERS_reg_21_51_inst : DFF_X1 port map( D => n6064, CK => CLK, Q => 
                           n19993, QN => n15418);
   REGISTERS_reg_21_50_inst : DFF_X1 port map( D => n6063, CK => CLK, Q => 
                           n19992, QN => n15419);
   REGISTERS_reg_21_49_inst : DFF_X1 port map( D => n6062, CK => CLK, Q => 
                           n19991, QN => n15420);
   REGISTERS_reg_21_48_inst : DFF_X1 port map( D => n6061, CK => CLK, Q => 
                           n19990, QN => n15421);
   REGISTERS_reg_21_47_inst : DFF_X1 port map( D => n6060, CK => CLK, Q => 
                           n19989, QN => n15422);
   REGISTERS_reg_21_46_inst : DFF_X1 port map( D => n6059, CK => CLK, Q => 
                           n19988, QN => n15423);
   REGISTERS_reg_21_45_inst : DFF_X1 port map( D => n6058, CK => CLK, Q => 
                           n19987, QN => n15424);
   REGISTERS_reg_21_44_inst : DFF_X1 port map( D => n6057, CK => CLK, Q => 
                           n19986, QN => n15425);
   REGISTERS_reg_21_43_inst : DFF_X1 port map( D => n6056, CK => CLK, Q => 
                           n19985, QN => n15426);
   REGISTERS_reg_21_42_inst : DFF_X1 port map( D => n6055, CK => CLK, Q => 
                           n19984, QN => n15427);
   REGISTERS_reg_21_41_inst : DFF_X1 port map( D => n6054, CK => CLK, Q => 
                           n19983, QN => n15428);
   REGISTERS_reg_21_40_inst : DFF_X1 port map( D => n6053, CK => CLK, Q => 
                           n19982, QN => n15429);
   REGISTERS_reg_21_39_inst : DFF_X1 port map( D => n6052, CK => CLK, Q => 
                           n19981, QN => n15430);
   REGISTERS_reg_21_38_inst : DFF_X1 port map( D => n6051, CK => CLK, Q => 
                           n19980, QN => n15431);
   REGISTERS_reg_21_37_inst : DFF_X1 port map( D => n6050, CK => CLK, Q => 
                           n19979, QN => n15432);
   REGISTERS_reg_21_36_inst : DFF_X1 port map( D => n6049, CK => CLK, Q => 
                           n19978, QN => n15433);
   REGISTERS_reg_21_35_inst : DFF_X1 port map( D => n6048, CK => CLK, Q => 
                           n19977, QN => n15434);
   REGISTERS_reg_21_34_inst : DFF_X1 port map( D => n6047, CK => CLK, Q => 
                           n19976, QN => n15435);
   REGISTERS_reg_21_33_inst : DFF_X1 port map( D => n6046, CK => CLK, Q => 
                           n19975, QN => n15436);
   REGISTERS_reg_21_32_inst : DFF_X1 port map( D => n6045, CK => CLK, Q => 
                           n19974, QN => n15437);
   REGISTERS_reg_21_31_inst : DFF_X1 port map( D => n6044, CK => CLK, Q => 
                           n19973, QN => n15438);
   REGISTERS_reg_21_30_inst : DFF_X1 port map( D => n6043, CK => CLK, Q => 
                           n19972, QN => n15439);
   REGISTERS_reg_21_29_inst : DFF_X1 port map( D => n6042, CK => CLK, Q => 
                           n19971, QN => n15440);
   REGISTERS_reg_21_28_inst : DFF_X1 port map( D => n6041, CK => CLK, Q => 
                           n19970, QN => n15441);
   REGISTERS_reg_21_27_inst : DFF_X1 port map( D => n6040, CK => CLK, Q => 
                           n19969, QN => n15442);
   REGISTERS_reg_21_26_inst : DFF_X1 port map( D => n6039, CK => CLK, Q => 
                           n19968, QN => n15443);
   REGISTERS_reg_21_25_inst : DFF_X1 port map( D => n6038, CK => CLK, Q => 
                           n19967, QN => n15444);
   REGISTERS_reg_21_24_inst : DFF_X1 port map( D => n6037, CK => CLK, Q => 
                           n19966, QN => n15445);
   REGISTERS_reg_21_23_inst : DFF_X1 port map( D => n6036, CK => CLK, Q => 
                           n19965, QN => n15446);
   REGISTERS_reg_21_22_inst : DFF_X1 port map( D => n6035, CK => CLK, Q => 
                           n19964, QN => n15447);
   REGISTERS_reg_21_21_inst : DFF_X1 port map( D => n6034, CK => CLK, Q => 
                           n19963, QN => n15448);
   REGISTERS_reg_21_20_inst : DFF_X1 port map( D => n6033, CK => CLK, Q => 
                           n19962, QN => n15449);
   REGISTERS_reg_21_19_inst : DFF_X1 port map( D => n6032, CK => CLK, Q => 
                           n19961, QN => n15450);
   REGISTERS_reg_21_18_inst : DFF_X1 port map( D => n6031, CK => CLK, Q => 
                           n19960, QN => n15451);
   REGISTERS_reg_21_17_inst : DFF_X1 port map( D => n6030, CK => CLK, Q => 
                           n19959, QN => n15452);
   REGISTERS_reg_21_16_inst : DFF_X1 port map( D => n6029, CK => CLK, Q => 
                           n19958, QN => n15453);
   REGISTERS_reg_21_15_inst : DFF_X1 port map( D => n6028, CK => CLK, Q => 
                           n19957, QN => n15454);
   REGISTERS_reg_21_14_inst : DFF_X1 port map( D => n6027, CK => CLK, Q => 
                           n19956, QN => n15455);
   REGISTERS_reg_21_13_inst : DFF_X1 port map( D => n6026, CK => CLK, Q => 
                           n19955, QN => n15456);
   REGISTERS_reg_21_12_inst : DFF_X1 port map( D => n6025, CK => CLK, Q => 
                           n19954, QN => n15457);
   REGISTERS_reg_21_11_inst : DFF_X1 port map( D => n6024, CK => CLK, Q => 
                           n19953, QN => n15458);
   REGISTERS_reg_21_10_inst : DFF_X1 port map( D => n6023, CK => CLK, Q => 
                           n19952, QN => n15459);
   REGISTERS_reg_21_9_inst : DFF_X1 port map( D => n6022, CK => CLK, Q => 
                           n19951, QN => n15460);
   REGISTERS_reg_21_8_inst : DFF_X1 port map( D => n6021, CK => CLK, Q => 
                           n19950, QN => n15461);
   REGISTERS_reg_21_7_inst : DFF_X1 port map( D => n6020, CK => CLK, Q => 
                           n19949, QN => n15462);
   REGISTERS_reg_21_6_inst : DFF_X1 port map( D => n6019, CK => CLK, Q => 
                           n19948, QN => n15463);
   REGISTERS_reg_21_5_inst : DFF_X1 port map( D => n6018, CK => CLK, Q => 
                           n19947, QN => n15464);
   REGISTERS_reg_21_4_inst : DFF_X1 port map( D => n6017, CK => CLK, Q => 
                           n19946, QN => n15465);
   REGISTERS_reg_21_3_inst : DFF_X1 port map( D => n6016, CK => CLK, Q => 
                           n19945, QN => n15466);
   REGISTERS_reg_21_2_inst : DFF_X1 port map( D => n6015, CK => CLK, Q => 
                           n19944, QN => n15467);
   REGISTERS_reg_21_1_inst : DFF_X1 port map( D => n6014, CK => CLK, Q => 
                           n19943, QN => n15468);
   REGISTERS_reg_21_0_inst : DFF_X1 port map( D => n6013, CK => CLK, Q => 
                           n19942, QN => n15469);
   REGISTERS_reg_20_59_inst : DFF_X1 port map( D => n6136, CK => CLK, Q => 
                           n18621, QN => n15344);
   REGISTERS_reg_20_58_inst : DFF_X1 port map( D => n6135, CK => CLK, Q => 
                           n18641, QN => n15345);
   REGISTERS_reg_20_57_inst : DFF_X1 port map( D => n6134, CK => CLK, Q => 
                           n18661, QN => n15346);
   REGISTERS_reg_20_56_inst : DFF_X1 port map( D => n6133, CK => CLK, Q => 
                           n18681, QN => n15347);
   REGISTERS_reg_20_55_inst : DFF_X1 port map( D => n6132, CK => CLK, Q => 
                           n18701, QN => n15348);
   REGISTERS_reg_20_54_inst : DFF_X1 port map( D => n6131, CK => CLK, Q => 
                           n18721, QN => n15349);
   REGISTERS_reg_20_53_inst : DFF_X1 port map( D => n6130, CK => CLK, Q => 
                           n18741, QN => n15350);
   REGISTERS_reg_20_52_inst : DFF_X1 port map( D => n6129, CK => CLK, Q => 
                           n18761, QN => n15351);
   REGISTERS_reg_20_51_inst : DFF_X1 port map( D => n6128, CK => CLK, Q => 
                           n18781, QN => n15352);
   REGISTERS_reg_20_50_inst : DFF_X1 port map( D => n6127, CK => CLK, Q => 
                           n18801, QN => n15353);
   REGISTERS_reg_20_49_inst : DFF_X1 port map( D => n6126, CK => CLK, Q => 
                           n18821, QN => n15354);
   REGISTERS_reg_20_48_inst : DFF_X1 port map( D => n6125, CK => CLK, Q => 
                           n18841, QN => n15355);
   REGISTERS_reg_20_47_inst : DFF_X1 port map( D => n6124, CK => CLK, Q => 
                           n18861, QN => n15356);
   REGISTERS_reg_20_46_inst : DFF_X1 port map( D => n6123, CK => CLK, Q => 
                           n18881, QN => n15357);
   REGISTERS_reg_20_45_inst : DFF_X1 port map( D => n6122, CK => CLK, Q => 
                           n18901, QN => n15358);
   REGISTERS_reg_20_44_inst : DFF_X1 port map( D => n6121, CK => CLK, Q => 
                           n18921, QN => n15359);
   REGISTERS_reg_20_43_inst : DFF_X1 port map( D => n6120, CK => CLK, Q => 
                           n18941, QN => n15360);
   REGISTERS_reg_20_42_inst : DFF_X1 port map( D => n6119, CK => CLK, Q => 
                           n18961, QN => n15361);
   REGISTERS_reg_20_41_inst : DFF_X1 port map( D => n6118, CK => CLK, Q => 
                           n18981, QN => n15362);
   REGISTERS_reg_20_40_inst : DFF_X1 port map( D => n6117, CK => CLK, Q => 
                           n19001, QN => n15363);
   REGISTERS_reg_20_39_inst : DFF_X1 port map( D => n6116, CK => CLK, Q => 
                           n19021, QN => n15364);
   REGISTERS_reg_20_38_inst : DFF_X1 port map( D => n6115, CK => CLK, Q => 
                           n19041, QN => n15365);
   REGISTERS_reg_20_37_inst : DFF_X1 port map( D => n6114, CK => CLK, Q => 
                           n19061, QN => n15366);
   REGISTERS_reg_20_36_inst : DFF_X1 port map( D => n6113, CK => CLK, Q => 
                           n19081, QN => n15367);
   REGISTERS_reg_20_35_inst : DFF_X1 port map( D => n6112, CK => CLK, Q => 
                           n19101, QN => n15368);
   REGISTERS_reg_20_34_inst : DFF_X1 port map( D => n6111, CK => CLK, Q => 
                           n19121, QN => n15369);
   REGISTERS_reg_20_33_inst : DFF_X1 port map( D => n6110, CK => CLK, Q => 
                           n19141, QN => n15370);
   REGISTERS_reg_20_32_inst : DFF_X1 port map( D => n6109, CK => CLK, Q => 
                           n19161, QN => n15371);
   REGISTERS_reg_20_31_inst : DFF_X1 port map( D => n6108, CK => CLK, Q => 
                           n19181, QN => n15372);
   REGISTERS_reg_20_30_inst : DFF_X1 port map( D => n6107, CK => CLK, Q => 
                           n19201, QN => n15373);
   REGISTERS_reg_20_29_inst : DFF_X1 port map( D => n6106, CK => CLK, Q => 
                           n19221, QN => n15374);
   REGISTERS_reg_20_28_inst : DFF_X1 port map( D => n6105, CK => CLK, Q => 
                           n19241, QN => n15375);
   REGISTERS_reg_20_27_inst : DFF_X1 port map( D => n6104, CK => CLK, Q => 
                           n19261, QN => n15376);
   REGISTERS_reg_20_26_inst : DFF_X1 port map( D => n6103, CK => CLK, Q => 
                           n19281, QN => n15377);
   REGISTERS_reg_20_25_inst : DFF_X1 port map( D => n6102, CK => CLK, Q => 
                           n19301, QN => n15378);
   REGISTERS_reg_20_24_inst : DFF_X1 port map( D => n6101, CK => CLK, Q => 
                           n19321, QN => n15379);
   REGISTERS_reg_20_23_inst : DFF_X1 port map( D => n6100, CK => CLK, Q => 
                           n19341, QN => n15380);
   REGISTERS_reg_20_22_inst : DFF_X1 port map( D => n6099, CK => CLK, Q => 
                           n19361, QN => n15381);
   REGISTERS_reg_20_21_inst : DFF_X1 port map( D => n6098, CK => CLK, Q => 
                           n19381, QN => n15382);
   REGISTERS_reg_20_20_inst : DFF_X1 port map( D => n6097, CK => CLK, Q => 
                           n19401, QN => n15383);
   REGISTERS_reg_20_19_inst : DFF_X1 port map( D => n6096, CK => CLK, Q => 
                           n19421, QN => n15384);
   REGISTERS_reg_20_18_inst : DFF_X1 port map( D => n6095, CK => CLK, Q => 
                           n19441, QN => n15385);
   REGISTERS_reg_20_17_inst : DFF_X1 port map( D => n6094, CK => CLK, Q => 
                           n19461, QN => n15386);
   REGISTERS_reg_20_16_inst : DFF_X1 port map( D => n6093, CK => CLK, Q => 
                           n19481, QN => n15387);
   REGISTERS_reg_20_15_inst : DFF_X1 port map( D => n6092, CK => CLK, Q => 
                           n19501, QN => n15388);
   REGISTERS_reg_20_14_inst : DFF_X1 port map( D => n6091, CK => CLK, Q => 
                           n19521, QN => n15389);
   REGISTERS_reg_20_13_inst : DFF_X1 port map( D => n6090, CK => CLK, Q => 
                           n19541, QN => n15390);
   REGISTERS_reg_20_12_inst : DFF_X1 port map( D => n6089, CK => CLK, Q => 
                           n19561, QN => n15391);
   REGISTERS_reg_20_11_inst : DFF_X1 port map( D => n6088, CK => CLK, Q => 
                           n19581, QN => n15392);
   REGISTERS_reg_20_10_inst : DFF_X1 port map( D => n6087, CK => CLK, Q => 
                           n19601, QN => n15393);
   REGISTERS_reg_20_9_inst : DFF_X1 port map( D => n6086, CK => CLK, Q => 
                           n19621, QN => n15394);
   REGISTERS_reg_20_8_inst : DFF_X1 port map( D => n6085, CK => CLK, Q => 
                           n19641, QN => n15395);
   REGISTERS_reg_20_7_inst : DFF_X1 port map( D => n6084, CK => CLK, Q => 
                           n19661, QN => n15396);
   REGISTERS_reg_20_6_inst : DFF_X1 port map( D => n6083, CK => CLK, Q => 
                           n19681, QN => n15397);
   REGISTERS_reg_20_5_inst : DFF_X1 port map( D => n6082, CK => CLK, Q => 
                           n19701, QN => n15398);
   REGISTERS_reg_20_4_inst : DFF_X1 port map( D => n6081, CK => CLK, Q => 
                           n19721, QN => n15399);
   REGISTERS_reg_20_3_inst : DFF_X1 port map( D => n6080, CK => CLK, Q => 
                           n19741, QN => n15400);
   REGISTERS_reg_20_2_inst : DFF_X1 port map( D => n6079, CK => CLK, Q => 
                           n19761, QN => n15401);
   REGISTERS_reg_20_1_inst : DFF_X1 port map( D => n6078, CK => CLK, Q => 
                           n19781, QN => n15402);
   REGISTERS_reg_20_0_inst : DFF_X1 port map( D => n6077, CK => CLK, Q => 
                           n19801, QN => n15403);
   REGISTERS_reg_19_59_inst : DFF_X1 port map( D => n6200, CK => CLK, Q => 
                           n19941, QN => n15278);
   REGISTERS_reg_19_58_inst : DFF_X1 port map( D => n6199, CK => CLK, Q => 
                           n19940, QN => n15279);
   REGISTERS_reg_19_57_inst : DFF_X1 port map( D => n6198, CK => CLK, Q => 
                           n19939, QN => n15280);
   REGISTERS_reg_19_56_inst : DFF_X1 port map( D => n6197, CK => CLK, Q => 
                           n19938, QN => n15281);
   REGISTERS_reg_19_55_inst : DFF_X1 port map( D => n6196, CK => CLK, Q => 
                           n19937, QN => n15282);
   REGISTERS_reg_19_54_inst : DFF_X1 port map( D => n6195, CK => CLK, Q => 
                           n19936, QN => n15283);
   REGISTERS_reg_19_53_inst : DFF_X1 port map( D => n6194, CK => CLK, Q => 
                           n19935, QN => n15284);
   REGISTERS_reg_19_52_inst : DFF_X1 port map( D => n6193, CK => CLK, Q => 
                           n19934, QN => n15285);
   REGISTERS_reg_19_51_inst : DFF_X1 port map( D => n6192, CK => CLK, Q => 
                           n19933, QN => n15286);
   REGISTERS_reg_19_50_inst : DFF_X1 port map( D => n6191, CK => CLK, Q => 
                           n19932, QN => n15287);
   REGISTERS_reg_19_49_inst : DFF_X1 port map( D => n6190, CK => CLK, Q => 
                           n19931, QN => n15288);
   REGISTERS_reg_19_48_inst : DFF_X1 port map( D => n6189, CK => CLK, Q => 
                           n19930, QN => n15289);
   REGISTERS_reg_19_47_inst : DFF_X1 port map( D => n6188, CK => CLK, Q => 
                           n19929, QN => n15290);
   REGISTERS_reg_19_46_inst : DFF_X1 port map( D => n6187, CK => CLK, Q => 
                           n19928, QN => n15291);
   REGISTERS_reg_19_45_inst : DFF_X1 port map( D => n6186, CK => CLK, Q => 
                           n19927, QN => n15292);
   REGISTERS_reg_19_44_inst : DFF_X1 port map( D => n6185, CK => CLK, Q => 
                           n19926, QN => n15293);
   REGISTERS_reg_19_43_inst : DFF_X1 port map( D => n6184, CK => CLK, Q => 
                           n19925, QN => n15294);
   REGISTERS_reg_19_42_inst : DFF_X1 port map( D => n6183, CK => CLK, Q => 
                           n19924, QN => n15295);
   REGISTERS_reg_19_41_inst : DFF_X1 port map( D => n6182, CK => CLK, Q => 
                           n19923, QN => n15296);
   REGISTERS_reg_19_40_inst : DFF_X1 port map( D => n6181, CK => CLK, Q => 
                           n19922, QN => n15297);
   REGISTERS_reg_19_39_inst : DFF_X1 port map( D => n6180, CK => CLK, Q => 
                           n19921, QN => n15298);
   REGISTERS_reg_19_38_inst : DFF_X1 port map( D => n6179, CK => CLK, Q => 
                           n19920, QN => n15299);
   REGISTERS_reg_19_37_inst : DFF_X1 port map( D => n6178, CK => CLK, Q => 
                           n19919, QN => n15300);
   REGISTERS_reg_19_36_inst : DFF_X1 port map( D => n6177, CK => CLK, Q => 
                           n19918, QN => n15301);
   REGISTERS_reg_19_35_inst : DFF_X1 port map( D => n6176, CK => CLK, Q => 
                           n19917, QN => n15302);
   REGISTERS_reg_19_34_inst : DFF_X1 port map( D => n6175, CK => CLK, Q => 
                           n19916, QN => n15303);
   REGISTERS_reg_19_33_inst : DFF_X1 port map( D => n6174, CK => CLK, Q => 
                           n19915, QN => n15304);
   REGISTERS_reg_19_32_inst : DFF_X1 port map( D => n6173, CK => CLK, Q => 
                           n19914, QN => n15305);
   REGISTERS_reg_19_31_inst : DFF_X1 port map( D => n6172, CK => CLK, Q => 
                           n19913, QN => n15306);
   REGISTERS_reg_19_30_inst : DFF_X1 port map( D => n6171, CK => CLK, Q => 
                           n19912, QN => n15307);
   REGISTERS_reg_19_29_inst : DFF_X1 port map( D => n6170, CK => CLK, Q => 
                           n19911, QN => n15308);
   REGISTERS_reg_19_28_inst : DFF_X1 port map( D => n6169, CK => CLK, Q => 
                           n19910, QN => n15309);
   REGISTERS_reg_19_27_inst : DFF_X1 port map( D => n6168, CK => CLK, Q => 
                           n19909, QN => n15310);
   REGISTERS_reg_19_26_inst : DFF_X1 port map( D => n6167, CK => CLK, Q => 
                           n19908, QN => n15311);
   REGISTERS_reg_19_25_inst : DFF_X1 port map( D => n6166, CK => CLK, Q => 
                           n19907, QN => n15312);
   REGISTERS_reg_19_24_inst : DFF_X1 port map( D => n6165, CK => CLK, Q => 
                           n19906, QN => n15313);
   REGISTERS_reg_19_23_inst : DFF_X1 port map( D => n6164, CK => CLK, Q => 
                           n19905, QN => n15314);
   REGISTERS_reg_19_22_inst : DFF_X1 port map( D => n6163, CK => CLK, Q => 
                           n19904, QN => n15315);
   REGISTERS_reg_19_21_inst : DFF_X1 port map( D => n6162, CK => CLK, Q => 
                           n19903, QN => n15316);
   REGISTERS_reg_19_20_inst : DFF_X1 port map( D => n6161, CK => CLK, Q => 
                           n19902, QN => n15317);
   REGISTERS_reg_19_19_inst : DFF_X1 port map( D => n6160, CK => CLK, Q => 
                           n19901, QN => n15318);
   REGISTERS_reg_19_18_inst : DFF_X1 port map( D => n6159, CK => CLK, Q => 
                           n19900, QN => n15319);
   REGISTERS_reg_19_17_inst : DFF_X1 port map( D => n6158, CK => CLK, Q => 
                           n19899, QN => n15320);
   REGISTERS_reg_19_16_inst : DFF_X1 port map( D => n6157, CK => CLK, Q => 
                           n19898, QN => n15321);
   REGISTERS_reg_19_15_inst : DFF_X1 port map( D => n6156, CK => CLK, Q => 
                           n19897, QN => n15322);
   REGISTERS_reg_19_14_inst : DFF_X1 port map( D => n6155, CK => CLK, Q => 
                           n19896, QN => n15323);
   REGISTERS_reg_19_13_inst : DFF_X1 port map( D => n6154, CK => CLK, Q => 
                           n19895, QN => n15324);
   REGISTERS_reg_19_12_inst : DFF_X1 port map( D => n6153, CK => CLK, Q => 
                           n19894, QN => n15325);
   REGISTERS_reg_19_11_inst : DFF_X1 port map( D => n6152, CK => CLK, Q => 
                           n19893, QN => n15326);
   REGISTERS_reg_19_10_inst : DFF_X1 port map( D => n6151, CK => CLK, Q => 
                           n19892, QN => n15327);
   REGISTERS_reg_19_9_inst : DFF_X1 port map( D => n6150, CK => CLK, Q => 
                           n19891, QN => n15328);
   REGISTERS_reg_19_8_inst : DFF_X1 port map( D => n6149, CK => CLK, Q => 
                           n19890, QN => n15329);
   REGISTERS_reg_19_7_inst : DFF_X1 port map( D => n6148, CK => CLK, Q => 
                           n19889, QN => n15330);
   REGISTERS_reg_19_6_inst : DFF_X1 port map( D => n6147, CK => CLK, Q => 
                           n19888, QN => n15331);
   REGISTERS_reg_19_5_inst : DFF_X1 port map( D => n6146, CK => CLK, Q => 
                           n19887, QN => n15332);
   REGISTERS_reg_19_4_inst : DFF_X1 port map( D => n6145, CK => CLK, Q => 
                           n19886, QN => n15333);
   REGISTERS_reg_19_3_inst : DFF_X1 port map( D => n6144, CK => CLK, Q => 
                           n19885, QN => n15334);
   REGISTERS_reg_19_2_inst : DFF_X1 port map( D => n6143, CK => CLK, Q => 
                           n19884, QN => n15335);
   REGISTERS_reg_19_1_inst : DFF_X1 port map( D => n6142, CK => CLK, Q => 
                           n19883, QN => n15336);
   REGISTERS_reg_19_0_inst : DFF_X1 port map( D => n6141, CK => CLK, Q => 
                           n19882, QN => n15337);
   REGISTERS_reg_18_59_inst : DFF_X1 port map( D => n6264, CK => CLK, Q => 
                           n8838, QN => n15212);
   REGISTERS_reg_18_58_inst : DFF_X1 port map( D => n6263, CK => CLK, Q => 
                           n8840, QN => n15213);
   REGISTERS_reg_18_57_inst : DFF_X1 port map( D => n6262, CK => CLK, Q => 
                           n8842, QN => n15214);
   REGISTERS_reg_18_56_inst : DFF_X1 port map( D => n6261, CK => CLK, Q => 
                           n8844, QN => n15215);
   REGISTERS_reg_18_55_inst : DFF_X1 port map( D => n6260, CK => CLK, Q => 
                           n8846, QN => n15216);
   REGISTERS_reg_18_54_inst : DFF_X1 port map( D => n6259, CK => CLK, Q => 
                           n8848, QN => n15217);
   REGISTERS_reg_18_53_inst : DFF_X1 port map( D => n6258, CK => CLK, Q => 
                           n8850, QN => n15218);
   REGISTERS_reg_18_52_inst : DFF_X1 port map( D => n6257, CK => CLK, Q => 
                           n8852, QN => n15219);
   REGISTERS_reg_18_51_inst : DFF_X1 port map( D => n6256, CK => CLK, Q => 
                           n8854, QN => n15220);
   REGISTERS_reg_18_50_inst : DFF_X1 port map( D => n6255, CK => CLK, Q => 
                           n8856, QN => n15221);
   REGISTERS_reg_18_49_inst : DFF_X1 port map( D => n6254, CK => CLK, Q => 
                           n8858, QN => n15222);
   REGISTERS_reg_18_48_inst : DFF_X1 port map( D => n6253, CK => CLK, Q => 
                           n8860, QN => n15223);
   REGISTERS_reg_18_47_inst : DFF_X1 port map( D => n6252, CK => CLK, Q => 
                           n8862, QN => n15224);
   REGISTERS_reg_18_46_inst : DFF_X1 port map( D => n6251, CK => CLK, Q => 
                           n8864, QN => n15225);
   REGISTERS_reg_18_45_inst : DFF_X1 port map( D => n6250, CK => CLK, Q => 
                           n8866, QN => n15226);
   REGISTERS_reg_18_44_inst : DFF_X1 port map( D => n6249, CK => CLK, Q => 
                           n8868, QN => n15227);
   REGISTERS_reg_18_43_inst : DFF_X1 port map( D => n6248, CK => CLK, Q => 
                           n8870, QN => n15228);
   REGISTERS_reg_18_42_inst : DFF_X1 port map( D => n6247, CK => CLK, Q => 
                           n8872, QN => n15229);
   REGISTERS_reg_18_41_inst : DFF_X1 port map( D => n6246, CK => CLK, Q => 
                           n8874, QN => n15230);
   REGISTERS_reg_18_40_inst : DFF_X1 port map( D => n6245, CK => CLK, Q => 
                           n8876, QN => n15231);
   REGISTERS_reg_18_39_inst : DFF_X1 port map( D => n6244, CK => CLK, Q => 
                           n8878, QN => n15232);
   REGISTERS_reg_18_38_inst : DFF_X1 port map( D => n6243, CK => CLK, Q => 
                           n8880, QN => n15233);
   REGISTERS_reg_18_37_inst : DFF_X1 port map( D => n6242, CK => CLK, Q => 
                           n8882, QN => n15234);
   REGISTERS_reg_18_36_inst : DFF_X1 port map( D => n6241, CK => CLK, Q => 
                           n8884, QN => n15235);
   REGISTERS_reg_18_35_inst : DFF_X1 port map( D => n6240, CK => CLK, Q => 
                           n8886, QN => n15236);
   REGISTERS_reg_18_34_inst : DFF_X1 port map( D => n6239, CK => CLK, Q => 
                           n8888, QN => n15237);
   REGISTERS_reg_18_33_inst : DFF_X1 port map( D => n6238, CK => CLK, Q => 
                           n8890, QN => n15238);
   REGISTERS_reg_18_32_inst : DFF_X1 port map( D => n6237, CK => CLK, Q => 
                           n8892, QN => n15239);
   REGISTERS_reg_18_31_inst : DFF_X1 port map( D => n6236, CK => CLK, Q => 
                           n8894, QN => n15240);
   REGISTERS_reg_18_30_inst : DFF_X1 port map( D => n6235, CK => CLK, Q => 
                           n8896, QN => n15241);
   REGISTERS_reg_18_29_inst : DFF_X1 port map( D => n6234, CK => CLK, Q => 
                           n8898, QN => n15242);
   REGISTERS_reg_18_28_inst : DFF_X1 port map( D => n6233, CK => CLK, Q => 
                           n8900, QN => n15243);
   REGISTERS_reg_18_27_inst : DFF_X1 port map( D => n6232, CK => CLK, Q => 
                           n8902, QN => n15244);
   REGISTERS_reg_18_26_inst : DFF_X1 port map( D => n6231, CK => CLK, Q => 
                           n8904, QN => n15245);
   REGISTERS_reg_18_25_inst : DFF_X1 port map( D => n6230, CK => CLK, Q => 
                           n8906, QN => n15246);
   REGISTERS_reg_18_24_inst : DFF_X1 port map( D => n6229, CK => CLK, Q => 
                           n8908, QN => n15247);
   REGISTERS_reg_18_23_inst : DFF_X1 port map( D => n6228, CK => CLK, Q => 
                           n8910, QN => n15248);
   REGISTERS_reg_18_22_inst : DFF_X1 port map( D => n6227, CK => CLK, Q => 
                           n8912, QN => n15249);
   REGISTERS_reg_18_21_inst : DFF_X1 port map( D => n6226, CK => CLK, Q => 
                           n8914, QN => n15250);
   REGISTERS_reg_18_20_inst : DFF_X1 port map( D => n6225, CK => CLK, Q => 
                           n8916, QN => n15251);
   REGISTERS_reg_18_19_inst : DFF_X1 port map( D => n6224, CK => CLK, Q => 
                           n8918, QN => n15252);
   REGISTERS_reg_18_18_inst : DFF_X1 port map( D => n6223, CK => CLK, Q => 
                           n8920, QN => n15253);
   REGISTERS_reg_18_17_inst : DFF_X1 port map( D => n6222, CK => CLK, Q => 
                           n8922, QN => n15254);
   REGISTERS_reg_18_16_inst : DFF_X1 port map( D => n6221, CK => CLK, Q => 
                           n8924, QN => n15255);
   REGISTERS_reg_18_15_inst : DFF_X1 port map( D => n6220, CK => CLK, Q => 
                           n8926, QN => n15256);
   REGISTERS_reg_18_14_inst : DFF_X1 port map( D => n6219, CK => CLK, Q => 
                           n8928, QN => n15257);
   REGISTERS_reg_18_13_inst : DFF_X1 port map( D => n6218, CK => CLK, Q => 
                           n8930, QN => n15258);
   REGISTERS_reg_18_12_inst : DFF_X1 port map( D => n6217, CK => CLK, Q => 
                           n8932, QN => n15259);
   REGISTERS_reg_18_11_inst : DFF_X1 port map( D => n6216, CK => CLK, Q => 
                           n8934, QN => n15260);
   REGISTERS_reg_18_10_inst : DFF_X1 port map( D => n6215, CK => CLK, Q => 
                           n8936, QN => n15261);
   REGISTERS_reg_18_9_inst : DFF_X1 port map( D => n6214, CK => CLK, Q => n8938
                           , QN => n15262);
   REGISTERS_reg_18_8_inst : DFF_X1 port map( D => n6213, CK => CLK, Q => n8940
                           , QN => n15263);
   REGISTERS_reg_18_7_inst : DFF_X1 port map( D => n6212, CK => CLK, Q => n8942
                           , QN => n15264);
   REGISTERS_reg_18_6_inst : DFF_X1 port map( D => n6211, CK => CLK, Q => n8944
                           , QN => n15265);
   REGISTERS_reg_18_5_inst : DFF_X1 port map( D => n6210, CK => CLK, Q => n8946
                           , QN => n15266);
   REGISTERS_reg_18_4_inst : DFF_X1 port map( D => n6209, CK => CLK, Q => n8948
                           , QN => n15267);
   REGISTERS_reg_18_3_inst : DFF_X1 port map( D => n6208, CK => CLK, Q => n8950
                           , QN => n15268);
   REGISTERS_reg_18_2_inst : DFF_X1 port map( D => n6207, CK => CLK, Q => n8952
                           , QN => n15269);
   REGISTERS_reg_18_1_inst : DFF_X1 port map( D => n6206, CK => CLK, Q => n8954
                           , QN => n15270);
   REGISTERS_reg_18_0_inst : DFF_X1 port map( D => n6205, CK => CLK, Q => n8956
                           , QN => n15271);
   REGISTERS_reg_24_59_inst : DFF_X1 port map( D => n5880, CK => CLK, Q => 
                           n19881, QN => n15609);
   REGISTERS_reg_24_58_inst : DFF_X1 port map( D => n5879, CK => CLK, Q => 
                           n19880, QN => n15610);
   REGISTERS_reg_24_57_inst : DFF_X1 port map( D => n5878, CK => CLK, Q => 
                           n19879, QN => n15611);
   REGISTERS_reg_24_56_inst : DFF_X1 port map( D => n5877, CK => CLK, Q => 
                           n19878, QN => n15612);
   REGISTERS_reg_24_55_inst : DFF_X1 port map( D => n5876, CK => CLK, Q => 
                           n19877, QN => n15613);
   REGISTERS_reg_24_54_inst : DFF_X1 port map( D => n5875, CK => CLK, Q => 
                           n19876, QN => n15614);
   REGISTERS_reg_24_53_inst : DFF_X1 port map( D => n5874, CK => CLK, Q => 
                           n19875, QN => n15615);
   REGISTERS_reg_24_52_inst : DFF_X1 port map( D => n5873, CK => CLK, Q => 
                           n19874, QN => n15616);
   REGISTERS_reg_24_51_inst : DFF_X1 port map( D => n5872, CK => CLK, Q => 
                           n19873, QN => n15617);
   REGISTERS_reg_24_50_inst : DFF_X1 port map( D => n5871, CK => CLK, Q => 
                           n19872, QN => n15618);
   REGISTERS_reg_24_49_inst : DFF_X1 port map( D => n5870, CK => CLK, Q => 
                           n19871, QN => n15619);
   REGISTERS_reg_24_48_inst : DFF_X1 port map( D => n5869, CK => CLK, Q => 
                           n19870, QN => n15620);
   REGISTERS_reg_24_47_inst : DFF_X1 port map( D => n5868, CK => CLK, Q => 
                           n19869, QN => n15621);
   REGISTERS_reg_24_46_inst : DFF_X1 port map( D => n5867, CK => CLK, Q => 
                           n19868, QN => n15622);
   REGISTERS_reg_24_45_inst : DFF_X1 port map( D => n5866, CK => CLK, Q => 
                           n19867, QN => n15623);
   REGISTERS_reg_24_44_inst : DFF_X1 port map( D => n5865, CK => CLK, Q => 
                           n19866, QN => n15624);
   REGISTERS_reg_24_43_inst : DFF_X1 port map( D => n5864, CK => CLK, Q => 
                           n19865, QN => n15625);
   REGISTERS_reg_24_42_inst : DFF_X1 port map( D => n5863, CK => CLK, Q => 
                           n19864, QN => n15626);
   REGISTERS_reg_24_41_inst : DFF_X1 port map( D => n5862, CK => CLK, Q => 
                           n19863, QN => n15627);
   REGISTERS_reg_24_40_inst : DFF_X1 port map( D => n5861, CK => CLK, Q => 
                           n19862, QN => n15628);
   REGISTERS_reg_24_39_inst : DFF_X1 port map( D => n5860, CK => CLK, Q => 
                           n19861, QN => n15629);
   REGISTERS_reg_24_38_inst : DFF_X1 port map( D => n5859, CK => CLK, Q => 
                           n19860, QN => n15630);
   REGISTERS_reg_24_37_inst : DFF_X1 port map( D => n5858, CK => CLK, Q => 
                           n19859, QN => n15631);
   REGISTERS_reg_24_36_inst : DFF_X1 port map( D => n5857, CK => CLK, Q => 
                           n19858, QN => n15632);
   REGISTERS_reg_24_35_inst : DFF_X1 port map( D => n5856, CK => CLK, Q => 
                           n19857, QN => n15633);
   REGISTERS_reg_24_34_inst : DFF_X1 port map( D => n5855, CK => CLK, Q => 
                           n19856, QN => n15634);
   REGISTERS_reg_24_33_inst : DFF_X1 port map( D => n5854, CK => CLK, Q => 
                           n19855, QN => n15635);
   REGISTERS_reg_24_32_inst : DFF_X1 port map( D => n5853, CK => CLK, Q => 
                           n19854, QN => n15636);
   REGISTERS_reg_24_31_inst : DFF_X1 port map( D => n5852, CK => CLK, Q => 
                           n19853, QN => n15637);
   REGISTERS_reg_24_30_inst : DFF_X1 port map( D => n5851, CK => CLK, Q => 
                           n19852, QN => n15638);
   REGISTERS_reg_24_29_inst : DFF_X1 port map( D => n5850, CK => CLK, Q => 
                           n19851, QN => n15639);
   REGISTERS_reg_24_28_inst : DFF_X1 port map( D => n5849, CK => CLK, Q => 
                           n19850, QN => n15640);
   REGISTERS_reg_24_27_inst : DFF_X1 port map( D => n5848, CK => CLK, Q => 
                           n19849, QN => n15641);
   REGISTERS_reg_24_26_inst : DFF_X1 port map( D => n5847, CK => CLK, Q => 
                           n19848, QN => n15642);
   REGISTERS_reg_24_25_inst : DFF_X1 port map( D => n5846, CK => CLK, Q => 
                           n19847, QN => n15643);
   REGISTERS_reg_24_24_inst : DFF_X1 port map( D => n5845, CK => CLK, Q => 
                           n19846, QN => n15644);
   REGISTERS_reg_24_23_inst : DFF_X1 port map( D => n5844, CK => CLK, Q => 
                           n19845, QN => n15645);
   REGISTERS_reg_24_22_inst : DFF_X1 port map( D => n5843, CK => CLK, Q => 
                           n19844, QN => n15646);
   REGISTERS_reg_24_21_inst : DFF_X1 port map( D => n5842, CK => CLK, Q => 
                           n19843, QN => n15647);
   REGISTERS_reg_24_20_inst : DFF_X1 port map( D => n5841, CK => CLK, Q => 
                           n19842, QN => n15648);
   REGISTERS_reg_24_19_inst : DFF_X1 port map( D => n5840, CK => CLK, Q => 
                           n19841, QN => n15649);
   REGISTERS_reg_24_18_inst : DFF_X1 port map( D => n5839, CK => CLK, Q => 
                           n19840, QN => n15650);
   REGISTERS_reg_24_17_inst : DFF_X1 port map( D => n5838, CK => CLK, Q => 
                           n19839, QN => n15651);
   REGISTERS_reg_24_16_inst : DFF_X1 port map( D => n5837, CK => CLK, Q => 
                           n19838, QN => n15652);
   REGISTERS_reg_24_15_inst : DFF_X1 port map( D => n5836, CK => CLK, Q => 
                           n19837, QN => n15653);
   REGISTERS_reg_24_14_inst : DFF_X1 port map( D => n5835, CK => CLK, Q => 
                           n19836, QN => n15654);
   REGISTERS_reg_24_13_inst : DFF_X1 port map( D => n5834, CK => CLK, Q => 
                           n19835, QN => n15655);
   REGISTERS_reg_24_12_inst : DFF_X1 port map( D => n5833, CK => CLK, Q => 
                           n19834, QN => n15656);
   REGISTERS_reg_24_11_inst : DFF_X1 port map( D => n5832, CK => CLK, Q => 
                           n19833, QN => n15657);
   REGISTERS_reg_24_10_inst : DFF_X1 port map( D => n5831, CK => CLK, Q => 
                           n19832, QN => n15658);
   REGISTERS_reg_24_9_inst : DFF_X1 port map( D => n5830, CK => CLK, Q => 
                           n19831, QN => n15659);
   REGISTERS_reg_24_8_inst : DFF_X1 port map( D => n5829, CK => CLK, Q => 
                           n19830, QN => n15660);
   REGISTERS_reg_24_7_inst : DFF_X1 port map( D => n5828, CK => CLK, Q => 
                           n19829, QN => n15661);
   REGISTERS_reg_24_6_inst : DFF_X1 port map( D => n5827, CK => CLK, Q => 
                           n19828, QN => n15662);
   REGISTERS_reg_24_5_inst : DFF_X1 port map( D => n5826, CK => CLK, Q => 
                           n19827, QN => n15663);
   REGISTERS_reg_24_4_inst : DFF_X1 port map( D => n5825, CK => CLK, Q => 
                           n19826, QN => n15664);
   REGISTERS_reg_24_3_inst : DFF_X1 port map( D => n5824, CK => CLK, Q => 
                           n19825, QN => n15665);
   REGISTERS_reg_24_2_inst : DFF_X1 port map( D => n5823, CK => CLK, Q => 
                           n19824, QN => n15666);
   REGISTERS_reg_24_1_inst : DFF_X1 port map( D => n5822, CK => CLK, Q => 
                           n19823, QN => n15667);
   REGISTERS_reg_24_0_inst : DFF_X1 port map( D => n5821, CK => CLK, Q => 
                           n19822, QN => n15668);
   REGISTERS_reg_17_59_inst : DFF_X1 port map( D => n6328, CK => CLK, Q => 
                           n18634, QN => n15145);
   REGISTERS_reg_17_58_inst : DFF_X1 port map( D => n6327, CK => CLK, Q => 
                           n18654, QN => n15146);
   REGISTERS_reg_17_57_inst : DFF_X1 port map( D => n6326, CK => CLK, Q => 
                           n18674, QN => n15147);
   REGISTERS_reg_17_56_inst : DFF_X1 port map( D => n6325, CK => CLK, Q => 
                           n18694, QN => n15148);
   REGISTERS_reg_17_55_inst : DFF_X1 port map( D => n6324, CK => CLK, Q => 
                           n18714, QN => n15149);
   REGISTERS_reg_17_54_inst : DFF_X1 port map( D => n6323, CK => CLK, Q => 
                           n18734, QN => n15150);
   REGISTERS_reg_17_53_inst : DFF_X1 port map( D => n6322, CK => CLK, Q => 
                           n18754, QN => n15151);
   REGISTERS_reg_17_52_inst : DFF_X1 port map( D => n6321, CK => CLK, Q => 
                           n18774, QN => n15152);
   REGISTERS_reg_17_51_inst : DFF_X1 port map( D => n6320, CK => CLK, Q => 
                           n18794, QN => n15153);
   REGISTERS_reg_17_50_inst : DFF_X1 port map( D => n6319, CK => CLK, Q => 
                           n18814, QN => n15154);
   REGISTERS_reg_17_49_inst : DFF_X1 port map( D => n6318, CK => CLK, Q => 
                           n18834, QN => n15155);
   REGISTERS_reg_17_48_inst : DFF_X1 port map( D => n6317, CK => CLK, Q => 
                           n18854, QN => n15156);
   REGISTERS_reg_17_47_inst : DFF_X1 port map( D => n6316, CK => CLK, Q => 
                           n18874, QN => n15157);
   REGISTERS_reg_17_46_inst : DFF_X1 port map( D => n6315, CK => CLK, Q => 
                           n18894, QN => n15158);
   REGISTERS_reg_17_45_inst : DFF_X1 port map( D => n6314, CK => CLK, Q => 
                           n18914, QN => n15159);
   REGISTERS_reg_17_44_inst : DFF_X1 port map( D => n6313, CK => CLK, Q => 
                           n18934, QN => n15160);
   REGISTERS_reg_17_43_inst : DFF_X1 port map( D => n6312, CK => CLK, Q => 
                           n18954, QN => n15161);
   REGISTERS_reg_17_42_inst : DFF_X1 port map( D => n6311, CK => CLK, Q => 
                           n18974, QN => n15162);
   REGISTERS_reg_17_41_inst : DFF_X1 port map( D => n6310, CK => CLK, Q => 
                           n18994, QN => n15163);
   REGISTERS_reg_17_40_inst : DFF_X1 port map( D => n6309, CK => CLK, Q => 
                           n19014, QN => n15164);
   REGISTERS_reg_17_39_inst : DFF_X1 port map( D => n6308, CK => CLK, Q => 
                           n19034, QN => n15165);
   REGISTERS_reg_17_38_inst : DFF_X1 port map( D => n6307, CK => CLK, Q => 
                           n19054, QN => n15166);
   REGISTERS_reg_17_37_inst : DFF_X1 port map( D => n6306, CK => CLK, Q => 
                           n19074, QN => n15167);
   REGISTERS_reg_17_36_inst : DFF_X1 port map( D => n6305, CK => CLK, Q => 
                           n19094, QN => n15168);
   REGISTERS_reg_17_35_inst : DFF_X1 port map( D => n6304, CK => CLK, Q => 
                           n19114, QN => n15169);
   REGISTERS_reg_17_34_inst : DFF_X1 port map( D => n6303, CK => CLK, Q => 
                           n19134, QN => n15170);
   REGISTERS_reg_17_33_inst : DFF_X1 port map( D => n6302, CK => CLK, Q => 
                           n19154, QN => n15171);
   REGISTERS_reg_17_32_inst : DFF_X1 port map( D => n6301, CK => CLK, Q => 
                           n19174, QN => n15172);
   REGISTERS_reg_17_31_inst : DFF_X1 port map( D => n6300, CK => CLK, Q => 
                           n19194, QN => n15173);
   REGISTERS_reg_17_30_inst : DFF_X1 port map( D => n6299, CK => CLK, Q => 
                           n19214, QN => n15174);
   REGISTERS_reg_17_29_inst : DFF_X1 port map( D => n6298, CK => CLK, Q => 
                           n19234, QN => n15175);
   REGISTERS_reg_17_28_inst : DFF_X1 port map( D => n6297, CK => CLK, Q => 
                           n19254, QN => n15176);
   REGISTERS_reg_17_27_inst : DFF_X1 port map( D => n6296, CK => CLK, Q => 
                           n19274, QN => n15177);
   REGISTERS_reg_17_26_inst : DFF_X1 port map( D => n6295, CK => CLK, Q => 
                           n19294, QN => n15178);
   REGISTERS_reg_17_25_inst : DFF_X1 port map( D => n6294, CK => CLK, Q => 
                           n19314, QN => n15179);
   REGISTERS_reg_17_24_inst : DFF_X1 port map( D => n6293, CK => CLK, Q => 
                           n19334, QN => n15180);
   REGISTERS_reg_17_23_inst : DFF_X1 port map( D => n6292, CK => CLK, Q => 
                           n19354, QN => n15181);
   REGISTERS_reg_17_22_inst : DFF_X1 port map( D => n6291, CK => CLK, Q => 
                           n19374, QN => n15182);
   REGISTERS_reg_17_21_inst : DFF_X1 port map( D => n6290, CK => CLK, Q => 
                           n19394, QN => n15183);
   REGISTERS_reg_17_20_inst : DFF_X1 port map( D => n6289, CK => CLK, Q => 
                           n19414, QN => n15184);
   REGISTERS_reg_17_19_inst : DFF_X1 port map( D => n6288, CK => CLK, Q => 
                           n19434, QN => n15185);
   REGISTERS_reg_17_18_inst : DFF_X1 port map( D => n6287, CK => CLK, Q => 
                           n19454, QN => n15186);
   REGISTERS_reg_17_17_inst : DFF_X1 port map( D => n6286, CK => CLK, Q => 
                           n19474, QN => n15187);
   REGISTERS_reg_17_16_inst : DFF_X1 port map( D => n6285, CK => CLK, Q => 
                           n19494, QN => n15188);
   REGISTERS_reg_17_15_inst : DFF_X1 port map( D => n6284, CK => CLK, Q => 
                           n19514, QN => n15189);
   REGISTERS_reg_17_14_inst : DFF_X1 port map( D => n6283, CK => CLK, Q => 
                           n19534, QN => n15190);
   REGISTERS_reg_17_13_inst : DFF_X1 port map( D => n6282, CK => CLK, Q => 
                           n19554, QN => n15191);
   REGISTERS_reg_17_12_inst : DFF_X1 port map( D => n6281, CK => CLK, Q => 
                           n19574, QN => n15192);
   REGISTERS_reg_17_11_inst : DFF_X1 port map( D => n6280, CK => CLK, Q => 
                           n19594, QN => n15193);
   REGISTERS_reg_17_10_inst : DFF_X1 port map( D => n6279, CK => CLK, Q => 
                           n19614, QN => n15194);
   REGISTERS_reg_17_9_inst : DFF_X1 port map( D => n6278, CK => CLK, Q => 
                           n19634, QN => n15195);
   REGISTERS_reg_17_8_inst : DFF_X1 port map( D => n6277, CK => CLK, Q => 
                           n19654, QN => n15196);
   REGISTERS_reg_17_7_inst : DFF_X1 port map( D => n6276, CK => CLK, Q => 
                           n19674, QN => n15197);
   REGISTERS_reg_17_6_inst : DFF_X1 port map( D => n6275, CK => CLK, Q => 
                           n19694, QN => n15198);
   REGISTERS_reg_17_5_inst : DFF_X1 port map( D => n6274, CK => CLK, Q => 
                           n19714, QN => n15199);
   REGISTERS_reg_17_4_inst : DFF_X1 port map( D => n6273, CK => CLK, Q => 
                           n19734, QN => n15200);
   REGISTERS_reg_17_3_inst : DFF_X1 port map( D => n6272, CK => CLK, Q => 
                           n19754, QN => n15201);
   REGISTERS_reg_17_2_inst : DFF_X1 port map( D => n6271, CK => CLK, Q => 
                           n19774, QN => n15202);
   REGISTERS_reg_17_1_inst : DFF_X1 port map( D => n6270, CK => CLK, Q => 
                           n19794, QN => n15203);
   REGISTERS_reg_17_0_inst : DFF_X1 port map( D => n6269, CK => CLK, Q => 
                           n19814, QN => n15204);
   REGISTERS_reg_16_59_inst : DFF_X1 port map( D => n6392, CK => CLK, Q => 
                           n8589, QN => n15078);
   REGISTERS_reg_16_58_inst : DFF_X1 port map( D => n6391, CK => CLK, Q => 
                           n8593, QN => n15079);
   REGISTERS_reg_16_57_inst : DFF_X1 port map( D => n6390, CK => CLK, Q => 
                           n8597, QN => n15080);
   REGISTERS_reg_16_56_inst : DFF_X1 port map( D => n6389, CK => CLK, Q => 
                           n8601, QN => n15081);
   REGISTERS_reg_16_55_inst : DFF_X1 port map( D => n6388, CK => CLK, Q => 
                           n8605, QN => n15082);
   REGISTERS_reg_16_54_inst : DFF_X1 port map( D => n6387, CK => CLK, Q => 
                           n8609, QN => n15083);
   REGISTERS_reg_16_53_inst : DFF_X1 port map( D => n6386, CK => CLK, Q => 
                           n8613, QN => n15084);
   REGISTERS_reg_16_52_inst : DFF_X1 port map( D => n6385, CK => CLK, Q => 
                           n8617, QN => n15085);
   REGISTERS_reg_16_51_inst : DFF_X1 port map( D => n6384, CK => CLK, Q => 
                           n8621, QN => n15086);
   REGISTERS_reg_16_50_inst : DFF_X1 port map( D => n6383, CK => CLK, Q => 
                           n8625, QN => n15087);
   REGISTERS_reg_16_49_inst : DFF_X1 port map( D => n6382, CK => CLK, Q => 
                           n8629, QN => n15088);
   REGISTERS_reg_16_48_inst : DFF_X1 port map( D => n6381, CK => CLK, Q => 
                           n8633, QN => n15089);
   REGISTERS_reg_16_47_inst : DFF_X1 port map( D => n6380, CK => CLK, Q => 
                           n8637, QN => n15090);
   REGISTERS_reg_16_46_inst : DFF_X1 port map( D => n6379, CK => CLK, Q => 
                           n8641, QN => n15091);
   REGISTERS_reg_16_45_inst : DFF_X1 port map( D => n6378, CK => CLK, Q => 
                           n8645, QN => n15092);
   REGISTERS_reg_16_44_inst : DFF_X1 port map( D => n6377, CK => CLK, Q => 
                           n8649, QN => n15093);
   REGISTERS_reg_16_43_inst : DFF_X1 port map( D => n6376, CK => CLK, Q => 
                           n8653, QN => n15094);
   REGISTERS_reg_16_42_inst : DFF_X1 port map( D => n6375, CK => CLK, Q => 
                           n8657, QN => n15095);
   REGISTERS_reg_16_41_inst : DFF_X1 port map( D => n6374, CK => CLK, Q => 
                           n8661, QN => n15096);
   REGISTERS_reg_16_40_inst : DFF_X1 port map( D => n6373, CK => CLK, Q => 
                           n8665, QN => n15097);
   REGISTERS_reg_16_39_inst : DFF_X1 port map( D => n6372, CK => CLK, Q => 
                           n8669, QN => n15098);
   REGISTERS_reg_16_38_inst : DFF_X1 port map( D => n6371, CK => CLK, Q => 
                           n8673, QN => n15099);
   REGISTERS_reg_16_37_inst : DFF_X1 port map( D => n6370, CK => CLK, Q => 
                           n8677, QN => n15100);
   REGISTERS_reg_16_36_inst : DFF_X1 port map( D => n6369, CK => CLK, Q => 
                           n8681, QN => n15101);
   REGISTERS_reg_16_35_inst : DFF_X1 port map( D => n6368, CK => CLK, Q => 
                           n8685, QN => n15102);
   REGISTERS_reg_16_34_inst : DFF_X1 port map( D => n6367, CK => CLK, Q => 
                           n8689, QN => n15103);
   REGISTERS_reg_16_33_inst : DFF_X1 port map( D => n6366, CK => CLK, Q => 
                           n8693, QN => n15104);
   REGISTERS_reg_16_32_inst : DFF_X1 port map( D => n6365, CK => CLK, Q => 
                           n8697, QN => n15105);
   REGISTERS_reg_16_31_inst : DFF_X1 port map( D => n6364, CK => CLK, Q => 
                           n8701, QN => n15106);
   REGISTERS_reg_16_30_inst : DFF_X1 port map( D => n6363, CK => CLK, Q => 
                           n8705, QN => n15107);
   REGISTERS_reg_16_29_inst : DFF_X1 port map( D => n6362, CK => CLK, Q => 
                           n8709, QN => n15108);
   REGISTERS_reg_16_28_inst : DFF_X1 port map( D => n6361, CK => CLK, Q => 
                           n8713, QN => n15109);
   REGISTERS_reg_16_27_inst : DFF_X1 port map( D => n6360, CK => CLK, Q => 
                           n8717, QN => n15110);
   REGISTERS_reg_16_26_inst : DFF_X1 port map( D => n6359, CK => CLK, Q => 
                           n8721, QN => n15111);
   REGISTERS_reg_16_25_inst : DFF_X1 port map( D => n6358, CK => CLK, Q => 
                           n8725, QN => n15112);
   REGISTERS_reg_16_24_inst : DFF_X1 port map( D => n6357, CK => CLK, Q => 
                           n8729, QN => n15113);
   REGISTERS_reg_16_23_inst : DFF_X1 port map( D => n6356, CK => CLK, Q => 
                           n8733, QN => n15114);
   REGISTERS_reg_16_22_inst : DFF_X1 port map( D => n6355, CK => CLK, Q => 
                           n8737, QN => n15115);
   REGISTERS_reg_16_21_inst : DFF_X1 port map( D => n6354, CK => CLK, Q => 
                           n8741, QN => n15116);
   REGISTERS_reg_16_20_inst : DFF_X1 port map( D => n6353, CK => CLK, Q => 
                           n8745, QN => n15117);
   REGISTERS_reg_16_19_inst : DFF_X1 port map( D => n6352, CK => CLK, Q => 
                           n8749, QN => n15118);
   REGISTERS_reg_16_18_inst : DFF_X1 port map( D => n6351, CK => CLK, Q => 
                           n8753, QN => n15119);
   REGISTERS_reg_16_17_inst : DFF_X1 port map( D => n6350, CK => CLK, Q => 
                           n8757, QN => n15120);
   REGISTERS_reg_16_16_inst : DFF_X1 port map( D => n6349, CK => CLK, Q => 
                           n8761, QN => n15121);
   REGISTERS_reg_16_15_inst : DFF_X1 port map( D => n6348, CK => CLK, Q => 
                           n8765, QN => n15122);
   REGISTERS_reg_16_14_inst : DFF_X1 port map( D => n6347, CK => CLK, Q => 
                           n8769, QN => n15123);
   REGISTERS_reg_16_13_inst : DFF_X1 port map( D => n6346, CK => CLK, Q => 
                           n8773, QN => n15124);
   REGISTERS_reg_16_12_inst : DFF_X1 port map( D => n6345, CK => CLK, Q => 
                           n8777, QN => n15125);
   REGISTERS_reg_16_11_inst : DFF_X1 port map( D => n6344, CK => CLK, Q => 
                           n8781, QN => n15126);
   REGISTERS_reg_16_10_inst : DFF_X1 port map( D => n6343, CK => CLK, Q => 
                           n8785, QN => n15127);
   REGISTERS_reg_16_9_inst : DFF_X1 port map( D => n6342, CK => CLK, Q => n8789
                           , QN => n15128);
   REGISTERS_reg_16_8_inst : DFF_X1 port map( D => n6341, CK => CLK, Q => n8793
                           , QN => n15129);
   REGISTERS_reg_16_7_inst : DFF_X1 port map( D => n6340, CK => CLK, Q => n8797
                           , QN => n15130);
   REGISTERS_reg_16_6_inst : DFF_X1 port map( D => n6339, CK => CLK, Q => n8801
                           , QN => n15131);
   REGISTERS_reg_16_5_inst : DFF_X1 port map( D => n6338, CK => CLK, Q => n8805
                           , QN => n15132);
   REGISTERS_reg_16_4_inst : DFF_X1 port map( D => n6337, CK => CLK, Q => n8809
                           , QN => n15133);
   REGISTERS_reg_16_3_inst : DFF_X1 port map( D => n6336, CK => CLK, Q => n8813
                           , QN => n15134);
   REGISTERS_reg_16_2_inst : DFF_X1 port map( D => n6335, CK => CLK, Q => n8817
                           , QN => n15135);
   REGISTERS_reg_16_1_inst : DFF_X1 port map( D => n6334, CK => CLK, Q => n8821
                           , QN => n15136);
   REGISTERS_reg_16_0_inst : DFF_X1 port map( D => n6333, CK => CLK, Q => n8825
                           , QN => n15137);
   OUT2_reg_63_inst : DFF_X1 port map( D => n5308, CK => CLK, Q => OUT2_63_port
                           , QN => n19821);
   U13048 : NOR3_X1 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n20984,
                           ZN => n18520);
   U13049 : NOR3_X1 port map( A1 => n20984, A2 => ADD_RD2(2), A3 => n18538, ZN 
                           => n18531);
   U13050 : NOR3_X1 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n20984,
                           ZN => n17320);
   U13051 : NOR3_X1 port map( A1 => n20984, A2 => ADD_RD1(2), A3 => n17337, ZN 
                           => n17330);
   U13052 : NOR3_X1 port map( A1 => n20984, A2 => ADD_RD1(1), A3 => n17338, ZN 
                           => n17313);
   U13053 : NOR3_X1 port map( A1 => n18539, A2 => n20984, A3 => n18538, ZN => 
                           n18512);
   U13054 : NOR3_X1 port map( A1 => n20984, A2 => ADD_RD2(1), A3 => n18539, ZN 
                           => n18514);
   U13055 : BUF_X1 port map( A => n13941, Z => n21719);
   U13056 : BUF_X1 port map( A => n13941, Z => n21720);
   U13057 : BUF_X1 port map( A => n13941, Z => n21721);
   U13058 : BUF_X1 port map( A => n13941, Z => n21722);
   U13059 : BUF_X1 port map( A => n21317, Z => n21319);
   U13060 : BUF_X1 port map( A => n21724, Z => n21726);
   U13061 : BUF_X1 port map( A => n21317, Z => n21320);
   U13062 : BUF_X1 port map( A => n21317, Z => n21321);
   U13063 : BUF_X1 port map( A => n21318, Z => n21322);
   U13064 : BUF_X1 port map( A => n21318, Z => n21323);
   U13065 : BUF_X1 port map( A => n21724, Z => n21727);
   U13066 : BUF_X1 port map( A => n21724, Z => n21728);
   U13067 : BUF_X1 port map( A => n21725, Z => n21729);
   U13068 : BUF_X1 port map( A => n21725, Z => n21730);
   U13069 : BUF_X1 port map( A => n16071, Z => n21116);
   U13070 : BUF_X1 port map( A => n16071, Z => n21117);
   U13071 : BUF_X1 port map( A => n16071, Z => n21118);
   U13072 : BUF_X1 port map( A => n16071, Z => n21119);
   U13073 : BUF_X1 port map( A => n16071, Z => n21120);
   U13074 : BUF_X1 port map( A => n16005, Z => n21129);
   U13075 : BUF_X1 port map( A => n16005, Z => n21130);
   U13076 : BUF_X1 port map( A => n16005, Z => n21131);
   U13077 : BUF_X1 port map( A => n16005, Z => n21132);
   U13078 : BUF_X1 port map( A => n16005, Z => n21133);
   U13079 : BUF_X1 port map( A => n15939, Z => n21142);
   U13080 : BUF_X1 port map( A => n15939, Z => n21143);
   U13081 : BUF_X1 port map( A => n15939, Z => n21144);
   U13082 : BUF_X1 port map( A => n15939, Z => n21145);
   U13083 : BUF_X1 port map( A => n15939, Z => n21146);
   U13084 : BUF_X1 port map( A => n15873, Z => n21155);
   U13085 : BUF_X1 port map( A => n15873, Z => n21156);
   U13086 : BUF_X1 port map( A => n15873, Z => n21157);
   U13087 : BUF_X1 port map( A => n15873, Z => n21158);
   U13088 : BUF_X1 port map( A => n15873, Z => n21159);
   U13089 : BUF_X1 port map( A => n15807, Z => n21168);
   U13090 : BUF_X1 port map( A => n15807, Z => n21169);
   U13091 : BUF_X1 port map( A => n15807, Z => n21170);
   U13092 : BUF_X1 port map( A => n15807, Z => n21171);
   U13093 : BUF_X1 port map( A => n15807, Z => n21172);
   U13094 : BUF_X1 port map( A => n15741, Z => n21181);
   U13095 : BUF_X1 port map( A => n15741, Z => n21182);
   U13096 : BUF_X1 port map( A => n15741, Z => n21183);
   U13097 : BUF_X1 port map( A => n15741, Z => n21184);
   U13098 : BUF_X1 port map( A => n15741, Z => n21185);
   U13099 : BUF_X1 port map( A => n15672, Z => n21194);
   U13100 : BUF_X1 port map( A => n15672, Z => n21195);
   U13101 : BUF_X1 port map( A => n15672, Z => n21196);
   U13102 : BUF_X1 port map( A => n15672, Z => n21197);
   U13103 : BUF_X1 port map( A => n15672, Z => n21198);
   U13104 : BUF_X1 port map( A => n15605, Z => n21207);
   U13105 : BUF_X1 port map( A => n15605, Z => n21208);
   U13106 : BUF_X1 port map( A => n15605, Z => n21209);
   U13107 : BUF_X1 port map( A => n15605, Z => n21210);
   U13108 : BUF_X1 port map( A => n15605, Z => n21211);
   U13109 : BUF_X1 port map( A => n15539, Z => n21220);
   U13110 : BUF_X1 port map( A => n15539, Z => n21221);
   U13111 : BUF_X1 port map( A => n15539, Z => n21222);
   U13112 : BUF_X1 port map( A => n15539, Z => n21223);
   U13113 : BUF_X1 port map( A => n15539, Z => n21224);
   U13114 : BUF_X1 port map( A => n15472, Z => n21233);
   U13115 : BUF_X1 port map( A => n15472, Z => n21234);
   U13116 : BUF_X1 port map( A => n15472, Z => n21235);
   U13117 : BUF_X1 port map( A => n15472, Z => n21236);
   U13118 : BUF_X1 port map( A => n15472, Z => n21237);
   U13119 : BUF_X1 port map( A => n15406, Z => n21246);
   U13120 : BUF_X1 port map( A => n15406, Z => n21247);
   U13121 : BUF_X1 port map( A => n15406, Z => n21248);
   U13122 : BUF_X1 port map( A => n15406, Z => n21249);
   U13123 : BUF_X1 port map( A => n15406, Z => n21250);
   U13124 : BUF_X1 port map( A => n15340, Z => n21259);
   U13125 : BUF_X1 port map( A => n15340, Z => n21260);
   U13126 : BUF_X1 port map( A => n15340, Z => n21261);
   U13127 : BUF_X1 port map( A => n15340, Z => n21262);
   U13128 : BUF_X1 port map( A => n15340, Z => n21263);
   U13129 : BUF_X1 port map( A => n15274, Z => n21272);
   U13130 : BUF_X1 port map( A => n15274, Z => n21273);
   U13131 : BUF_X1 port map( A => n15274, Z => n21274);
   U13132 : BUF_X1 port map( A => n15274, Z => n21275);
   U13133 : BUF_X1 port map( A => n15274, Z => n21276);
   U13134 : BUF_X1 port map( A => n15208, Z => n21285);
   U13135 : BUF_X1 port map( A => n15208, Z => n21286);
   U13136 : BUF_X1 port map( A => n15208, Z => n21287);
   U13137 : BUF_X1 port map( A => n15208, Z => n21288);
   U13138 : BUF_X1 port map( A => n15208, Z => n21289);
   U13139 : BUF_X1 port map( A => n15141, Z => n21298);
   U13140 : BUF_X1 port map( A => n15141, Z => n21299);
   U13141 : BUF_X1 port map( A => n15141, Z => n21300);
   U13142 : BUF_X1 port map( A => n15141, Z => n21301);
   U13143 : BUF_X1 port map( A => n15141, Z => n21302);
   U13144 : BUF_X1 port map( A => n15074, Z => n21311);
   U13145 : BUF_X1 port map( A => n15074, Z => n21312);
   U13146 : BUF_X1 port map( A => n15074, Z => n21313);
   U13147 : BUF_X1 port map( A => n15074, Z => n21314);
   U13148 : BUF_X1 port map( A => n15074, Z => n21315);
   U13149 : BUF_X1 port map( A => n15007, Z => n21324);
   U13150 : BUF_X1 port map( A => n15007, Z => n21325);
   U13151 : BUF_X1 port map( A => n15007, Z => n21326);
   U13152 : BUF_X1 port map( A => n15007, Z => n21327);
   U13153 : BUF_X1 port map( A => n15007, Z => n21328);
   U13154 : BUF_X1 port map( A => n14941, Z => n21337);
   U13155 : BUF_X1 port map( A => n14941, Z => n21338);
   U13156 : BUF_X1 port map( A => n14941, Z => n21339);
   U13157 : BUF_X1 port map( A => n14941, Z => n21340);
   U13158 : BUF_X1 port map( A => n14941, Z => n21341);
   U13159 : BUF_X1 port map( A => n14875, Z => n21350);
   U13160 : BUF_X1 port map( A => n14875, Z => n21351);
   U13161 : BUF_X1 port map( A => n14875, Z => n21352);
   U13162 : BUF_X1 port map( A => n14875, Z => n21353);
   U13163 : BUF_X1 port map( A => n14875, Z => n21354);
   U13164 : BUF_X1 port map( A => n14809, Z => n21363);
   U13165 : BUF_X1 port map( A => n14809, Z => n21364);
   U13166 : BUF_X1 port map( A => n14809, Z => n21365);
   U13167 : BUF_X1 port map( A => n14809, Z => n21366);
   U13168 : BUF_X1 port map( A => n14809, Z => n21367);
   U13169 : BUF_X1 port map( A => n14743, Z => n21376);
   U13170 : BUF_X1 port map( A => n14743, Z => n21377);
   U13171 : BUF_X1 port map( A => n14743, Z => n21378);
   U13172 : BUF_X1 port map( A => n14743, Z => n21379);
   U13173 : BUF_X1 port map( A => n14743, Z => n21380);
   U13174 : BUF_X1 port map( A => n14677, Z => n21389);
   U13175 : BUF_X1 port map( A => n14677, Z => n21390);
   U13176 : BUF_X1 port map( A => n14677, Z => n21391);
   U13177 : BUF_X1 port map( A => n14677, Z => n21392);
   U13178 : BUF_X1 port map( A => n14677, Z => n21393);
   U13179 : BUF_X1 port map( A => n14610, Z => n21402);
   U13180 : BUF_X1 port map( A => n14610, Z => n21403);
   U13181 : BUF_X1 port map( A => n14610, Z => n21404);
   U13182 : BUF_X1 port map( A => n14610, Z => n21405);
   U13183 : BUF_X1 port map( A => n14610, Z => n21406);
   U13184 : BUF_X1 port map( A => n14543, Z => n21415);
   U13185 : BUF_X1 port map( A => n14543, Z => n21416);
   U13186 : BUF_X1 port map( A => n14543, Z => n21417);
   U13187 : BUF_X1 port map( A => n14543, Z => n21418);
   U13188 : BUF_X1 port map( A => n14543, Z => n21419);
   U13189 : BUF_X1 port map( A => n14477, Z => n21428);
   U13190 : BUF_X1 port map( A => n14477, Z => n21429);
   U13191 : BUF_X1 port map( A => n14477, Z => n21430);
   U13192 : BUF_X1 port map( A => n14477, Z => n21431);
   U13193 : BUF_X1 port map( A => n14477, Z => n21432);
   U13194 : BUF_X1 port map( A => n14407, Z => n21441);
   U13195 : BUF_X1 port map( A => n14407, Z => n21442);
   U13196 : BUF_X1 port map( A => n14407, Z => n21443);
   U13197 : BUF_X1 port map( A => n14407, Z => n21444);
   U13198 : BUF_X1 port map( A => n14407, Z => n21445);
   U13199 : BUF_X1 port map( A => n14341, Z => n21454);
   U13200 : BUF_X1 port map( A => n14341, Z => n21455);
   U13201 : BUF_X1 port map( A => n14341, Z => n21456);
   U13202 : BUF_X1 port map( A => n14341, Z => n21457);
   U13203 : BUF_X1 port map( A => n14341, Z => n21458);
   U13204 : BUF_X1 port map( A => n14274, Z => n21467);
   U13205 : BUF_X1 port map( A => n14274, Z => n21468);
   U13206 : BUF_X1 port map( A => n14274, Z => n21469);
   U13207 : BUF_X1 port map( A => n14274, Z => n21470);
   U13208 : BUF_X1 port map( A => n14274, Z => n21471);
   U13209 : BUF_X1 port map( A => n14208, Z => n21480);
   U13210 : BUF_X1 port map( A => n14208, Z => n21481);
   U13211 : BUF_X1 port map( A => n14208, Z => n21482);
   U13212 : BUF_X1 port map( A => n14208, Z => n21483);
   U13213 : BUF_X1 port map( A => n14208, Z => n21484);
   U13214 : BUF_X1 port map( A => n14141, Z => n21493);
   U13215 : BUF_X1 port map( A => n14141, Z => n21494);
   U13216 : BUF_X1 port map( A => n14141, Z => n21495);
   U13217 : BUF_X1 port map( A => n14141, Z => n21496);
   U13218 : BUF_X1 port map( A => n14141, Z => n21497);
   U13219 : BUF_X1 port map( A => n14074, Z => n21506);
   U13220 : BUF_X1 port map( A => n14074, Z => n21507);
   U13221 : BUF_X1 port map( A => n14074, Z => n21508);
   U13222 : BUF_X1 port map( A => n14074, Z => n21509);
   U13223 : BUF_X1 port map( A => n14074, Z => n21510);
   U13224 : BUF_X1 port map( A => n13941, Z => n21718);
   U13225 : BUF_X1 port map( A => n17350, Z => n20881);
   U13226 : BUF_X1 port map( A => n17350, Z => n20882);
   U13227 : BUF_X1 port map( A => n17350, Z => n20883);
   U13228 : BUF_X1 port map( A => n17350, Z => n20884);
   U13229 : BUF_X1 port map( A => n21080, Z => n21084);
   U13230 : BUF_X1 port map( A => n21079, Z => n21083);
   U13231 : BUF_X1 port map( A => n21079, Z => n21082);
   U13232 : BUF_X1 port map( A => n20982, Z => n20984);
   U13233 : BUF_X1 port map( A => n21122, Z => n21124);
   U13234 : BUF_X1 port map( A => n21135, Z => n21137);
   U13235 : BUF_X1 port map( A => n21148, Z => n21150);
   U13236 : BUF_X1 port map( A => n21161, Z => n21163);
   U13237 : BUF_X1 port map( A => n21174, Z => n21176);
   U13238 : BUF_X1 port map( A => n21187, Z => n21189);
   U13239 : BUF_X1 port map( A => n21200, Z => n21202);
   U13240 : BUF_X1 port map( A => n21213, Z => n21215);
   U13241 : BUF_X1 port map( A => n21226, Z => n21228);
   U13242 : BUF_X1 port map( A => n21239, Z => n21241);
   U13243 : BUF_X1 port map( A => n21252, Z => n21254);
   U13244 : BUF_X1 port map( A => n21265, Z => n21267);
   U13245 : BUF_X1 port map( A => n21278, Z => n21280);
   U13246 : BUF_X1 port map( A => n21291, Z => n21293);
   U13247 : BUF_X1 port map( A => n21304, Z => n21306);
   U13248 : BUF_X1 port map( A => n21330, Z => n21332);
   U13249 : BUF_X1 port map( A => n21343, Z => n21345);
   U13250 : BUF_X1 port map( A => n21356, Z => n21358);
   U13251 : BUF_X1 port map( A => n21369, Z => n21371);
   U13252 : BUF_X1 port map( A => n21382, Z => n21384);
   U13253 : BUF_X1 port map( A => n21395, Z => n21397);
   U13254 : BUF_X1 port map( A => n21408, Z => n21410);
   U13255 : BUF_X1 port map( A => n21421, Z => n21423);
   U13256 : BUF_X1 port map( A => n21434, Z => n21436);
   U13257 : BUF_X1 port map( A => n21447, Z => n21449);
   U13258 : BUF_X1 port map( A => n21460, Z => n21462);
   U13259 : BUF_X1 port map( A => n21473, Z => n21475);
   U13260 : BUF_X1 port map( A => n21486, Z => n21488);
   U13261 : BUF_X1 port map( A => n21499, Z => n21501);
   U13262 : BUF_X1 port map( A => n21512, Z => n21514);
   U13263 : BUF_X1 port map( A => n16084, Z => n21086);
   U13264 : BUF_X1 port map( A => n16084, Z => n21087);
   U13265 : BUF_X1 port map( A => n16084, Z => n21088);
   U13266 : BUF_X1 port map( A => n16084, Z => n21089);
   U13267 : BUF_X1 port map( A => n16084, Z => n21090);
   U13268 : BUF_X1 port map( A => n21122, Z => n21125);
   U13269 : BUF_X1 port map( A => n21122, Z => n21126);
   U13270 : BUF_X1 port map( A => n21123, Z => n21127);
   U13271 : BUF_X1 port map( A => n21123, Z => n21128);
   U13272 : BUF_X1 port map( A => n21135, Z => n21138);
   U13273 : BUF_X1 port map( A => n21135, Z => n21139);
   U13274 : BUF_X1 port map( A => n21136, Z => n21140);
   U13275 : BUF_X1 port map( A => n21136, Z => n21141);
   U13276 : BUF_X1 port map( A => n21148, Z => n21151);
   U13277 : BUF_X1 port map( A => n21148, Z => n21152);
   U13278 : BUF_X1 port map( A => n21149, Z => n21153);
   U13279 : BUF_X1 port map( A => n21149, Z => n21154);
   U13280 : BUF_X1 port map( A => n21161, Z => n21164);
   U13281 : BUF_X1 port map( A => n21161, Z => n21165);
   U13282 : BUF_X1 port map( A => n21162, Z => n21166);
   U13283 : BUF_X1 port map( A => n21162, Z => n21167);
   U13284 : BUF_X1 port map( A => n21174, Z => n21177);
   U13285 : BUF_X1 port map( A => n21174, Z => n21178);
   U13286 : BUF_X1 port map( A => n21175, Z => n21179);
   U13287 : BUF_X1 port map( A => n21175, Z => n21180);
   U13288 : BUF_X1 port map( A => n21187, Z => n21190);
   U13289 : BUF_X1 port map( A => n21187, Z => n21191);
   U13290 : BUF_X1 port map( A => n21188, Z => n21192);
   U13291 : BUF_X1 port map( A => n21188, Z => n21193);
   U13292 : BUF_X1 port map( A => n21200, Z => n21203);
   U13293 : BUF_X1 port map( A => n21200, Z => n21204);
   U13294 : BUF_X1 port map( A => n21201, Z => n21205);
   U13295 : BUF_X1 port map( A => n21201, Z => n21206);
   U13296 : BUF_X1 port map( A => n21213, Z => n21216);
   U13297 : BUF_X1 port map( A => n21213, Z => n21217);
   U13298 : BUF_X1 port map( A => n21214, Z => n21218);
   U13299 : BUF_X1 port map( A => n21214, Z => n21219);
   U13300 : BUF_X1 port map( A => n21226, Z => n21229);
   U13301 : BUF_X1 port map( A => n21226, Z => n21230);
   U13302 : BUF_X1 port map( A => n21227, Z => n21231);
   U13303 : BUF_X1 port map( A => n21227, Z => n21232);
   U13304 : BUF_X1 port map( A => n21239, Z => n21242);
   U13305 : BUF_X1 port map( A => n21239, Z => n21243);
   U13306 : BUF_X1 port map( A => n21240, Z => n21244);
   U13307 : BUF_X1 port map( A => n21240, Z => n21245);
   U13308 : BUF_X1 port map( A => n21252, Z => n21255);
   U13309 : BUF_X1 port map( A => n21252, Z => n21256);
   U13310 : BUF_X1 port map( A => n21253, Z => n21257);
   U13311 : BUF_X1 port map( A => n21253, Z => n21258);
   U13312 : BUF_X1 port map( A => n21265, Z => n21268);
   U13313 : BUF_X1 port map( A => n21265, Z => n21269);
   U13314 : BUF_X1 port map( A => n21266, Z => n21270);
   U13315 : BUF_X1 port map( A => n21266, Z => n21271);
   U13316 : BUF_X1 port map( A => n21278, Z => n21281);
   U13317 : BUF_X1 port map( A => n21278, Z => n21282);
   U13318 : BUF_X1 port map( A => n21279, Z => n21283);
   U13319 : BUF_X1 port map( A => n21279, Z => n21284);
   U13320 : BUF_X1 port map( A => n21291, Z => n21294);
   U13321 : BUF_X1 port map( A => n21291, Z => n21295);
   U13322 : BUF_X1 port map( A => n21292, Z => n21296);
   U13323 : BUF_X1 port map( A => n21292, Z => n21297);
   U13324 : BUF_X1 port map( A => n21304, Z => n21307);
   U13325 : BUF_X1 port map( A => n21304, Z => n21308);
   U13326 : BUF_X1 port map( A => n21305, Z => n21309);
   U13327 : BUF_X1 port map( A => n21305, Z => n21310);
   U13328 : BUF_X1 port map( A => n21330, Z => n21333);
   U13329 : BUF_X1 port map( A => n21330, Z => n21334);
   U13330 : BUF_X1 port map( A => n21331, Z => n21335);
   U13331 : BUF_X1 port map( A => n21331, Z => n21336);
   U13332 : BUF_X1 port map( A => n21343, Z => n21346);
   U13333 : BUF_X1 port map( A => n21343, Z => n21347);
   U13334 : BUF_X1 port map( A => n21344, Z => n21348);
   U13335 : BUF_X1 port map( A => n21344, Z => n21349);
   U13336 : BUF_X1 port map( A => n21356, Z => n21359);
   U13337 : BUF_X1 port map( A => n21356, Z => n21360);
   U13338 : BUF_X1 port map( A => n21357, Z => n21361);
   U13339 : BUF_X1 port map( A => n21357, Z => n21362);
   U13340 : BUF_X1 port map( A => n21369, Z => n21372);
   U13341 : BUF_X1 port map( A => n21369, Z => n21373);
   U13342 : BUF_X1 port map( A => n21370, Z => n21374);
   U13343 : BUF_X1 port map( A => n21370, Z => n21375);
   U13344 : BUF_X1 port map( A => n21382, Z => n21385);
   U13345 : BUF_X1 port map( A => n21382, Z => n21386);
   U13346 : BUF_X1 port map( A => n21383, Z => n21387);
   U13347 : BUF_X1 port map( A => n21383, Z => n21388);
   U13348 : BUF_X1 port map( A => n21395, Z => n21398);
   U13349 : BUF_X1 port map( A => n21395, Z => n21399);
   U13350 : BUF_X1 port map( A => n21396, Z => n21400);
   U13351 : BUF_X1 port map( A => n21396, Z => n21401);
   U13352 : BUF_X1 port map( A => n21408, Z => n21411);
   U13353 : BUF_X1 port map( A => n21408, Z => n21412);
   U13354 : BUF_X1 port map( A => n21409, Z => n21413);
   U13355 : BUF_X1 port map( A => n21409, Z => n21414);
   U13356 : BUF_X1 port map( A => n21421, Z => n21424);
   U13357 : BUF_X1 port map( A => n21421, Z => n21425);
   U13358 : BUF_X1 port map( A => n21422, Z => n21426);
   U13359 : BUF_X1 port map( A => n21422, Z => n21427);
   U13360 : BUF_X1 port map( A => n21434, Z => n21437);
   U13361 : BUF_X1 port map( A => n21434, Z => n21438);
   U13362 : BUF_X1 port map( A => n21435, Z => n21439);
   U13363 : BUF_X1 port map( A => n21435, Z => n21440);
   U13364 : BUF_X1 port map( A => n21447, Z => n21450);
   U13365 : BUF_X1 port map( A => n21447, Z => n21451);
   U13366 : BUF_X1 port map( A => n21448, Z => n21452);
   U13367 : BUF_X1 port map( A => n21448, Z => n21453);
   U13368 : BUF_X1 port map( A => n21460, Z => n21463);
   U13369 : BUF_X1 port map( A => n21460, Z => n21464);
   U13370 : BUF_X1 port map( A => n21461, Z => n21465);
   U13371 : BUF_X1 port map( A => n21461, Z => n21466);
   U13372 : BUF_X1 port map( A => n21473, Z => n21476);
   U13373 : BUF_X1 port map( A => n21473, Z => n21477);
   U13374 : BUF_X1 port map( A => n21474, Z => n21478);
   U13375 : BUF_X1 port map( A => n21474, Z => n21479);
   U13376 : BUF_X1 port map( A => n21486, Z => n21489);
   U13377 : BUF_X1 port map( A => n21486, Z => n21490);
   U13378 : BUF_X1 port map( A => n21487, Z => n21491);
   U13379 : BUF_X1 port map( A => n21487, Z => n21492);
   U13380 : BUF_X1 port map( A => n21499, Z => n21502);
   U13381 : BUF_X1 port map( A => n21499, Z => n21503);
   U13382 : BUF_X1 port map( A => n21500, Z => n21504);
   U13383 : BUF_X1 port map( A => n21500, Z => n21505);
   U13384 : BUF_X1 port map( A => n21512, Z => n21515);
   U13385 : BUF_X1 port map( A => n21512, Z => n21516);
   U13386 : BUF_X1 port map( A => n21513, Z => n21517);
   U13387 : BUF_X1 port map( A => n21513, Z => n21518);
   U13388 : BUF_X1 port map( A => n21079, Z => n21081);
   U13389 : BUF_X1 port map( A => n20982, Z => n20988);
   U13390 : BUF_X1 port map( A => n20982, Z => n20986);
   U13391 : BUF_X1 port map( A => n20982, Z => n20985);
   U13392 : BUF_X1 port map( A => n20982, Z => n20987);
   U13393 : BUF_X1 port map( A => n20982, Z => n20989);
   U13394 : BUF_X1 port map( A => n20983, Z => n20993);
   U13395 : BUF_X1 port map( A => n20983, Z => n20992);
   U13396 : BUF_X1 port map( A => n20983, Z => n20991);
   U13397 : BUF_X1 port map( A => n20983, Z => n20990);
   U13398 : NAND2_X1 port map( A1 => n21523, A2 => n21124, ZN => n16071);
   U13399 : NAND2_X1 port map( A1 => n21525, A2 => n21137, ZN => n16005);
   U13400 : NAND2_X1 port map( A1 => n21525, A2 => n21150, ZN => n15939);
   U13401 : NAND2_X1 port map( A1 => n21525, A2 => n21163, ZN => n15873);
   U13402 : NAND2_X1 port map( A1 => n21525, A2 => n21176, ZN => n15807);
   U13403 : NAND2_X1 port map( A1 => n21525, A2 => n21189, ZN => n15741);
   U13404 : NAND2_X1 port map( A1 => n21525, A2 => n21202, ZN => n15672);
   U13405 : NAND2_X1 port map( A1 => n21525, A2 => n21215, ZN => n15605);
   U13406 : NAND2_X1 port map( A1 => n21525, A2 => n21228, ZN => n15539);
   U13407 : NAND2_X1 port map( A1 => n21525, A2 => n21241, ZN => n15472);
   U13408 : NAND2_X1 port map( A1 => n21525, A2 => n21254, ZN => n15406);
   U13409 : NAND2_X1 port map( A1 => n21525, A2 => n21267, ZN => n15340);
   U13410 : NAND2_X1 port map( A1 => n21525, A2 => n21280, ZN => n15274);
   U13411 : NAND2_X1 port map( A1 => n21525, A2 => n21293, ZN => n15208);
   U13412 : NAND2_X1 port map( A1 => n21524, A2 => n21306, ZN => n15141);
   U13413 : NAND2_X1 port map( A1 => n21524, A2 => n21319, ZN => n15074);
   U13414 : NAND2_X1 port map( A1 => n21524, A2 => n21332, ZN => n15007);
   U13415 : NAND2_X1 port map( A1 => n21524, A2 => n21345, ZN => n14941);
   U13416 : NAND2_X1 port map( A1 => n21524, A2 => n21358, ZN => n14875);
   U13417 : NAND2_X1 port map( A1 => n21524, A2 => n21371, ZN => n14809);
   U13418 : NAND2_X1 port map( A1 => n21524, A2 => n21384, ZN => n14743);
   U13419 : NAND2_X1 port map( A1 => n21524, A2 => n21397, ZN => n14677);
   U13420 : NAND2_X1 port map( A1 => n21524, A2 => n21410, ZN => n14610);
   U13421 : NAND2_X1 port map( A1 => n21524, A2 => n21423, ZN => n14543);
   U13422 : NAND2_X1 port map( A1 => n21523, A2 => n21436, ZN => n14477);
   U13423 : NAND2_X1 port map( A1 => n21523, A2 => n21449, ZN => n14407);
   U13424 : NAND2_X1 port map( A1 => n21524, A2 => n21462, ZN => n14341);
   U13425 : NAND2_X1 port map( A1 => n21523, A2 => n21475, ZN => n14274);
   U13426 : NAND2_X1 port map( A1 => n21523, A2 => n21488, ZN => n14208);
   U13427 : NAND2_X1 port map( A1 => n21524, A2 => n21501, ZN => n14141);
   U13428 : NAND2_X1 port map( A1 => n21523, A2 => n21514, ZN => n14074);
   U13429 : BUF_X1 port map( A => n17350, Z => n20880);
   U13430 : BUF_X1 port map( A => n21080, Z => n21085);
   U13431 : NAND2_X1 port map( A1 => n21524, A2 => n21726, ZN => n13941);
   U13432 : BUF_X1 port map( A => n13939, Z => n21724);
   U13433 : BUF_X1 port map( A => n15072, Z => n21317);
   U13434 : BUF_X1 port map( A => n13939, Z => n21725);
   U13435 : BUF_X1 port map( A => n15072, Z => n21318);
   U13436 : BUF_X1 port map( A => n17363, Z => n20820);
   U13437 : BUF_X1 port map( A => n17363, Z => n20821);
   U13438 : BUF_X1 port map( A => n17363, Z => n20822);
   U13439 : BUF_X1 port map( A => n17363, Z => n20823);
   U13440 : BUF_X1 port map( A => n17363, Z => n20824);
   U13441 : BUF_X1 port map( A => n16097, Z => n21025);
   U13442 : BUF_X1 port map( A => n16097, Z => n21026);
   U13443 : BUF_X1 port map( A => n16097, Z => n21027);
   U13444 : BUF_X1 port map( A => n16097, Z => n21028);
   U13445 : BUF_X1 port map( A => n16097, Z => n21029);
   U13446 : BUF_X1 port map( A => n17348, Z => n20892);
   U13447 : BUF_X1 port map( A => n17377, Z => n20772);
   U13448 : BUF_X1 port map( A => n17348, Z => n20893);
   U13449 : BUF_X1 port map( A => n17377, Z => n20773);
   U13450 : BUF_X1 port map( A => n17348, Z => n20894);
   U13451 : BUF_X1 port map( A => n17377, Z => n20774);
   U13452 : BUF_X1 port map( A => n17348, Z => n20895);
   U13453 : BUF_X1 port map( A => n17377, Z => n20775);
   U13454 : BUF_X1 port map( A => n17348, Z => n20896);
   U13455 : BUF_X1 port map( A => n17377, Z => n20776);
   U13456 : BUF_X1 port map( A => n16081, Z => n21098);
   U13457 : BUF_X1 port map( A => n16081, Z => n21099);
   U13458 : BUF_X1 port map( A => n16081, Z => n21100);
   U13459 : BUF_X1 port map( A => n16081, Z => n21101);
   U13460 : BUF_X1 port map( A => n16081, Z => n21102);
   U13461 : BUF_X1 port map( A => n17373, Z => n20790);
   U13462 : BUF_X1 port map( A => n17387, Z => n20724);
   U13463 : BUF_X1 port map( A => n17373, Z => n20791);
   U13464 : BUF_X1 port map( A => n17387, Z => n20725);
   U13465 : BUF_X1 port map( A => n17373, Z => n20792);
   U13466 : BUF_X1 port map( A => n17387, Z => n20726);
   U13467 : BUF_X1 port map( A => n17373, Z => n20793);
   U13468 : BUF_X1 port map( A => n17387, Z => n20727);
   U13469 : BUF_X1 port map( A => n17373, Z => n20794);
   U13470 : BUF_X1 port map( A => n17387, Z => n20728);
   U13471 : BUF_X1 port map( A => n16112, Z => n20964);
   U13472 : BUF_X1 port map( A => n16107, Z => n20995);
   U13473 : BUF_X1 port map( A => n16122, Z => n20916);
   U13474 : BUF_X1 port map( A => n16107, Z => n20996);
   U13475 : BUF_X1 port map( A => n16112, Z => n20965);
   U13476 : BUF_X1 port map( A => n16122, Z => n20917);
   U13477 : BUF_X1 port map( A => n16107, Z => n20997);
   U13478 : BUF_X1 port map( A => n16112, Z => n20966);
   U13479 : BUF_X1 port map( A => n16122, Z => n20918);
   U13480 : BUF_X1 port map( A => n16107, Z => n20998);
   U13481 : BUF_X1 port map( A => n16112, Z => n20967);
   U13482 : BUF_X1 port map( A => n16122, Z => n20919);
   U13483 : BUF_X1 port map( A => n16107, Z => n20999);
   U13484 : BUF_X1 port map( A => n16112, Z => n20968);
   U13485 : BUF_X1 port map( A => n16122, Z => n20920);
   U13486 : BUF_X1 port map( A => n17353, Z => n20868);
   U13487 : BUF_X1 port map( A => n17358, Z => n20844);
   U13488 : BUF_X1 port map( A => n17382, Z => n20748);
   U13489 : BUF_X1 port map( A => n17353, Z => n20869);
   U13490 : BUF_X1 port map( A => n17358, Z => n20845);
   U13491 : BUF_X1 port map( A => n17382, Z => n20749);
   U13492 : BUF_X1 port map( A => n17353, Z => n20870);
   U13493 : BUF_X1 port map( A => n17358, Z => n20846);
   U13494 : BUF_X1 port map( A => n17382, Z => n20750);
   U13495 : BUF_X1 port map( A => n17353, Z => n20871);
   U13496 : BUF_X1 port map( A => n17358, Z => n20847);
   U13497 : BUF_X1 port map( A => n17382, Z => n20751);
   U13498 : BUF_X1 port map( A => n17353, Z => n20872);
   U13499 : BUF_X1 port map( A => n17358, Z => n20848);
   U13500 : BUF_X1 port map( A => n17382, Z => n20752);
   U13501 : BUF_X1 port map( A => n16092, Z => n21049);
   U13502 : BUF_X1 port map( A => n16117, Z => n20940);
   U13503 : BUF_X1 port map( A => n16092, Z => n21050);
   U13504 : BUF_X1 port map( A => n16117, Z => n20941);
   U13505 : BUF_X1 port map( A => n16092, Z => n21051);
   U13506 : BUF_X1 port map( A => n16117, Z => n20942);
   U13507 : BUF_X1 port map( A => n16092, Z => n21052);
   U13508 : BUF_X1 port map( A => n16117, Z => n20943);
   U13509 : BUF_X1 port map( A => n16092, Z => n21053);
   U13510 : BUF_X1 port map( A => n16117, Z => n20944);
   U13511 : BUF_X1 port map( A => n17360, Z => n20833);
   U13512 : BUF_X1 port map( A => n17345, Z => n20905);
   U13513 : BUF_X1 port map( A => n17355, Z => n20857);
   U13514 : BUF_X1 port map( A => n17370, Z => n20803);
   U13515 : BUF_X1 port map( A => n17360, Z => n20834);
   U13516 : BUF_X1 port map( A => n17345, Z => n20906);
   U13517 : BUF_X1 port map( A => n17355, Z => n20858);
   U13518 : BUF_X1 port map( A => n17370, Z => n20804);
   U13519 : BUF_X1 port map( A => n17360, Z => n20835);
   U13520 : BUF_X1 port map( A => n17345, Z => n20907);
   U13521 : BUF_X1 port map( A => n17355, Z => n20859);
   U13522 : BUF_X1 port map( A => n17370, Z => n20805);
   U13523 : BUF_X1 port map( A => n17360, Z => n20836);
   U13524 : BUF_X1 port map( A => n17345, Z => n20908);
   U13525 : BUF_X1 port map( A => n17355, Z => n20860);
   U13526 : BUF_X1 port map( A => n17370, Z => n20806);
   U13527 : BUF_X1 port map( A => n16087, Z => n21077);
   U13528 : BUF_X1 port map( A => n16094, Z => n21038);
   U13529 : BUF_X1 port map( A => n16078, Z => n21111);
   U13530 : BUF_X1 port map( A => n16089, Z => n21062);
   U13531 : BUF_X1 port map( A => n16104, Z => n21008);
   U13532 : BUF_X1 port map( A => n16087, Z => n21076);
   U13533 : BUF_X1 port map( A => n16094, Z => n21039);
   U13534 : BUF_X1 port map( A => n16078, Z => n21112);
   U13535 : BUF_X1 port map( A => n16089, Z => n21063);
   U13536 : BUF_X1 port map( A => n16104, Z => n21009);
   U13537 : BUF_X1 port map( A => n16087, Z => n21075);
   U13538 : BUF_X1 port map( A => n16094, Z => n21040);
   U13539 : BUF_X1 port map( A => n16078, Z => n21113);
   U13540 : BUF_X1 port map( A => n16089, Z => n21064);
   U13541 : BUF_X1 port map( A => n16104, Z => n21010);
   U13542 : BUF_X1 port map( A => n16087, Z => n21074);
   U13543 : BUF_X1 port map( A => n16094, Z => n21041);
   U13544 : BUF_X1 port map( A => n16078, Z => n21114);
   U13545 : BUF_X1 port map( A => n16089, Z => n21065);
   U13546 : BUF_X1 port map( A => n16104, Z => n21011);
   U13547 : BUF_X1 port map( A => n17379, Z => n20761);
   U13548 : BUF_X1 port map( A => n17374, Z => n20785);
   U13549 : BUF_X1 port map( A => n17384, Z => n20737);
   U13550 : BUF_X1 port map( A => n17379, Z => n20762);
   U13551 : BUF_X1 port map( A => n17374, Z => n20786);
   U13552 : BUF_X1 port map( A => n17384, Z => n20738);
   U13553 : BUF_X1 port map( A => n17379, Z => n20763);
   U13554 : BUF_X1 port map( A => n17374, Z => n20787);
   U13555 : BUF_X1 port map( A => n17384, Z => n20739);
   U13556 : BUF_X1 port map( A => n17379, Z => n20764);
   U13557 : BUF_X1 port map( A => n17374, Z => n20788);
   U13558 : BUF_X1 port map( A => n17384, Z => n20740);
   U13559 : BUF_X1 port map( A => n16114, Z => n20953);
   U13560 : BUF_X1 port map( A => n16109, Z => n20977);
   U13561 : BUF_X1 port map( A => n16119, Z => n20929);
   U13562 : BUF_X1 port map( A => n16114, Z => n20954);
   U13563 : BUF_X1 port map( A => n16109, Z => n20978);
   U13564 : BUF_X1 port map( A => n16119, Z => n20930);
   U13565 : BUF_X1 port map( A => n16114, Z => n20955);
   U13566 : BUF_X1 port map( A => n16109, Z => n20979);
   U13567 : BUF_X1 port map( A => n16119, Z => n20931);
   U13568 : BUF_X1 port map( A => n16114, Z => n20956);
   U13569 : BUF_X1 port map( A => n16109, Z => n20980);
   U13570 : BUF_X1 port map( A => n16119, Z => n20932);
   U13571 : BUF_X1 port map( A => n17364, Z => n20814);
   U13572 : BUF_X1 port map( A => n17364, Z => n20815);
   U13573 : BUF_X1 port map( A => n17364, Z => n20816);
   U13574 : BUF_X1 port map( A => n17364, Z => n20817);
   U13575 : BUF_X1 port map( A => n17364, Z => n20818);
   U13576 : BUF_X1 port map( A => n16098, Z => n21019);
   U13577 : BUF_X1 port map( A => n16098, Z => n21020);
   U13578 : BUF_X1 port map( A => n16098, Z => n21021);
   U13579 : BUF_X1 port map( A => n16098, Z => n21022);
   U13580 : BUF_X1 port map( A => n16098, Z => n21023);
   U13581 : BUF_X1 port map( A => n17349, Z => n20886);
   U13582 : BUF_X1 port map( A => n17349, Z => n20887);
   U13583 : BUF_X1 port map( A => n17349, Z => n20888);
   U13584 : BUF_X1 port map( A => n17349, Z => n20889);
   U13585 : BUF_X1 port map( A => n17349, Z => n20890);
   U13586 : BUF_X1 port map( A => n17378, Z => n20766);
   U13587 : BUF_X1 port map( A => n17388, Z => n20718);
   U13588 : BUF_X1 port map( A => n17378, Z => n20767);
   U13589 : BUF_X1 port map( A => n17388, Z => n20719);
   U13590 : BUF_X1 port map( A => n17378, Z => n20768);
   U13591 : BUF_X1 port map( A => n17388, Z => n20720);
   U13592 : BUF_X1 port map( A => n17378, Z => n20769);
   U13593 : BUF_X1 port map( A => n17388, Z => n20721);
   U13594 : BUF_X1 port map( A => n17378, Z => n20770);
   U13595 : BUF_X1 port map( A => n17388, Z => n20722);
   U13596 : BUF_X1 port map( A => n16082, Z => n21092);
   U13597 : BUF_X1 port map( A => n16113, Z => n20958);
   U13598 : BUF_X1 port map( A => n16123, Z => n20910);
   U13599 : BUF_X1 port map( A => n16082, Z => n21093);
   U13600 : BUF_X1 port map( A => n16113, Z => n20959);
   U13601 : BUF_X1 port map( A => n16123, Z => n20911);
   U13602 : BUF_X1 port map( A => n16082, Z => n21094);
   U13603 : BUF_X1 port map( A => n16113, Z => n20960);
   U13604 : BUF_X1 port map( A => n16123, Z => n20912);
   U13605 : BUF_X1 port map( A => n16082, Z => n21095);
   U13606 : BUF_X1 port map( A => n16113, Z => n20961);
   U13607 : BUF_X1 port map( A => n16123, Z => n20913);
   U13608 : BUF_X1 port map( A => n16082, Z => n21096);
   U13609 : BUF_X1 port map( A => n16113, Z => n20962);
   U13610 : BUF_X1 port map( A => n16123, Z => n20914);
   U13611 : BUF_X1 port map( A => n17354, Z => n20862);
   U13612 : BUF_X1 port map( A => n17383, Z => n20742);
   U13613 : BUF_X1 port map( A => n17354, Z => n20863);
   U13614 : BUF_X1 port map( A => n17383, Z => n20743);
   U13615 : BUF_X1 port map( A => n17354, Z => n20864);
   U13616 : BUF_X1 port map( A => n17383, Z => n20744);
   U13617 : BUF_X1 port map( A => n17354, Z => n20865);
   U13618 : BUF_X1 port map( A => n17383, Z => n20745);
   U13619 : BUF_X1 port map( A => n17354, Z => n20866);
   U13620 : BUF_X1 port map( A => n17383, Z => n20746);
   U13621 : BUF_X1 port map( A => n17359, Z => n20838);
   U13622 : BUF_X1 port map( A => n17359, Z => n20839);
   U13623 : BUF_X1 port map( A => n17359, Z => n20840);
   U13624 : BUF_X1 port map( A => n17359, Z => n20841);
   U13625 : BUF_X1 port map( A => n17359, Z => n20842);
   U13626 : BUF_X1 port map( A => n16093, Z => n21043);
   U13627 : BUF_X1 port map( A => n16118, Z => n20934);
   U13628 : BUF_X1 port map( A => n16093, Z => n21044);
   U13629 : BUF_X1 port map( A => n16118, Z => n20935);
   U13630 : BUF_X1 port map( A => n16093, Z => n21045);
   U13631 : BUF_X1 port map( A => n16118, Z => n20936);
   U13632 : BUF_X1 port map( A => n16093, Z => n21046);
   U13633 : BUF_X1 port map( A => n16118, Z => n20937);
   U13634 : BUF_X1 port map( A => n16093, Z => n21047);
   U13635 : BUF_X1 port map( A => n16118, Z => n20938);
   U13636 : BUF_X1 port map( A => n17365, Z => n20808);
   U13637 : BUF_X1 port map( A => n17365, Z => n20809);
   U13638 : BUF_X1 port map( A => n17365, Z => n20810);
   U13639 : BUF_X1 port map( A => n17365, Z => n20811);
   U13640 : BUF_X1 port map( A => n17365, Z => n20812);
   U13641 : BUF_X1 port map( A => n16099, Z => n21013);
   U13642 : BUF_X1 port map( A => n16099, Z => n21014);
   U13643 : BUF_X1 port map( A => n16099, Z => n21015);
   U13644 : BUF_X1 port map( A => n16099, Z => n21016);
   U13645 : BUF_X1 port map( A => n16099, Z => n21017);
   U13646 : NAND2_X1 port map( A1 => n18512, A2 => n18515, ZN => n17350);
   U13647 : BUF_X1 port map( A => n21519, Z => n21521);
   U13648 : BUF_X1 port map( A => n21519, Z => n21522);
   U13649 : BUF_X1 port map( A => n21519, Z => n21523);
   U13650 : BUF_X1 port map( A => n21520, Z => n21525);
   U13651 : BUF_X1 port map( A => n21520, Z => n21524);
   U13652 : BUF_X1 port map( A => n17361, Z => n20826);
   U13653 : BUF_X1 port map( A => n17346, Z => n20898);
   U13654 : BUF_X1 port map( A => n17351, Z => n20874);
   U13655 : BUF_X1 port map( A => n17371, Z => n20796);
   U13656 : BUF_X1 port map( A => n17385, Z => n20730);
   U13657 : BUF_X1 port map( A => n17361, Z => n20827);
   U13658 : BUF_X1 port map( A => n17346, Z => n20899);
   U13659 : BUF_X1 port map( A => n17351, Z => n20875);
   U13660 : BUF_X1 port map( A => n17371, Z => n20797);
   U13661 : BUF_X1 port map( A => n17385, Z => n20731);
   U13662 : BUF_X1 port map( A => n17361, Z => n20828);
   U13663 : BUF_X1 port map( A => n17346, Z => n20900);
   U13664 : BUF_X1 port map( A => n17351, Z => n20876);
   U13665 : BUF_X1 port map( A => n17371, Z => n20798);
   U13666 : BUF_X1 port map( A => n17385, Z => n20732);
   U13667 : BUF_X1 port map( A => n17361, Z => n20829);
   U13668 : BUF_X1 port map( A => n17346, Z => n20901);
   U13669 : BUF_X1 port map( A => n17351, Z => n20877);
   U13670 : BUF_X1 port map( A => n17371, Z => n20799);
   U13671 : BUF_X1 port map( A => n17385, Z => n20733);
   U13672 : BUF_X1 port map( A => n17361, Z => n20830);
   U13673 : BUF_X1 port map( A => n17346, Z => n20902);
   U13674 : BUF_X1 port map( A => n17351, Z => n20878);
   U13675 : BUF_X1 port map( A => n17371, Z => n20800);
   U13676 : BUF_X1 port map( A => n17385, Z => n20734);
   U13677 : BUF_X1 port map( A => n16088, Z => n21067);
   U13678 : BUF_X1 port map( A => n16095, Z => n21031);
   U13679 : BUF_X1 port map( A => n16079, Z => n21104);
   U13680 : BUF_X1 port map( A => n16105, Z => n21001);
   U13681 : BUF_X1 port map( A => n16120, Z => n20922);
   U13682 : BUF_X1 port map( A => n16088, Z => n21068);
   U13683 : BUF_X1 port map( A => n16095, Z => n21032);
   U13684 : BUF_X1 port map( A => n16079, Z => n21105);
   U13685 : BUF_X1 port map( A => n16105, Z => n21002);
   U13686 : BUF_X1 port map( A => n16120, Z => n20923);
   U13687 : BUF_X1 port map( A => n16088, Z => n21069);
   U13688 : BUF_X1 port map( A => n16095, Z => n21033);
   U13689 : BUF_X1 port map( A => n16079, Z => n21106);
   U13690 : BUF_X1 port map( A => n16105, Z => n21003);
   U13691 : BUF_X1 port map( A => n16120, Z => n20924);
   U13692 : BUF_X1 port map( A => n16088, Z => n21070);
   U13693 : BUF_X1 port map( A => n16095, Z => n21034);
   U13694 : BUF_X1 port map( A => n16079, Z => n21107);
   U13695 : BUF_X1 port map( A => n16105, Z => n21004);
   U13696 : BUF_X1 port map( A => n16120, Z => n20925);
   U13697 : BUF_X1 port map( A => n16088, Z => n21071);
   U13698 : BUF_X1 port map( A => n16095, Z => n21035);
   U13699 : BUF_X1 port map( A => n16079, Z => n21108);
   U13700 : BUF_X1 port map( A => n16105, Z => n21005);
   U13701 : BUF_X1 port map( A => n16120, Z => n20926);
   U13702 : BUF_X1 port map( A => n17356, Z => n20850);
   U13703 : BUF_X1 port map( A => n17380, Z => n20754);
   U13704 : BUF_X1 port map( A => n17375, Z => n20778);
   U13705 : BUF_X1 port map( A => n17356, Z => n20851);
   U13706 : BUF_X1 port map( A => n17380, Z => n20755);
   U13707 : BUF_X1 port map( A => n17375, Z => n20779);
   U13708 : BUF_X1 port map( A => n17356, Z => n20852);
   U13709 : BUF_X1 port map( A => n17380, Z => n20756);
   U13710 : BUF_X1 port map( A => n17375, Z => n20780);
   U13711 : BUF_X1 port map( A => n17356, Z => n20853);
   U13712 : BUF_X1 port map( A => n17380, Z => n20757);
   U13713 : BUF_X1 port map( A => n17375, Z => n20781);
   U13714 : BUF_X1 port map( A => n17356, Z => n20854);
   U13715 : BUF_X1 port map( A => n17380, Z => n20758);
   U13716 : BUF_X1 port map( A => n17375, Z => n20782);
   U13717 : BUF_X1 port map( A => n16090, Z => n21055);
   U13718 : BUF_X1 port map( A => n16115, Z => n20946);
   U13719 : BUF_X1 port map( A => n16110, Z => n20970);
   U13720 : BUF_X1 port map( A => n16090, Z => n21056);
   U13721 : BUF_X1 port map( A => n16115, Z => n20947);
   U13722 : BUF_X1 port map( A => n16110, Z => n20971);
   U13723 : BUF_X1 port map( A => n16090, Z => n21057);
   U13724 : BUF_X1 port map( A => n16115, Z => n20948);
   U13725 : BUF_X1 port map( A => n16110, Z => n20972);
   U13726 : BUF_X1 port map( A => n16090, Z => n21058);
   U13727 : BUF_X1 port map( A => n16115, Z => n20949);
   U13728 : BUF_X1 port map( A => n16110, Z => n20973);
   U13729 : BUF_X1 port map( A => n16090, Z => n21059);
   U13730 : BUF_X1 port map( A => n16115, Z => n20950);
   U13731 : BUF_X1 port map( A => n16110, Z => n20974);
   U13732 : AND2_X1 port map( A1 => n17311, A2 => n17314, ZN => n16084);
   U13733 : BUF_X1 port map( A => n16087, Z => n21073);
   U13734 : BUF_X1 port map( A => n17345, Z => n20904);
   U13735 : BUF_X1 port map( A => n17355, Z => n20856);
   U13736 : BUF_X1 port map( A => n17370, Z => n20802);
   U13737 : BUF_X1 port map( A => n16094, Z => n21037);
   U13738 : BUF_X1 port map( A => n16078, Z => n21110);
   U13739 : BUF_X1 port map( A => n16089, Z => n21061);
   U13740 : BUF_X1 port map( A => n17360, Z => n20832);
   U13741 : BUF_X1 port map( A => n16104, Z => n21007);
   U13742 : BUF_X1 port map( A => n17379, Z => n20760);
   U13743 : BUF_X1 port map( A => n17374, Z => n20784);
   U13744 : BUF_X1 port map( A => n17384, Z => n20736);
   U13745 : BUF_X1 port map( A => n16114, Z => n20952);
   U13746 : BUF_X1 port map( A => n16109, Z => n20976);
   U13747 : BUF_X1 port map( A => n16119, Z => n20928);
   U13748 : OAI21_X1 port map( B1 => n14070, B2 => n14071, A => n21521, ZN => 
                           n13939);
   U13749 : OAI21_X1 port map( B1 => n14071, B2 => n15138, A => n21522, ZN => 
                           n15072);
   U13750 : BUF_X1 port map( A => n16108, Z => n20982);
   U13751 : BUF_X1 port map( A => n16108, Z => n20983);
   U13752 : BUF_X1 port map( A => n14475, Z => n21434);
   U13753 : BUF_X1 port map( A => n14339, Z => n21460);
   U13754 : BUF_X1 port map( A => n14206, Z => n21486);
   U13755 : BUF_X1 port map( A => n14405, Z => n21447);
   U13756 : BUF_X1 port map( A => n14272, Z => n21473);
   U13757 : BUF_X1 port map( A => n14139, Z => n21499);
   U13758 : BUF_X1 port map( A => n16069, Z => n21122);
   U13759 : BUF_X1 port map( A => n16003, Z => n21135);
   U13760 : BUF_X1 port map( A => n15937, Z => n21148);
   U13761 : BUF_X1 port map( A => n15871, Z => n21161);
   U13762 : BUF_X1 port map( A => n15805, Z => n21174);
   U13763 : BUF_X1 port map( A => n15739, Z => n21187);
   U13764 : BUF_X1 port map( A => n15670, Z => n21200);
   U13765 : BUF_X1 port map( A => n15603, Z => n21213);
   U13766 : BUF_X1 port map( A => n15537, Z => n21226);
   U13767 : BUF_X1 port map( A => n15470, Z => n21239);
   U13768 : BUF_X1 port map( A => n15404, Z => n21252);
   U13769 : BUF_X1 port map( A => n15338, Z => n21265);
   U13770 : BUF_X1 port map( A => n15272, Z => n21278);
   U13771 : BUF_X1 port map( A => n15206, Z => n21291);
   U13772 : BUF_X1 port map( A => n15139, Z => n21304);
   U13773 : BUF_X1 port map( A => n15005, Z => n21330);
   U13774 : BUF_X1 port map( A => n14939, Z => n21343);
   U13775 : BUF_X1 port map( A => n14873, Z => n21356);
   U13776 : BUF_X1 port map( A => n14807, Z => n21369);
   U13777 : BUF_X1 port map( A => n14741, Z => n21382);
   U13778 : BUF_X1 port map( A => n14675, Z => n21395);
   U13779 : BUF_X1 port map( A => n14608, Z => n21408);
   U13780 : BUF_X1 port map( A => n14541, Z => n21421);
   U13781 : BUF_X1 port map( A => n14072, Z => n21512);
   U13782 : BUF_X1 port map( A => n16085, Z => n21079);
   U13783 : BUF_X1 port map( A => n14475, Z => n21435);
   U13784 : BUF_X1 port map( A => n14339, Z => n21461);
   U13785 : BUF_X1 port map( A => n14206, Z => n21487);
   U13786 : BUF_X1 port map( A => n14405, Z => n21448);
   U13787 : BUF_X1 port map( A => n14272, Z => n21474);
   U13788 : BUF_X1 port map( A => n14139, Z => n21500);
   U13789 : BUF_X1 port map( A => n16069, Z => n21123);
   U13790 : BUF_X1 port map( A => n16003, Z => n21136);
   U13791 : BUF_X1 port map( A => n15937, Z => n21149);
   U13792 : BUF_X1 port map( A => n15871, Z => n21162);
   U13793 : BUF_X1 port map( A => n15805, Z => n21175);
   U13794 : BUF_X1 port map( A => n15739, Z => n21188);
   U13795 : BUF_X1 port map( A => n15670, Z => n21201);
   U13796 : BUF_X1 port map( A => n15603, Z => n21214);
   U13797 : BUF_X1 port map( A => n15537, Z => n21227);
   U13798 : BUF_X1 port map( A => n15470, Z => n21240);
   U13799 : BUF_X1 port map( A => n15404, Z => n21253);
   U13800 : BUF_X1 port map( A => n15338, Z => n21266);
   U13801 : BUF_X1 port map( A => n15272, Z => n21279);
   U13802 : BUF_X1 port map( A => n15206, Z => n21292);
   U13803 : BUF_X1 port map( A => n15139, Z => n21305);
   U13804 : BUF_X1 port map( A => n15005, Z => n21331);
   U13805 : BUF_X1 port map( A => n14939, Z => n21344);
   U13806 : BUF_X1 port map( A => n14873, Z => n21357);
   U13807 : BUF_X1 port map( A => n14807, Z => n21370);
   U13808 : BUF_X1 port map( A => n14741, Z => n21383);
   U13809 : BUF_X1 port map( A => n14675, Z => n21396);
   U13810 : BUF_X1 port map( A => n14608, Z => n21409);
   U13811 : BUF_X1 port map( A => n14541, Z => n21422);
   U13812 : BUF_X1 port map( A => n14072, Z => n21513);
   U13813 : BUF_X1 port map( A => n16085, Z => n21080);
   U13814 : NOR3_X1 port map( A1 => n17338, A2 => n20984, A3 => n17337, ZN => 
                           n17311);
   U13815 : NOR3_X1 port map( A1 => n18534, A2 => n18535, A3 => n18532, ZN => 
                           n18515);
   U13816 : NOR3_X1 port map( A1 => n17333, A2 => n17334, A3 => n17331, ZN => 
                           n17314);
   U13817 : NAND2_X1 port map( A1 => n17425, A2 => n17426, ZN => n5305);
   U13818 : NOR4_X1 port map( A1 => n17435, A2 => n17436, A3 => n17437, A4 => 
                           n17438, ZN => n17425);
   U13819 : NOR4_X1 port map( A1 => n17427, A2 => n17428, A3 => n17429, A4 => 
                           n17430, ZN => n17426);
   U13820 : OAI221_X1 port map( B1 => n14480, B2 => n20741, C1 => n15876, C2 =>
                           n20735, A => n17442, ZN => n17435);
   U13821 : NAND2_X1 port map( A1 => n17407, A2 => n17408, ZN => n5306);
   U13822 : NOR4_X1 port map( A1 => n17417, A2 => n17418, A3 => n17419, A4 => 
                           n17420, ZN => n17407);
   U13823 : NOR4_X1 port map( A1 => n17409, A2 => n17410, A3 => n17411, A4 => 
                           n17412, ZN => n17408);
   U13824 : OAI221_X1 port map( B1 => n14479, B2 => n20741, C1 => n15875, C2 =>
                           n20735, A => n17424, ZN => n17417);
   U13825 : NAND2_X1 port map( A1 => n17389, A2 => n17390, ZN => n5307);
   U13826 : NOR4_X1 port map( A1 => n17399, A2 => n17400, A3 => n17401, A4 => 
                           n17402, ZN => n17389);
   U13827 : NOR4_X1 port map( A1 => n17391, A2 => n17392, A3 => n17393, A4 => 
                           n17394, ZN => n17390);
   U13828 : OAI221_X1 port map( B1 => n14478, B2 => n20741, C1 => n15874, C2 =>
                           n20735, A => n17406, ZN => n17399);
   U13829 : NAND2_X1 port map( A1 => n17339, A2 => n17340, ZN => n5308);
   U13830 : NOR4_X1 port map( A1 => n17366, A2 => n17367, A3 => n17368, A4 => 
                           n17369, ZN => n17339);
   U13831 : NOR4_X1 port map( A1 => n17341, A2 => n17342, A3 => n17343, A4 => 
                           n17344, ZN => n17340);
   U13832 : OAI221_X1 port map( B1 => n14476, B2 => n20741, C1 => n15872, C2 =>
                           n20735, A => n17386, ZN => n17366);
   U13833 : NAND2_X1 port map( A1 => n17075, A2 => n17076, ZN => n5333);
   U13834 : NOR4_X1 port map( A1 => n17085, A2 => n17086, A3 => n17087, A4 => 
                           n17088, ZN => n17075);
   U13835 : NOR4_X1 port map( A1 => n17077, A2 => n17078, A3 => n17079, A4 => 
                           n17080, ZN => n17076);
   U13836 : OAI221_X1 port map( B1 => n14528, B2 => n20929, C1 => n15924, C2 =>
                           n20923, A => n17092, ZN => n17085);
   U13837 : NAND2_X1 port map( A1 => n17056, A2 => n17057, ZN => n5335);
   U13838 : NOR4_X1 port map( A1 => n17066, A2 => n17067, A3 => n17068, A4 => 
                           n17069, ZN => n17056);
   U13839 : NOR4_X1 port map( A1 => n17058, A2 => n17059, A3 => n17060, A4 => 
                           n17061, ZN => n17057);
   U13840 : OAI221_X1 port map( B1 => n14527, B2 => n20929, C1 => n15923, C2 =>
                           n20923, A => n17073, ZN => n17066);
   U13841 : NAND2_X1 port map( A1 => n17037, A2 => n17038, ZN => n5337);
   U13842 : NOR4_X1 port map( A1 => n17047, A2 => n17048, A3 => n17049, A4 => 
                           n17050, ZN => n17037);
   U13843 : NOR4_X1 port map( A1 => n17039, A2 => n17040, A3 => n17041, A4 => 
                           n17042, ZN => n17038);
   U13844 : OAI221_X1 port map( B1 => n14526, B2 => n20929, C1 => n15922, C2 =>
                           n20923, A => n17054, ZN => n17047);
   U13845 : NAND2_X1 port map( A1 => n17018, A2 => n17019, ZN => n5339);
   U13846 : NOR4_X1 port map( A1 => n17028, A2 => n17029, A3 => n17030, A4 => 
                           n17031, ZN => n17018);
   U13847 : NOR4_X1 port map( A1 => n17020, A2 => n17021, A3 => n17022, A4 => 
                           n17023, ZN => n17019);
   U13848 : OAI221_X1 port map( B1 => n14525, B2 => n20929, C1 => n15921, C2 =>
                           n20923, A => n17035, ZN => n17028);
   U13849 : NAND2_X1 port map( A1 => n16999, A2 => n17000, ZN => n5341);
   U13850 : NOR4_X1 port map( A1 => n17009, A2 => n17010, A3 => n17011, A4 => 
                           n17012, ZN => n16999);
   U13851 : NOR4_X1 port map( A1 => n17001, A2 => n17002, A3 => n17003, A4 => 
                           n17004, ZN => n17000);
   U13852 : OAI221_X1 port map( B1 => n14524, B2 => n20929, C1 => n15920, C2 =>
                           n20923, A => n17016, ZN => n17009);
   U13853 : NAND2_X1 port map( A1 => n16980, A2 => n16981, ZN => n5343);
   U13854 : NOR4_X1 port map( A1 => n16990, A2 => n16991, A3 => n16992, A4 => 
                           n16993, ZN => n16980);
   U13855 : NOR4_X1 port map( A1 => n16982, A2 => n16983, A3 => n16984, A4 => 
                           n16985, ZN => n16981);
   U13856 : OAI221_X1 port map( B1 => n14523, B2 => n20929, C1 => n15919, C2 =>
                           n20923, A => n16997, ZN => n16990);
   U13857 : NAND2_X1 port map( A1 => n16961, A2 => n16962, ZN => n5345);
   U13858 : NOR4_X1 port map( A1 => n16971, A2 => n16972, A3 => n16973, A4 => 
                           n16974, ZN => n16961);
   U13859 : NOR4_X1 port map( A1 => n16963, A2 => n16964, A3 => n16965, A4 => 
                           n16966, ZN => n16962);
   U13860 : OAI221_X1 port map( B1 => n14522, B2 => n20929, C1 => n15918, C2 =>
                           n20923, A => n16978, ZN => n16971);
   U13861 : NAND2_X1 port map( A1 => n16942, A2 => n16943, ZN => n5347);
   U13862 : NOR4_X1 port map( A1 => n16952, A2 => n16953, A3 => n16954, A4 => 
                           n16955, ZN => n16942);
   U13863 : NOR4_X1 port map( A1 => n16944, A2 => n16945, A3 => n16946, A4 => 
                           n16947, ZN => n16943);
   U13864 : OAI221_X1 port map( B1 => n14521, B2 => n20929, C1 => n15917, C2 =>
                           n20923, A => n16959, ZN => n16952);
   U13865 : NAND2_X1 port map( A1 => n16923, A2 => n16924, ZN => n5349);
   U13866 : NOR4_X1 port map( A1 => n16933, A2 => n16934, A3 => n16935, A4 => 
                           n16936, ZN => n16923);
   U13867 : NOR4_X1 port map( A1 => n16925, A2 => n16926, A3 => n16927, A4 => 
                           n16928, ZN => n16924);
   U13868 : OAI221_X1 port map( B1 => n14520, B2 => n20929, C1 => n15916, C2 =>
                           n20923, A => n16940, ZN => n16933);
   U13869 : NAND2_X1 port map( A1 => n16904, A2 => n16905, ZN => n5351);
   U13870 : NOR4_X1 port map( A1 => n16914, A2 => n16915, A3 => n16916, A4 => 
                           n16917, ZN => n16904);
   U13871 : NOR4_X1 port map( A1 => n16906, A2 => n16907, A3 => n16908, A4 => 
                           n16909, ZN => n16905);
   U13872 : OAI221_X1 port map( B1 => n14519, B2 => n20929, C1 => n15915, C2 =>
                           n20923, A => n16921, ZN => n16914);
   U13873 : NAND2_X1 port map( A1 => n16885, A2 => n16886, ZN => n5353);
   U13874 : NOR4_X1 port map( A1 => n16895, A2 => n16896, A3 => n16897, A4 => 
                           n16898, ZN => n16885);
   U13875 : NOR4_X1 port map( A1 => n16887, A2 => n16888, A3 => n16889, A4 => 
                           n16890, ZN => n16886);
   U13876 : OAI221_X1 port map( B1 => n14518, B2 => n20929, C1 => n15914, C2 =>
                           n20923, A => n16902, ZN => n16895);
   U13877 : NAND2_X1 port map( A1 => n16334, A2 => n16335, ZN => n5411);
   U13878 : NOR4_X1 port map( A1 => n16344, A2 => n16345, A3 => n16346, A4 => 
                           n16347, ZN => n16334);
   U13879 : NOR4_X1 port map( A1 => n16336, A2 => n16337, A3 => n16338, A4 => 
                           n16339, ZN => n16335);
   U13880 : OAI221_X1 port map( B1 => n14489, B2 => n20932, C1 => n15885, C2 =>
                           n20926, A => n16351, ZN => n16344);
   U13881 : NAND2_X1 port map( A1 => n18512, A2 => n18523, ZN => n17356);
   U13882 : NAND2_X1 port map( A1 => n15737, A2 => n15738, ZN => n14071);
   U13883 : NAND2_X1 port map( A1 => n17311, A2 => n17322, ZN => n16090);
   U13884 : NAND2_X1 port map( A1 => n18531, A2 => n18524, ZN => n17380);
   U13885 : NAND2_X1 port map( A1 => n18531, A2 => n18519, ZN => n17375);
   U13886 : NAND2_X1 port map( A1 => n17330, A2 => n17323, ZN => n16115);
   U13887 : NAND2_X1 port map( A1 => n17330, A2 => n17319, ZN => n16110);
   U13888 : NAND2_X1 port map( A1 => n18512, A2 => n18517, ZN => n17384);
   U13889 : NAND2_X1 port map( A1 => n18516, A2 => n18514, ZN => n17346);
   U13890 : NAND2_X1 port map( A1 => n18521, A2 => n18514, ZN => n17351);
   U13891 : NAND2_X1 port map( A1 => n18523, A2 => n18514, ZN => n17385);
   U13892 : NAND2_X1 port map( A1 => n17319, A2 => n17313, ZN => n16088);
   U13893 : NAND2_X1 port map( A1 => n17315, A2 => n17313, ZN => n16079);
   U13894 : NAND2_X1 port map( A1 => n17322, A2 => n17313, ZN => n16120);
   U13895 : NAND2_X1 port map( A1 => n17311, A2 => n17316, ZN => n16119);
   U13896 : NAND2_X1 port map( A1 => n18519, A2 => n18512, ZN => n17371);
   U13897 : NAND2_X1 port map( A1 => n18523, A2 => n18520, ZN => n17361);
   U13898 : NAND2_X1 port map( A1 => n17322, A2 => n17320, ZN => n16095);
   U13899 : NAND2_X1 port map( A1 => n18531, A2 => n18517, ZN => n17379);
   U13900 : NAND2_X1 port map( A1 => n18531, A2 => n18523, ZN => n17374);
   U13901 : NAND2_X1 port map( A1 => n17330, A2 => n17316, ZN => n16114);
   U13902 : NAND2_X1 port map( A1 => n17330, A2 => n17322, ZN => n16109);
   U13903 : NAND2_X1 port map( A1 => n17319, A2 => n17311, ZN => n16105);
   U13904 : BUF_X1 port map( A => n14068, Z => n21527);
   U13905 : BUF_X1 port map( A => n14066, Z => n21530);
   U13906 : BUF_X1 port map( A => n14064, Z => n21533);
   U13907 : BUF_X1 port map( A => n14062, Z => n21536);
   U13908 : BUF_X1 port map( A => n14060, Z => n21539);
   U13909 : BUF_X1 port map( A => n14058, Z => n21542);
   U13910 : BUF_X1 port map( A => n14056, Z => n21545);
   U13911 : BUF_X1 port map( A => n14054, Z => n21548);
   U13912 : BUF_X1 port map( A => n14052, Z => n21551);
   U13913 : BUF_X1 port map( A => n14050, Z => n21554);
   U13914 : BUF_X1 port map( A => n14048, Z => n21557);
   U13915 : BUF_X1 port map( A => n14046, Z => n21560);
   U13916 : BUF_X1 port map( A => n14044, Z => n21563);
   U13917 : BUF_X1 port map( A => n14042, Z => n21566);
   U13918 : BUF_X1 port map( A => n14040, Z => n21569);
   U13919 : BUF_X1 port map( A => n14038, Z => n21572);
   U13920 : BUF_X1 port map( A => n14036, Z => n21575);
   U13921 : BUF_X1 port map( A => n14034, Z => n21578);
   U13922 : BUF_X1 port map( A => n14032, Z => n21581);
   U13923 : BUF_X1 port map( A => n14030, Z => n21584);
   U13924 : BUF_X1 port map( A => n14028, Z => n21587);
   U13925 : BUF_X1 port map( A => n14026, Z => n21590);
   U13926 : BUF_X1 port map( A => n14024, Z => n21593);
   U13927 : BUF_X1 port map( A => n14022, Z => n21596);
   U13928 : BUF_X1 port map( A => n14020, Z => n21599);
   U13929 : BUF_X1 port map( A => n14018, Z => n21602);
   U13930 : BUF_X1 port map( A => n14016, Z => n21605);
   U13931 : BUF_X1 port map( A => n14014, Z => n21608);
   U13932 : BUF_X1 port map( A => n14012, Z => n21611);
   U13933 : BUF_X1 port map( A => n14010, Z => n21614);
   U13934 : BUF_X1 port map( A => n14008, Z => n21617);
   U13935 : BUF_X1 port map( A => n14006, Z => n21620);
   U13936 : BUF_X1 port map( A => n14004, Z => n21623);
   U13937 : BUF_X1 port map( A => n14002, Z => n21626);
   U13938 : BUF_X1 port map( A => n14000, Z => n21629);
   U13939 : BUF_X1 port map( A => n13998, Z => n21632);
   U13940 : BUF_X1 port map( A => n13996, Z => n21635);
   U13941 : BUF_X1 port map( A => n13994, Z => n21638);
   U13942 : BUF_X1 port map( A => n13992, Z => n21641);
   U13943 : BUF_X1 port map( A => n13990, Z => n21644);
   U13944 : BUF_X1 port map( A => n13988, Z => n21647);
   U13945 : BUF_X1 port map( A => n13986, Z => n21650);
   U13946 : BUF_X1 port map( A => n13984, Z => n21653);
   U13947 : BUF_X1 port map( A => n13982, Z => n21656);
   U13948 : BUF_X1 port map( A => n13980, Z => n21659);
   U13949 : BUF_X1 port map( A => n13978, Z => n21662);
   U13950 : BUF_X1 port map( A => n13976, Z => n21665);
   U13951 : BUF_X1 port map( A => n13974, Z => n21668);
   U13952 : BUF_X1 port map( A => n13972, Z => n21671);
   U13953 : BUF_X1 port map( A => n13970, Z => n21674);
   U13954 : BUF_X1 port map( A => n13968, Z => n21677);
   U13955 : BUF_X1 port map( A => n13966, Z => n21680);
   U13956 : BUF_X1 port map( A => n13964, Z => n21683);
   U13957 : BUF_X1 port map( A => n13962, Z => n21686);
   U13958 : BUF_X1 port map( A => n13960, Z => n21689);
   U13959 : BUF_X1 port map( A => n13958, Z => n21692);
   U13960 : BUF_X1 port map( A => n13956, Z => n21695);
   U13961 : BUF_X1 port map( A => n13954, Z => n21698);
   U13962 : BUF_X1 port map( A => n13952, Z => n21701);
   U13963 : BUF_X1 port map( A => n13950, Z => n21704);
   U13964 : BUF_X1 port map( A => n13948, Z => n21707);
   U13965 : BUF_X1 port map( A => n13946, Z => n21710);
   U13966 : BUF_X1 port map( A => n13944, Z => n21713);
   U13967 : BUF_X1 port map( A => n13942, Z => n21716);
   U13968 : BUF_X1 port map( A => n14068, Z => n21526);
   U13969 : BUF_X1 port map( A => n14066, Z => n21529);
   U13970 : BUF_X1 port map( A => n14064, Z => n21532);
   U13971 : BUF_X1 port map( A => n14062, Z => n21535);
   U13972 : BUF_X1 port map( A => n14060, Z => n21538);
   U13973 : BUF_X1 port map( A => n14058, Z => n21541);
   U13974 : BUF_X1 port map( A => n14056, Z => n21544);
   U13975 : BUF_X1 port map( A => n14054, Z => n21547);
   U13976 : BUF_X1 port map( A => n14052, Z => n21550);
   U13977 : BUF_X1 port map( A => n14050, Z => n21553);
   U13978 : BUF_X1 port map( A => n14048, Z => n21556);
   U13979 : BUF_X1 port map( A => n14046, Z => n21559);
   U13980 : BUF_X1 port map( A => n14044, Z => n21562);
   U13981 : BUF_X1 port map( A => n14042, Z => n21565);
   U13982 : BUF_X1 port map( A => n14040, Z => n21568);
   U13983 : BUF_X1 port map( A => n14038, Z => n21571);
   U13984 : BUF_X1 port map( A => n14036, Z => n21574);
   U13985 : BUF_X1 port map( A => n14034, Z => n21577);
   U13986 : BUF_X1 port map( A => n14032, Z => n21580);
   U13987 : BUF_X1 port map( A => n14030, Z => n21583);
   U13988 : BUF_X1 port map( A => n14028, Z => n21586);
   U13989 : BUF_X1 port map( A => n14026, Z => n21589);
   U13990 : BUF_X1 port map( A => n14024, Z => n21592);
   U13991 : BUF_X1 port map( A => n14022, Z => n21595);
   U13992 : BUF_X1 port map( A => n14020, Z => n21598);
   U13993 : BUF_X1 port map( A => n14018, Z => n21601);
   U13994 : BUF_X1 port map( A => n14016, Z => n21604);
   U13995 : BUF_X1 port map( A => n14014, Z => n21607);
   U13996 : BUF_X1 port map( A => n14012, Z => n21610);
   U13997 : BUF_X1 port map( A => n14010, Z => n21613);
   U13998 : BUF_X1 port map( A => n14008, Z => n21616);
   U13999 : BUF_X1 port map( A => n14006, Z => n21619);
   U14000 : BUF_X1 port map( A => n14004, Z => n21622);
   U14001 : BUF_X1 port map( A => n14002, Z => n21625);
   U14002 : BUF_X1 port map( A => n14000, Z => n21628);
   U14003 : BUF_X1 port map( A => n13998, Z => n21631);
   U14004 : BUF_X1 port map( A => n13996, Z => n21634);
   U14005 : BUF_X1 port map( A => n13994, Z => n21637);
   U14006 : BUF_X1 port map( A => n13992, Z => n21640);
   U14007 : BUF_X1 port map( A => n13990, Z => n21643);
   U14008 : BUF_X1 port map( A => n13988, Z => n21646);
   U14009 : BUF_X1 port map( A => n13986, Z => n21649);
   U14010 : BUF_X1 port map( A => n13984, Z => n21652);
   U14011 : BUF_X1 port map( A => n13982, Z => n21655);
   U14012 : BUF_X1 port map( A => n13980, Z => n21658);
   U14013 : BUF_X1 port map( A => n13978, Z => n21661);
   U14014 : BUF_X1 port map( A => n13976, Z => n21664);
   U14015 : BUF_X1 port map( A => n13974, Z => n21667);
   U14016 : BUF_X1 port map( A => n13972, Z => n21670);
   U14017 : BUF_X1 port map( A => n13970, Z => n21673);
   U14018 : BUF_X1 port map( A => n13968, Z => n21676);
   U14019 : BUF_X1 port map( A => n13966, Z => n21679);
   U14020 : BUF_X1 port map( A => n13964, Z => n21682);
   U14021 : BUF_X1 port map( A => n13962, Z => n21685);
   U14022 : BUF_X1 port map( A => n13960, Z => n21688);
   U14023 : BUF_X1 port map( A => n13958, Z => n21691);
   U14024 : BUF_X1 port map( A => n13956, Z => n21694);
   U14025 : BUF_X1 port map( A => n13954, Z => n21697);
   U14026 : BUF_X1 port map( A => n13952, Z => n21700);
   U14027 : BUF_X1 port map( A => n13950, Z => n21703);
   U14028 : BUF_X1 port map( A => n13948, Z => n21706);
   U14029 : BUF_X1 port map( A => n13946, Z => n21709);
   U14030 : BUF_X1 port map( A => n13944, Z => n21712);
   U14031 : BUF_X1 port map( A => n13942, Z => n21715);
   U14032 : NAND2_X1 port map( A1 => n18517, A2 => n18514, ZN => n17345);
   U14033 : NAND2_X1 port map( A1 => n18524, A2 => n18514, ZN => n17355);
   U14034 : NAND2_X1 port map( A1 => n17316, A2 => n17313, ZN => n16078);
   U14035 : NAND2_X1 port map( A1 => n17323, A2 => n17313, ZN => n16089);
   U14036 : OAI22_X1 port map( A1 => n21128, A2 => n16162, B1 => n21708, B2 => 
                           n21121, ZN => n5430);
   U14037 : OAI22_X1 port map( A1 => n21128, A2 => n16143, B1 => n21711, B2 => 
                           n21121, ZN => n5432);
   U14038 : OAI22_X1 port map( A1 => n21128, A2 => n16124, B1 => n21714, B2 => 
                           n21121, ZN => n5434);
   U14039 : OAI22_X1 port map( A1 => n21128, A2 => n16070, B1 => n21717, B2 => 
                           n21121, ZN => n5436);
   U14040 : OAI22_X1 port map( A1 => n21141, A2 => n16008, B1 => n21708, B2 => 
                           n21134, ZN => n5497);
   U14041 : OAI22_X1 port map( A1 => n21141, A2 => n16007, B1 => n21711, B2 => 
                           n21134, ZN => n5498);
   U14042 : OAI22_X1 port map( A1 => n21141, A2 => n16006, B1 => n21714, B2 => 
                           n21134, ZN => n5499);
   U14043 : OAI22_X1 port map( A1 => n21141, A2 => n16004, B1 => n21717, B2 => 
                           n21134, ZN => n5500);
   U14044 : OAI22_X1 port map( A1 => n21167, A2 => n15876, B1 => n21708, B2 => 
                           n21160, ZN => n5625);
   U14045 : OAI22_X1 port map( A1 => n21167, A2 => n15875, B1 => n21711, B2 => 
                           n21160, ZN => n5626);
   U14046 : OAI22_X1 port map( A1 => n21167, A2 => n15874, B1 => n21714, B2 => 
                           n21160, ZN => n5627);
   U14047 : OAI22_X1 port map( A1 => n21167, A2 => n15872, B1 => n21717, B2 => 
                           n21160, ZN => n5628);
   U14048 : OAI22_X1 port map( A1 => n21193, A2 => n15744, B1 => n21708, B2 => 
                           n21186, ZN => n5753);
   U14049 : OAI22_X1 port map( A1 => n21193, A2 => n15743, B1 => n21711, B2 => 
                           n21186, ZN => n5754);
   U14050 : OAI22_X1 port map( A1 => n21193, A2 => n15742, B1 => n21714, B2 => 
                           n21186, ZN => n5755);
   U14051 : OAI22_X1 port map( A1 => n21193, A2 => n15740, B1 => n21717, B2 => 
                           n21186, ZN => n5756);
   U14052 : OAI22_X1 port map( A1 => n21219, A2 => n15608, B1 => n21707, B2 => 
                           n21212, ZN => n5881);
   U14053 : OAI22_X1 port map( A1 => n21219, A2 => n15607, B1 => n21710, B2 => 
                           n21212, ZN => n5882);
   U14054 : OAI22_X1 port map( A1 => n21219, A2 => n15606, B1 => n21713, B2 => 
                           n21212, ZN => n5883);
   U14055 : OAI22_X1 port map( A1 => n21219, A2 => n15604, B1 => n21716, B2 => 
                           n21212, ZN => n5884);
   U14056 : OAI22_X1 port map( A1 => n21258, A2 => n15409, B1 => n21707, B2 => 
                           n21251, ZN => n6073);
   U14057 : OAI22_X1 port map( A1 => n21258, A2 => n15408, B1 => n21710, B2 => 
                           n21251, ZN => n6074);
   U14058 : OAI22_X1 port map( A1 => n21258, A2 => n15407, B1 => n21713, B2 => 
                           n21251, ZN => n6075);
   U14059 : OAI22_X1 port map( A1 => n21258, A2 => n15405, B1 => n21716, B2 => 
                           n21251, ZN => n6076);
   U14060 : OAI22_X1 port map( A1 => n21284, A2 => n15277, B1 => n21707, B2 => 
                           n21277, ZN => n6201);
   U14061 : OAI22_X1 port map( A1 => n21284, A2 => n15276, B1 => n21710, B2 => 
                           n21277, ZN => n6202);
   U14062 : OAI22_X1 port map( A1 => n21284, A2 => n15275, B1 => n21713, B2 => 
                           n21277, ZN => n6203);
   U14063 : OAI22_X1 port map( A1 => n21284, A2 => n15273, B1 => n21716, B2 => 
                           n21277, ZN => n6204);
   U14064 : OAI22_X1 port map( A1 => n21336, A2 => n15010, B1 => n21707, B2 => 
                           n21329, ZN => n6457);
   U14065 : OAI22_X1 port map( A1 => n21336, A2 => n15009, B1 => n21710, B2 => 
                           n21329, ZN => n6458);
   U14066 : OAI22_X1 port map( A1 => n21336, A2 => n15008, B1 => n21713, B2 => 
                           n21329, ZN => n6459);
   U14067 : OAI22_X1 port map( A1 => n21336, A2 => n15006, B1 => n21716, B2 => 
                           n21329, ZN => n6460);
   U14068 : OAI22_X1 port map( A1 => n21349, A2 => n14944, B1 => n21707, B2 => 
                           n21342, ZN => n6521);
   U14069 : OAI22_X1 port map( A1 => n21349, A2 => n14943, B1 => n21710, B2 => 
                           n21342, ZN => n6522);
   U14070 : OAI22_X1 port map( A1 => n21349, A2 => n14942, B1 => n21713, B2 => 
                           n21342, ZN => n6523);
   U14071 : OAI22_X1 port map( A1 => n21349, A2 => n14940, B1 => n21716, B2 => 
                           n21342, ZN => n6524);
   U14072 : OAI22_X1 port map( A1 => n21362, A2 => n14878, B1 => n21707, B2 => 
                           n21355, ZN => n6585);
   U14073 : OAI22_X1 port map( A1 => n21362, A2 => n14877, B1 => n21710, B2 => 
                           n21355, ZN => n6586);
   U14074 : OAI22_X1 port map( A1 => n21362, A2 => n14876, B1 => n21713, B2 => 
                           n21355, ZN => n6587);
   U14075 : OAI22_X1 port map( A1 => n21362, A2 => n14874, B1 => n21716, B2 => 
                           n21355, ZN => n6588);
   U14076 : OAI22_X1 port map( A1 => n21375, A2 => n14812, B1 => n21707, B2 => 
                           n21368, ZN => n6649);
   U14077 : OAI22_X1 port map( A1 => n21375, A2 => n14811, B1 => n21710, B2 => 
                           n21368, ZN => n6650);
   U14078 : OAI22_X1 port map( A1 => n21375, A2 => n14810, B1 => n21713, B2 => 
                           n21368, ZN => n6651);
   U14079 : OAI22_X1 port map( A1 => n21375, A2 => n14808, B1 => n21716, B2 => 
                           n21368, ZN => n6652);
   U14080 : OAI22_X1 port map( A1 => n21388, A2 => n14746, B1 => n21706, B2 => 
                           n21381, ZN => n6713);
   U14081 : OAI22_X1 port map( A1 => n21388, A2 => n14745, B1 => n21709, B2 => 
                           n21381, ZN => n6714);
   U14082 : OAI22_X1 port map( A1 => n21388, A2 => n14744, B1 => n21712, B2 => 
                           n21381, ZN => n6715);
   U14083 : OAI22_X1 port map( A1 => n21388, A2 => n14742, B1 => n21715, B2 => 
                           n21381, ZN => n6716);
   U14084 : OAI22_X1 port map( A1 => n21427, A2 => n14546, B1 => n21706, B2 => 
                           n21420, ZN => n6905);
   U14085 : OAI22_X1 port map( A1 => n21427, A2 => n14545, B1 => n21709, B2 => 
                           n21420, ZN => n6906);
   U14086 : OAI22_X1 port map( A1 => n21427, A2 => n14544, B1 => n21712, B2 => 
                           n21420, ZN => n6907);
   U14087 : OAI22_X1 port map( A1 => n21427, A2 => n14542, B1 => n21715, B2 => 
                           n21420, ZN => n6908);
   U14088 : OAI22_X1 port map( A1 => n21440, A2 => n14480, B1 => n21706, B2 => 
                           n21433, ZN => n6969);
   U14089 : OAI22_X1 port map( A1 => n21440, A2 => n14479, B1 => n21709, B2 => 
                           n21433, ZN => n6970);
   U14090 : OAI22_X1 port map( A1 => n21440, A2 => n14478, B1 => n21712, B2 => 
                           n21433, ZN => n6971);
   U14091 : OAI22_X1 port map( A1 => n21440, A2 => n14476, B1 => n21715, B2 => 
                           n21433, ZN => n6972);
   U14092 : OAI22_X1 port map( A1 => n21466, A2 => n14344, B1 => n21706, B2 => 
                           n21459, ZN => n7097);
   U14093 : OAI22_X1 port map( A1 => n21466, A2 => n14343, B1 => n21709, B2 => 
                           n21459, ZN => n7098);
   U14094 : OAI22_X1 port map( A1 => n21466, A2 => n14342, B1 => n21712, B2 => 
                           n21459, ZN => n7099);
   U14095 : OAI22_X1 port map( A1 => n21466, A2 => n14340, B1 => n21715, B2 => 
                           n21459, ZN => n7100);
   U14096 : OAI22_X1 port map( A1 => n21479, A2 => n14277, B1 => n21706, B2 => 
                           n21472, ZN => n7161);
   U14097 : OAI22_X1 port map( A1 => n21479, A2 => n14276, B1 => n21709, B2 => 
                           n21472, ZN => n7162);
   U14098 : OAI22_X1 port map( A1 => n21479, A2 => n14275, B1 => n21712, B2 => 
                           n21472, ZN => n7163);
   U14099 : OAI22_X1 port map( A1 => n21479, A2 => n14273, B1 => n21715, B2 => 
                           n21472, ZN => n7164);
   U14100 : OAI22_X1 port map( A1 => n21492, A2 => n14211, B1 => n21706, B2 => 
                           n21485, ZN => n7225);
   U14101 : OAI22_X1 port map( A1 => n21492, A2 => n14210, B1 => n21709, B2 => 
                           n21485, ZN => n7226);
   U14102 : OAI22_X1 port map( A1 => n21492, A2 => n14209, B1 => n21712, B2 => 
                           n21485, ZN => n7227);
   U14103 : OAI22_X1 port map( A1 => n21492, A2 => n14207, B1 => n21715, B2 => 
                           n21485, ZN => n7228);
   U14104 : OAI22_X1 port map( A1 => n21518, A2 => n14077, B1 => n21706, B2 => 
                           n21511, ZN => n7353);
   U14105 : OAI22_X1 port map( A1 => n21518, A2 => n14076, B1 => n21709, B2 => 
                           n21511, ZN => n7354);
   U14106 : OAI22_X1 port map( A1 => n21518, A2 => n14075, B1 => n21712, B2 => 
                           n21511, ZN => n7355);
   U14107 : OAI22_X1 port map( A1 => n21518, A2 => n14073, B1 => n21715, B2 => 
                           n21511, ZN => n7356);
   U14108 : NAND2_X1 port map( A1 => n18517, A2 => n18520, ZN => n17360);
   U14109 : NAND2_X1 port map( A1 => n17316, A2 => n17320, ZN => n16094);
   U14110 : NAND2_X1 port map( A1 => n18516, A2 => n18512, ZN => n17370);
   U14111 : OAI22_X1 port map( A1 => n21124, A2 => n17302, B1 => n21528, B2 => 
                           n21116, ZN => n5310);
   U14112 : OAI22_X1 port map( A1 => n21124, A2 => n17283, B1 => n21531, B2 => 
                           n21116, ZN => n5312);
   U14113 : OAI22_X1 port map( A1 => n21124, A2 => n17264, B1 => n21534, B2 => 
                           n21116, ZN => n5314);
   U14114 : OAI22_X1 port map( A1 => n21124, A2 => n17245, B1 => n21537, B2 => 
                           n21116, ZN => n5316);
   U14115 : OAI22_X1 port map( A1 => n21124, A2 => n17226, B1 => n21540, B2 => 
                           n21116, ZN => n5318);
   U14116 : OAI22_X1 port map( A1 => n21124, A2 => n17207, B1 => n21543, B2 => 
                           n21116, ZN => n5320);
   U14117 : OAI22_X1 port map( A1 => n21124, A2 => n17188, B1 => n21546, B2 => 
                           n21116, ZN => n5322);
   U14118 : OAI22_X1 port map( A1 => n21124, A2 => n17169, B1 => n21549, B2 => 
                           n21116, ZN => n5324);
   U14119 : OAI22_X1 port map( A1 => n21124, A2 => n17150, B1 => n21552, B2 => 
                           n21116, ZN => n5326);
   U14120 : OAI22_X1 port map( A1 => n21124, A2 => n17131, B1 => n21555, B2 => 
                           n21116, ZN => n5328);
   U14121 : OAI22_X1 port map( A1 => n21124, A2 => n17112, B1 => n21558, B2 => 
                           n21116, ZN => n5330);
   U14122 : OAI22_X1 port map( A1 => n21124, A2 => n17093, B1 => n21561, B2 => 
                           n21116, ZN => n5332);
   U14123 : OAI22_X1 port map( A1 => n21125, A2 => n17074, B1 => n21564, B2 => 
                           n21117, ZN => n5334);
   U14124 : OAI22_X1 port map( A1 => n21125, A2 => n17055, B1 => n21567, B2 => 
                           n21117, ZN => n5336);
   U14125 : OAI22_X1 port map( A1 => n21125, A2 => n17036, B1 => n21570, B2 => 
                           n21117, ZN => n5338);
   U14126 : OAI22_X1 port map( A1 => n21125, A2 => n17017, B1 => n21573, B2 => 
                           n21117, ZN => n5340);
   U14127 : OAI22_X1 port map( A1 => n21125, A2 => n16998, B1 => n21576, B2 => 
                           n21117, ZN => n5342);
   U14128 : OAI22_X1 port map( A1 => n21125, A2 => n16979, B1 => n21579, B2 => 
                           n21117, ZN => n5344);
   U14129 : OAI22_X1 port map( A1 => n21125, A2 => n16960, B1 => n21582, B2 => 
                           n21117, ZN => n5346);
   U14130 : OAI22_X1 port map( A1 => n21125, A2 => n16941, B1 => n21585, B2 => 
                           n21117, ZN => n5348);
   U14131 : OAI22_X1 port map( A1 => n21125, A2 => n16922, B1 => n21588, B2 => 
                           n21117, ZN => n5350);
   U14132 : OAI22_X1 port map( A1 => n21125, A2 => n16903, B1 => n21591, B2 => 
                           n21117, ZN => n5352);
   U14133 : OAI22_X1 port map( A1 => n21125, A2 => n16884, B1 => n21594, B2 => 
                           n21117, ZN => n5354);
   U14134 : OAI22_X1 port map( A1 => n21125, A2 => n16865, B1 => n21597, B2 => 
                           n21117, ZN => n5356);
   U14135 : OAI22_X1 port map( A1 => n21125, A2 => n16846, B1 => n21600, B2 => 
                           n21118, ZN => n5358);
   U14136 : OAI22_X1 port map( A1 => n21126, A2 => n16827, B1 => n21603, B2 => 
                           n21118, ZN => n5360);
   U14137 : OAI22_X1 port map( A1 => n21126, A2 => n16808, B1 => n21606, B2 => 
                           n21118, ZN => n5362);
   U14138 : OAI22_X1 port map( A1 => n21126, A2 => n16789, B1 => n21609, B2 => 
                           n21118, ZN => n5364);
   U14139 : OAI22_X1 port map( A1 => n21126, A2 => n16770, B1 => n21612, B2 => 
                           n21118, ZN => n5366);
   U14140 : OAI22_X1 port map( A1 => n21126, A2 => n16751, B1 => n21615, B2 => 
                           n21118, ZN => n5368);
   U14141 : OAI22_X1 port map( A1 => n21126, A2 => n16732, B1 => n21618, B2 => 
                           n21118, ZN => n5370);
   U14142 : OAI22_X1 port map( A1 => n21126, A2 => n16713, B1 => n21621, B2 => 
                           n21118, ZN => n5372);
   U14143 : OAI22_X1 port map( A1 => n21126, A2 => n16694, B1 => n21624, B2 => 
                           n21118, ZN => n5374);
   U14144 : OAI22_X1 port map( A1 => n21126, A2 => n16675, B1 => n21627, B2 => 
                           n21118, ZN => n5376);
   U14145 : OAI22_X1 port map( A1 => n21126, A2 => n16656, B1 => n21630, B2 => 
                           n21118, ZN => n5378);
   U14146 : OAI22_X1 port map( A1 => n21126, A2 => n16637, B1 => n21633, B2 => 
                           n21118, ZN => n5380);
   U14147 : OAI22_X1 port map( A1 => n21126, A2 => n16618, B1 => n21636, B2 => 
                           n21119, ZN => n5382);
   U14148 : OAI22_X1 port map( A1 => n21126, A2 => n16599, B1 => n21639, B2 => 
                           n21119, ZN => n5384);
   U14149 : OAI22_X1 port map( A1 => n21127, A2 => n16580, B1 => n21642, B2 => 
                           n21119, ZN => n5386);
   U14150 : OAI22_X1 port map( A1 => n21127, A2 => n16561, B1 => n21645, B2 => 
                           n21119, ZN => n5388);
   U14151 : OAI22_X1 port map( A1 => n21127, A2 => n16542, B1 => n21648, B2 => 
                           n21119, ZN => n5390);
   U14152 : OAI22_X1 port map( A1 => n21127, A2 => n16523, B1 => n21651, B2 => 
                           n21119, ZN => n5392);
   U14153 : OAI22_X1 port map( A1 => n21127, A2 => n16504, B1 => n21654, B2 => 
                           n21119, ZN => n5394);
   U14154 : OAI22_X1 port map( A1 => n21127, A2 => n16485, B1 => n21657, B2 => 
                           n21119, ZN => n5396);
   U14155 : OAI22_X1 port map( A1 => n21127, A2 => n16466, B1 => n21660, B2 => 
                           n21119, ZN => n5398);
   U14156 : OAI22_X1 port map( A1 => n21127, A2 => n16447, B1 => n21663, B2 => 
                           n21119, ZN => n5400);
   U14157 : OAI22_X1 port map( A1 => n21127, A2 => n16428, B1 => n21666, B2 => 
                           n21119, ZN => n5402);
   U14158 : OAI22_X1 port map( A1 => n21127, A2 => n16409, B1 => n21669, B2 => 
                           n21119, ZN => n5404);
   U14159 : OAI22_X1 port map( A1 => n21127, A2 => n16390, B1 => n21672, B2 => 
                           n21120, ZN => n5406);
   U14160 : OAI22_X1 port map( A1 => n21127, A2 => n16371, B1 => n21675, B2 => 
                           n21120, ZN => n5408);
   U14161 : OAI22_X1 port map( A1 => n21127, A2 => n16352, B1 => n21678, B2 => 
                           n21120, ZN => n5410);
   U14162 : OAI22_X1 port map( A1 => n21128, A2 => n16333, B1 => n21681, B2 => 
                           n21120, ZN => n5412);
   U14163 : OAI22_X1 port map( A1 => n21128, A2 => n16314, B1 => n21684, B2 => 
                           n21120, ZN => n5414);
   U14164 : OAI22_X1 port map( A1 => n21128, A2 => n16295, B1 => n21687, B2 => 
                           n21120, ZN => n5416);
   U14165 : OAI22_X1 port map( A1 => n21128, A2 => n16276, B1 => n21690, B2 => 
                           n21120, ZN => n5418);
   U14166 : OAI22_X1 port map( A1 => n21128, A2 => n16257, B1 => n21693, B2 => 
                           n21120, ZN => n5420);
   U14167 : OAI22_X1 port map( A1 => n21128, A2 => n16238, B1 => n21696, B2 => 
                           n21120, ZN => n5422);
   U14168 : OAI22_X1 port map( A1 => n21128, A2 => n16219, B1 => n21699, B2 => 
                           n21120, ZN => n5424);
   U14169 : OAI22_X1 port map( A1 => n21128, A2 => n16200, B1 => n21702, B2 => 
                           n21120, ZN => n5426);
   U14170 : OAI22_X1 port map( A1 => n21128, A2 => n16181, B1 => n21705, B2 => 
                           n21120, ZN => n5428);
   U14171 : OAI22_X1 port map( A1 => n21137, A2 => n16068, B1 => n21528, B2 => 
                           n21129, ZN => n5437);
   U14172 : OAI22_X1 port map( A1 => n21137, A2 => n16067, B1 => n21531, B2 => 
                           n21129, ZN => n5438);
   U14173 : OAI22_X1 port map( A1 => n21137, A2 => n16066, B1 => n21534, B2 => 
                           n21129, ZN => n5439);
   U14174 : OAI22_X1 port map( A1 => n21137, A2 => n16065, B1 => n21537, B2 => 
                           n21129, ZN => n5440);
   U14175 : OAI22_X1 port map( A1 => n21137, A2 => n16064, B1 => n21540, B2 => 
                           n21129, ZN => n5441);
   U14176 : OAI22_X1 port map( A1 => n21137, A2 => n16063, B1 => n21543, B2 => 
                           n21129, ZN => n5442);
   U14177 : OAI22_X1 port map( A1 => n21137, A2 => n16062, B1 => n21546, B2 => 
                           n21129, ZN => n5443);
   U14178 : OAI22_X1 port map( A1 => n21137, A2 => n16061, B1 => n21549, B2 => 
                           n21129, ZN => n5444);
   U14179 : OAI22_X1 port map( A1 => n21137, A2 => n16060, B1 => n21552, B2 => 
                           n21129, ZN => n5445);
   U14180 : OAI22_X1 port map( A1 => n21137, A2 => n16059, B1 => n21555, B2 => 
                           n21129, ZN => n5446);
   U14181 : OAI22_X1 port map( A1 => n21137, A2 => n16058, B1 => n21558, B2 => 
                           n21129, ZN => n5447);
   U14182 : OAI22_X1 port map( A1 => n21137, A2 => n16057, B1 => n21561, B2 => 
                           n21129, ZN => n5448);
   U14183 : OAI22_X1 port map( A1 => n21138, A2 => n16056, B1 => n21564, B2 => 
                           n21130, ZN => n5449);
   U14184 : OAI22_X1 port map( A1 => n21138, A2 => n16055, B1 => n21567, B2 => 
                           n21130, ZN => n5450);
   U14185 : OAI22_X1 port map( A1 => n21138, A2 => n16054, B1 => n21570, B2 => 
                           n21130, ZN => n5451);
   U14186 : OAI22_X1 port map( A1 => n21138, A2 => n16053, B1 => n21573, B2 => 
                           n21130, ZN => n5452);
   U14187 : OAI22_X1 port map( A1 => n21138, A2 => n16052, B1 => n21576, B2 => 
                           n21130, ZN => n5453);
   U14188 : OAI22_X1 port map( A1 => n21138, A2 => n16051, B1 => n21579, B2 => 
                           n21130, ZN => n5454);
   U14189 : OAI22_X1 port map( A1 => n21138, A2 => n16050, B1 => n21582, B2 => 
                           n21130, ZN => n5455);
   U14190 : OAI22_X1 port map( A1 => n21138, A2 => n16049, B1 => n21585, B2 => 
                           n21130, ZN => n5456);
   U14191 : OAI22_X1 port map( A1 => n21138, A2 => n16048, B1 => n21588, B2 => 
                           n21130, ZN => n5457);
   U14192 : OAI22_X1 port map( A1 => n21138, A2 => n16047, B1 => n21591, B2 => 
                           n21130, ZN => n5458);
   U14193 : OAI22_X1 port map( A1 => n21138, A2 => n16046, B1 => n21594, B2 => 
                           n21130, ZN => n5459);
   U14194 : OAI22_X1 port map( A1 => n21138, A2 => n16045, B1 => n21597, B2 => 
                           n21130, ZN => n5460);
   U14195 : OAI22_X1 port map( A1 => n21138, A2 => n16044, B1 => n21600, B2 => 
                           n21131, ZN => n5461);
   U14196 : OAI22_X1 port map( A1 => n21139, A2 => n16043, B1 => n21603, B2 => 
                           n21131, ZN => n5462);
   U14197 : OAI22_X1 port map( A1 => n21139, A2 => n16042, B1 => n21606, B2 => 
                           n21131, ZN => n5463);
   U14198 : OAI22_X1 port map( A1 => n21139, A2 => n16041, B1 => n21609, B2 => 
                           n21131, ZN => n5464);
   U14199 : OAI22_X1 port map( A1 => n21139, A2 => n16040, B1 => n21612, B2 => 
                           n21131, ZN => n5465);
   U14200 : OAI22_X1 port map( A1 => n21139, A2 => n16039, B1 => n21615, B2 => 
                           n21131, ZN => n5466);
   U14201 : OAI22_X1 port map( A1 => n21139, A2 => n16038, B1 => n21618, B2 => 
                           n21131, ZN => n5467);
   U14202 : OAI22_X1 port map( A1 => n21139, A2 => n16037, B1 => n21621, B2 => 
                           n21131, ZN => n5468);
   U14203 : OAI22_X1 port map( A1 => n21139, A2 => n16036, B1 => n21624, B2 => 
                           n21131, ZN => n5469);
   U14204 : OAI22_X1 port map( A1 => n21139, A2 => n16035, B1 => n21627, B2 => 
                           n21131, ZN => n5470);
   U14205 : OAI22_X1 port map( A1 => n21139, A2 => n16034, B1 => n21630, B2 => 
                           n21131, ZN => n5471);
   U14206 : OAI22_X1 port map( A1 => n21139, A2 => n16033, B1 => n21633, B2 => 
                           n21131, ZN => n5472);
   U14207 : OAI22_X1 port map( A1 => n21139, A2 => n16032, B1 => n21636, B2 => 
                           n21132, ZN => n5473);
   U14208 : OAI22_X1 port map( A1 => n21139, A2 => n16031, B1 => n21639, B2 => 
                           n21132, ZN => n5474);
   U14209 : OAI22_X1 port map( A1 => n21140, A2 => n16030, B1 => n21642, B2 => 
                           n21132, ZN => n5475);
   U14210 : OAI22_X1 port map( A1 => n21140, A2 => n16029, B1 => n21645, B2 => 
                           n21132, ZN => n5476);
   U14211 : OAI22_X1 port map( A1 => n21140, A2 => n16028, B1 => n21648, B2 => 
                           n21132, ZN => n5477);
   U14212 : OAI22_X1 port map( A1 => n21140, A2 => n16027, B1 => n21651, B2 => 
                           n21132, ZN => n5478);
   U14213 : OAI22_X1 port map( A1 => n21140, A2 => n16026, B1 => n21654, B2 => 
                           n21132, ZN => n5479);
   U14214 : OAI22_X1 port map( A1 => n21140, A2 => n16025, B1 => n21657, B2 => 
                           n21132, ZN => n5480);
   U14215 : OAI22_X1 port map( A1 => n21140, A2 => n16024, B1 => n21660, B2 => 
                           n21132, ZN => n5481);
   U14216 : OAI22_X1 port map( A1 => n21140, A2 => n16023, B1 => n21663, B2 => 
                           n21132, ZN => n5482);
   U14217 : OAI22_X1 port map( A1 => n21140, A2 => n16022, B1 => n21666, B2 => 
                           n21132, ZN => n5483);
   U14218 : OAI22_X1 port map( A1 => n21140, A2 => n16021, B1 => n21669, B2 => 
                           n21132, ZN => n5484);
   U14219 : OAI22_X1 port map( A1 => n21140, A2 => n16020, B1 => n21672, B2 => 
                           n21133, ZN => n5485);
   U14220 : OAI22_X1 port map( A1 => n21140, A2 => n16019, B1 => n21675, B2 => 
                           n21133, ZN => n5486);
   U14221 : OAI22_X1 port map( A1 => n21140, A2 => n16018, B1 => n21678, B2 => 
                           n21133, ZN => n5487);
   U14222 : OAI22_X1 port map( A1 => n21141, A2 => n16017, B1 => n21681, B2 => 
                           n21133, ZN => n5488);
   U14223 : OAI22_X1 port map( A1 => n21141, A2 => n16016, B1 => n21684, B2 => 
                           n21133, ZN => n5489);
   U14224 : OAI22_X1 port map( A1 => n21141, A2 => n16015, B1 => n21687, B2 => 
                           n21133, ZN => n5490);
   U14225 : OAI22_X1 port map( A1 => n21141, A2 => n16014, B1 => n21690, B2 => 
                           n21133, ZN => n5491);
   U14226 : OAI22_X1 port map( A1 => n21141, A2 => n16013, B1 => n21693, B2 => 
                           n21133, ZN => n5492);
   U14227 : OAI22_X1 port map( A1 => n21141, A2 => n16012, B1 => n21696, B2 => 
                           n21133, ZN => n5493);
   U14228 : OAI22_X1 port map( A1 => n21141, A2 => n16011, B1 => n21699, B2 => 
                           n21133, ZN => n5494);
   U14229 : OAI22_X1 port map( A1 => n21141, A2 => n16010, B1 => n21702, B2 => 
                           n21133, ZN => n5495);
   U14230 : OAI22_X1 port map( A1 => n21141, A2 => n16009, B1 => n21705, B2 => 
                           n21133, ZN => n5496);
   U14231 : OAI22_X1 port map( A1 => n21163, A2 => n15936, B1 => n21528, B2 => 
                           n21155, ZN => n5565);
   U14232 : OAI22_X1 port map( A1 => n21163, A2 => n15935, B1 => n21531, B2 => 
                           n21155, ZN => n5566);
   U14233 : OAI22_X1 port map( A1 => n21163, A2 => n15934, B1 => n21534, B2 => 
                           n21155, ZN => n5567);
   U14234 : OAI22_X1 port map( A1 => n21163, A2 => n15933, B1 => n21537, B2 => 
                           n21155, ZN => n5568);
   U14235 : OAI22_X1 port map( A1 => n21163, A2 => n15932, B1 => n21540, B2 => 
                           n21155, ZN => n5569);
   U14236 : OAI22_X1 port map( A1 => n21163, A2 => n15931, B1 => n21543, B2 => 
                           n21155, ZN => n5570);
   U14237 : OAI22_X1 port map( A1 => n21163, A2 => n15930, B1 => n21546, B2 => 
                           n21155, ZN => n5571);
   U14238 : OAI22_X1 port map( A1 => n21163, A2 => n15929, B1 => n21549, B2 => 
                           n21155, ZN => n5572);
   U14239 : OAI22_X1 port map( A1 => n21163, A2 => n15928, B1 => n21552, B2 => 
                           n21155, ZN => n5573);
   U14240 : OAI22_X1 port map( A1 => n21163, A2 => n15927, B1 => n21555, B2 => 
                           n21155, ZN => n5574);
   U14241 : OAI22_X1 port map( A1 => n21163, A2 => n15926, B1 => n21558, B2 => 
                           n21155, ZN => n5575);
   U14242 : OAI22_X1 port map( A1 => n21163, A2 => n15925, B1 => n21561, B2 => 
                           n21155, ZN => n5576);
   U14243 : OAI22_X1 port map( A1 => n21164, A2 => n15924, B1 => n21564, B2 => 
                           n21156, ZN => n5577);
   U14244 : OAI22_X1 port map( A1 => n21164, A2 => n15923, B1 => n21567, B2 => 
                           n21156, ZN => n5578);
   U14245 : OAI22_X1 port map( A1 => n21164, A2 => n15922, B1 => n21570, B2 => 
                           n21156, ZN => n5579);
   U14246 : OAI22_X1 port map( A1 => n21164, A2 => n15921, B1 => n21573, B2 => 
                           n21156, ZN => n5580);
   U14247 : OAI22_X1 port map( A1 => n21164, A2 => n15920, B1 => n21576, B2 => 
                           n21156, ZN => n5581);
   U14248 : OAI22_X1 port map( A1 => n21164, A2 => n15919, B1 => n21579, B2 => 
                           n21156, ZN => n5582);
   U14249 : OAI22_X1 port map( A1 => n21164, A2 => n15918, B1 => n21582, B2 => 
                           n21156, ZN => n5583);
   U14250 : OAI22_X1 port map( A1 => n21164, A2 => n15917, B1 => n21585, B2 => 
                           n21156, ZN => n5584);
   U14251 : OAI22_X1 port map( A1 => n21164, A2 => n15916, B1 => n21588, B2 => 
                           n21156, ZN => n5585);
   U14252 : OAI22_X1 port map( A1 => n21164, A2 => n15915, B1 => n21591, B2 => 
                           n21156, ZN => n5586);
   U14253 : OAI22_X1 port map( A1 => n21164, A2 => n15914, B1 => n21594, B2 => 
                           n21156, ZN => n5587);
   U14254 : OAI22_X1 port map( A1 => n21164, A2 => n15913, B1 => n21597, B2 => 
                           n21156, ZN => n5588);
   U14255 : OAI22_X1 port map( A1 => n21164, A2 => n15912, B1 => n21600, B2 => 
                           n21157, ZN => n5589);
   U14256 : OAI22_X1 port map( A1 => n21165, A2 => n15911, B1 => n21603, B2 => 
                           n21157, ZN => n5590);
   U14257 : OAI22_X1 port map( A1 => n21165, A2 => n15910, B1 => n21606, B2 => 
                           n21157, ZN => n5591);
   U14258 : OAI22_X1 port map( A1 => n21165, A2 => n15909, B1 => n21609, B2 => 
                           n21157, ZN => n5592);
   U14259 : OAI22_X1 port map( A1 => n21165, A2 => n15908, B1 => n21612, B2 => 
                           n21157, ZN => n5593);
   U14260 : OAI22_X1 port map( A1 => n21165, A2 => n15907, B1 => n21615, B2 => 
                           n21157, ZN => n5594);
   U14261 : OAI22_X1 port map( A1 => n21165, A2 => n15906, B1 => n21618, B2 => 
                           n21157, ZN => n5595);
   U14262 : OAI22_X1 port map( A1 => n21165, A2 => n15905, B1 => n21621, B2 => 
                           n21157, ZN => n5596);
   U14263 : OAI22_X1 port map( A1 => n21165, A2 => n15904, B1 => n21624, B2 => 
                           n21157, ZN => n5597);
   U14264 : OAI22_X1 port map( A1 => n21165, A2 => n15903, B1 => n21627, B2 => 
                           n21157, ZN => n5598);
   U14265 : OAI22_X1 port map( A1 => n21165, A2 => n15902, B1 => n21630, B2 => 
                           n21157, ZN => n5599);
   U14266 : OAI22_X1 port map( A1 => n21165, A2 => n15901, B1 => n21633, B2 => 
                           n21157, ZN => n5600);
   U14267 : OAI22_X1 port map( A1 => n21165, A2 => n15900, B1 => n21636, B2 => 
                           n21158, ZN => n5601);
   U14268 : OAI22_X1 port map( A1 => n21165, A2 => n15899, B1 => n21639, B2 => 
                           n21158, ZN => n5602);
   U14269 : OAI22_X1 port map( A1 => n21166, A2 => n15898, B1 => n21642, B2 => 
                           n21158, ZN => n5603);
   U14270 : OAI22_X1 port map( A1 => n21166, A2 => n15897, B1 => n21645, B2 => 
                           n21158, ZN => n5604);
   U14271 : OAI22_X1 port map( A1 => n21166, A2 => n15896, B1 => n21648, B2 => 
                           n21158, ZN => n5605);
   U14272 : OAI22_X1 port map( A1 => n21166, A2 => n15895, B1 => n21651, B2 => 
                           n21158, ZN => n5606);
   U14273 : OAI22_X1 port map( A1 => n21166, A2 => n15894, B1 => n21654, B2 => 
                           n21158, ZN => n5607);
   U14274 : OAI22_X1 port map( A1 => n21166, A2 => n15893, B1 => n21657, B2 => 
                           n21158, ZN => n5608);
   U14275 : OAI22_X1 port map( A1 => n21166, A2 => n15892, B1 => n21660, B2 => 
                           n21158, ZN => n5609);
   U14276 : OAI22_X1 port map( A1 => n21166, A2 => n15891, B1 => n21663, B2 => 
                           n21158, ZN => n5610);
   U14277 : OAI22_X1 port map( A1 => n21166, A2 => n15890, B1 => n21666, B2 => 
                           n21158, ZN => n5611);
   U14278 : OAI22_X1 port map( A1 => n21166, A2 => n15889, B1 => n21669, B2 => 
                           n21158, ZN => n5612);
   U14279 : OAI22_X1 port map( A1 => n21166, A2 => n15888, B1 => n21672, B2 => 
                           n21159, ZN => n5613);
   U14280 : OAI22_X1 port map( A1 => n21166, A2 => n15887, B1 => n21675, B2 => 
                           n21159, ZN => n5614);
   U14281 : OAI22_X1 port map( A1 => n21166, A2 => n15886, B1 => n21678, B2 => 
                           n21159, ZN => n5615);
   U14282 : OAI22_X1 port map( A1 => n21167, A2 => n15885, B1 => n21681, B2 => 
                           n21159, ZN => n5616);
   U14283 : OAI22_X1 port map( A1 => n21167, A2 => n15884, B1 => n21684, B2 => 
                           n21159, ZN => n5617);
   U14284 : OAI22_X1 port map( A1 => n21167, A2 => n15883, B1 => n21687, B2 => 
                           n21159, ZN => n5618);
   U14285 : OAI22_X1 port map( A1 => n21167, A2 => n15882, B1 => n21690, B2 => 
                           n21159, ZN => n5619);
   U14286 : OAI22_X1 port map( A1 => n21167, A2 => n15881, B1 => n21693, B2 => 
                           n21159, ZN => n5620);
   U14287 : OAI22_X1 port map( A1 => n21167, A2 => n15880, B1 => n21696, B2 => 
                           n21159, ZN => n5621);
   U14288 : OAI22_X1 port map( A1 => n21167, A2 => n15879, B1 => n21699, B2 => 
                           n21159, ZN => n5622);
   U14289 : OAI22_X1 port map( A1 => n21167, A2 => n15878, B1 => n21702, B2 => 
                           n21159, ZN => n5623);
   U14290 : OAI22_X1 port map( A1 => n21167, A2 => n15877, B1 => n21705, B2 => 
                           n21159, ZN => n5624);
   U14291 : OAI22_X1 port map( A1 => n21189, A2 => n15804, B1 => n21528, B2 => 
                           n21181, ZN => n5693);
   U14292 : OAI22_X1 port map( A1 => n21189, A2 => n15803, B1 => n21531, B2 => 
                           n21181, ZN => n5694);
   U14293 : OAI22_X1 port map( A1 => n21189, A2 => n15802, B1 => n21534, B2 => 
                           n21181, ZN => n5695);
   U14294 : OAI22_X1 port map( A1 => n21189, A2 => n15801, B1 => n21537, B2 => 
                           n21181, ZN => n5696);
   U14295 : OAI22_X1 port map( A1 => n21189, A2 => n15800, B1 => n21540, B2 => 
                           n21181, ZN => n5697);
   U14296 : OAI22_X1 port map( A1 => n21189, A2 => n15799, B1 => n21543, B2 => 
                           n21181, ZN => n5698);
   U14297 : OAI22_X1 port map( A1 => n21189, A2 => n15798, B1 => n21546, B2 => 
                           n21181, ZN => n5699);
   U14298 : OAI22_X1 port map( A1 => n21189, A2 => n15797, B1 => n21549, B2 => 
                           n21181, ZN => n5700);
   U14299 : OAI22_X1 port map( A1 => n21189, A2 => n15796, B1 => n21552, B2 => 
                           n21181, ZN => n5701);
   U14300 : OAI22_X1 port map( A1 => n21189, A2 => n15795, B1 => n21555, B2 => 
                           n21181, ZN => n5702);
   U14301 : OAI22_X1 port map( A1 => n21189, A2 => n15794, B1 => n21558, B2 => 
                           n21181, ZN => n5703);
   U14302 : OAI22_X1 port map( A1 => n21189, A2 => n15793, B1 => n21561, B2 => 
                           n21181, ZN => n5704);
   U14303 : OAI22_X1 port map( A1 => n21190, A2 => n15792, B1 => n21564, B2 => 
                           n21182, ZN => n5705);
   U14304 : OAI22_X1 port map( A1 => n21190, A2 => n15791, B1 => n21567, B2 => 
                           n21182, ZN => n5706);
   U14305 : OAI22_X1 port map( A1 => n21190, A2 => n15790, B1 => n21570, B2 => 
                           n21182, ZN => n5707);
   U14306 : OAI22_X1 port map( A1 => n21190, A2 => n15789, B1 => n21573, B2 => 
                           n21182, ZN => n5708);
   U14307 : OAI22_X1 port map( A1 => n21190, A2 => n15788, B1 => n21576, B2 => 
                           n21182, ZN => n5709);
   U14308 : OAI22_X1 port map( A1 => n21190, A2 => n15787, B1 => n21579, B2 => 
                           n21182, ZN => n5710);
   U14309 : OAI22_X1 port map( A1 => n21190, A2 => n15786, B1 => n21582, B2 => 
                           n21182, ZN => n5711);
   U14310 : OAI22_X1 port map( A1 => n21190, A2 => n15785, B1 => n21585, B2 => 
                           n21182, ZN => n5712);
   U14311 : OAI22_X1 port map( A1 => n21190, A2 => n15784, B1 => n21588, B2 => 
                           n21182, ZN => n5713);
   U14312 : OAI22_X1 port map( A1 => n21190, A2 => n15783, B1 => n21591, B2 => 
                           n21182, ZN => n5714);
   U14313 : OAI22_X1 port map( A1 => n21190, A2 => n15782, B1 => n21594, B2 => 
                           n21182, ZN => n5715);
   U14314 : OAI22_X1 port map( A1 => n21190, A2 => n15781, B1 => n21597, B2 => 
                           n21182, ZN => n5716);
   U14315 : OAI22_X1 port map( A1 => n21190, A2 => n15780, B1 => n21600, B2 => 
                           n21183, ZN => n5717);
   U14316 : OAI22_X1 port map( A1 => n21191, A2 => n15779, B1 => n21603, B2 => 
                           n21183, ZN => n5718);
   U14317 : OAI22_X1 port map( A1 => n21191, A2 => n15778, B1 => n21606, B2 => 
                           n21183, ZN => n5719);
   U14318 : OAI22_X1 port map( A1 => n21191, A2 => n15777, B1 => n21609, B2 => 
                           n21183, ZN => n5720);
   U14319 : OAI22_X1 port map( A1 => n21191, A2 => n15776, B1 => n21612, B2 => 
                           n21183, ZN => n5721);
   U14320 : OAI22_X1 port map( A1 => n21191, A2 => n15775, B1 => n21615, B2 => 
                           n21183, ZN => n5722);
   U14321 : OAI22_X1 port map( A1 => n21191, A2 => n15774, B1 => n21618, B2 => 
                           n21183, ZN => n5723);
   U14322 : OAI22_X1 port map( A1 => n21191, A2 => n15773, B1 => n21621, B2 => 
                           n21183, ZN => n5724);
   U14323 : OAI22_X1 port map( A1 => n21191, A2 => n15772, B1 => n21624, B2 => 
                           n21183, ZN => n5725);
   U14324 : OAI22_X1 port map( A1 => n21191, A2 => n15771, B1 => n21627, B2 => 
                           n21183, ZN => n5726);
   U14325 : OAI22_X1 port map( A1 => n21191, A2 => n15770, B1 => n21630, B2 => 
                           n21183, ZN => n5727);
   U14326 : OAI22_X1 port map( A1 => n21191, A2 => n15769, B1 => n21633, B2 => 
                           n21183, ZN => n5728);
   U14327 : OAI22_X1 port map( A1 => n21191, A2 => n15768, B1 => n21636, B2 => 
                           n21184, ZN => n5729);
   U14328 : OAI22_X1 port map( A1 => n21191, A2 => n15767, B1 => n21639, B2 => 
                           n21184, ZN => n5730);
   U14329 : OAI22_X1 port map( A1 => n21192, A2 => n15766, B1 => n21642, B2 => 
                           n21184, ZN => n5731);
   U14330 : OAI22_X1 port map( A1 => n21192, A2 => n15765, B1 => n21645, B2 => 
                           n21184, ZN => n5732);
   U14331 : OAI22_X1 port map( A1 => n21192, A2 => n15764, B1 => n21648, B2 => 
                           n21184, ZN => n5733);
   U14332 : OAI22_X1 port map( A1 => n21192, A2 => n15763, B1 => n21651, B2 => 
                           n21184, ZN => n5734);
   U14333 : OAI22_X1 port map( A1 => n21192, A2 => n15762, B1 => n21654, B2 => 
                           n21184, ZN => n5735);
   U14334 : OAI22_X1 port map( A1 => n21192, A2 => n15761, B1 => n21657, B2 => 
                           n21184, ZN => n5736);
   U14335 : OAI22_X1 port map( A1 => n21192, A2 => n15760, B1 => n21660, B2 => 
                           n21184, ZN => n5737);
   U14336 : OAI22_X1 port map( A1 => n21192, A2 => n15759, B1 => n21663, B2 => 
                           n21184, ZN => n5738);
   U14337 : OAI22_X1 port map( A1 => n21192, A2 => n15758, B1 => n21666, B2 => 
                           n21184, ZN => n5739);
   U14338 : OAI22_X1 port map( A1 => n21192, A2 => n15757, B1 => n21669, B2 => 
                           n21184, ZN => n5740);
   U14339 : OAI22_X1 port map( A1 => n21192, A2 => n15756, B1 => n21672, B2 => 
                           n21185, ZN => n5741);
   U14340 : OAI22_X1 port map( A1 => n21192, A2 => n15755, B1 => n21675, B2 => 
                           n21185, ZN => n5742);
   U14341 : OAI22_X1 port map( A1 => n21192, A2 => n15754, B1 => n21678, B2 => 
                           n21185, ZN => n5743);
   U14342 : OAI22_X1 port map( A1 => n21193, A2 => n15753, B1 => n21681, B2 => 
                           n21185, ZN => n5744);
   U14343 : OAI22_X1 port map( A1 => n21193, A2 => n15752, B1 => n21684, B2 => 
                           n21185, ZN => n5745);
   U14344 : OAI22_X1 port map( A1 => n21193, A2 => n15751, B1 => n21687, B2 => 
                           n21185, ZN => n5746);
   U14345 : OAI22_X1 port map( A1 => n21193, A2 => n15750, B1 => n21690, B2 => 
                           n21185, ZN => n5747);
   U14346 : OAI22_X1 port map( A1 => n21193, A2 => n15749, B1 => n21693, B2 => 
                           n21185, ZN => n5748);
   U14347 : OAI22_X1 port map( A1 => n21193, A2 => n15748, B1 => n21696, B2 => 
                           n21185, ZN => n5749);
   U14348 : OAI22_X1 port map( A1 => n21193, A2 => n15747, B1 => n21699, B2 => 
                           n21185, ZN => n5750);
   U14349 : OAI22_X1 port map( A1 => n21193, A2 => n15746, B1 => n21702, B2 => 
                           n21185, ZN => n5751);
   U14350 : OAI22_X1 port map( A1 => n21193, A2 => n15745, B1 => n21705, B2 => 
                           n21185, ZN => n5752);
   U14351 : NAND2_X1 port map( A1 => n17315, A2 => n17311, ZN => n16104);
   U14352 : OAI22_X1 port map( A1 => n21215, A2 => n15668, B1 => n21527, B2 => 
                           n21207, ZN => n5821);
   U14353 : OAI22_X1 port map( A1 => n21215, A2 => n15667, B1 => n21530, B2 => 
                           n21207, ZN => n5822);
   U14354 : OAI22_X1 port map( A1 => n21215, A2 => n15666, B1 => n21533, B2 => 
                           n21207, ZN => n5823);
   U14355 : OAI22_X1 port map( A1 => n21215, A2 => n15665, B1 => n21536, B2 => 
                           n21207, ZN => n5824);
   U14356 : OAI22_X1 port map( A1 => n21215, A2 => n15664, B1 => n21539, B2 => 
                           n21207, ZN => n5825);
   U14357 : OAI22_X1 port map( A1 => n21215, A2 => n15663, B1 => n21542, B2 => 
                           n21207, ZN => n5826);
   U14358 : OAI22_X1 port map( A1 => n21215, A2 => n15662, B1 => n21545, B2 => 
                           n21207, ZN => n5827);
   U14359 : OAI22_X1 port map( A1 => n21215, A2 => n15661, B1 => n21548, B2 => 
                           n21207, ZN => n5828);
   U14360 : OAI22_X1 port map( A1 => n21215, A2 => n15660, B1 => n21551, B2 => 
                           n21207, ZN => n5829);
   U14361 : OAI22_X1 port map( A1 => n21215, A2 => n15659, B1 => n21554, B2 => 
                           n21207, ZN => n5830);
   U14362 : OAI22_X1 port map( A1 => n21215, A2 => n15658, B1 => n21557, B2 => 
                           n21207, ZN => n5831);
   U14363 : OAI22_X1 port map( A1 => n21215, A2 => n15657, B1 => n21560, B2 => 
                           n21207, ZN => n5832);
   U14364 : OAI22_X1 port map( A1 => n21216, A2 => n15656, B1 => n21563, B2 => 
                           n21208, ZN => n5833);
   U14365 : OAI22_X1 port map( A1 => n21216, A2 => n15655, B1 => n21566, B2 => 
                           n21208, ZN => n5834);
   U14366 : OAI22_X1 port map( A1 => n21216, A2 => n15654, B1 => n21569, B2 => 
                           n21208, ZN => n5835);
   U14367 : OAI22_X1 port map( A1 => n21216, A2 => n15653, B1 => n21572, B2 => 
                           n21208, ZN => n5836);
   U14368 : OAI22_X1 port map( A1 => n21216, A2 => n15652, B1 => n21575, B2 => 
                           n21208, ZN => n5837);
   U14369 : OAI22_X1 port map( A1 => n21216, A2 => n15651, B1 => n21578, B2 => 
                           n21208, ZN => n5838);
   U14370 : OAI22_X1 port map( A1 => n21216, A2 => n15650, B1 => n21581, B2 => 
                           n21208, ZN => n5839);
   U14371 : OAI22_X1 port map( A1 => n21216, A2 => n15649, B1 => n21584, B2 => 
                           n21208, ZN => n5840);
   U14372 : OAI22_X1 port map( A1 => n21216, A2 => n15648, B1 => n21587, B2 => 
                           n21208, ZN => n5841);
   U14373 : OAI22_X1 port map( A1 => n21216, A2 => n15647, B1 => n21590, B2 => 
                           n21208, ZN => n5842);
   U14374 : OAI22_X1 port map( A1 => n21216, A2 => n15646, B1 => n21593, B2 => 
                           n21208, ZN => n5843);
   U14375 : OAI22_X1 port map( A1 => n21216, A2 => n15645, B1 => n21596, B2 => 
                           n21208, ZN => n5844);
   U14376 : OAI22_X1 port map( A1 => n21216, A2 => n15644, B1 => n21599, B2 => 
                           n21209, ZN => n5845);
   U14377 : OAI22_X1 port map( A1 => n21217, A2 => n15643, B1 => n21602, B2 => 
                           n21209, ZN => n5846);
   U14378 : OAI22_X1 port map( A1 => n21217, A2 => n15642, B1 => n21605, B2 => 
                           n21209, ZN => n5847);
   U14379 : OAI22_X1 port map( A1 => n21217, A2 => n15641, B1 => n21608, B2 => 
                           n21209, ZN => n5848);
   U14380 : OAI22_X1 port map( A1 => n21217, A2 => n15640, B1 => n21611, B2 => 
                           n21209, ZN => n5849);
   U14381 : OAI22_X1 port map( A1 => n21217, A2 => n15639, B1 => n21614, B2 => 
                           n21209, ZN => n5850);
   U14382 : OAI22_X1 port map( A1 => n21217, A2 => n15638, B1 => n21617, B2 => 
                           n21209, ZN => n5851);
   U14383 : OAI22_X1 port map( A1 => n21217, A2 => n15637, B1 => n21620, B2 => 
                           n21209, ZN => n5852);
   U14384 : OAI22_X1 port map( A1 => n21217, A2 => n15636, B1 => n21623, B2 => 
                           n21209, ZN => n5853);
   U14385 : OAI22_X1 port map( A1 => n21217, A2 => n15635, B1 => n21626, B2 => 
                           n21209, ZN => n5854);
   U14386 : OAI22_X1 port map( A1 => n21217, A2 => n15634, B1 => n21629, B2 => 
                           n21209, ZN => n5855);
   U14387 : OAI22_X1 port map( A1 => n21217, A2 => n15633, B1 => n21632, B2 => 
                           n21209, ZN => n5856);
   U14388 : OAI22_X1 port map( A1 => n21217, A2 => n15632, B1 => n21635, B2 => 
                           n21210, ZN => n5857);
   U14389 : OAI22_X1 port map( A1 => n21217, A2 => n15631, B1 => n21638, B2 => 
                           n21210, ZN => n5858);
   U14390 : OAI22_X1 port map( A1 => n21218, A2 => n15630, B1 => n21641, B2 => 
                           n21210, ZN => n5859);
   U14391 : OAI22_X1 port map( A1 => n21218, A2 => n15629, B1 => n21644, B2 => 
                           n21210, ZN => n5860);
   U14392 : OAI22_X1 port map( A1 => n21218, A2 => n15628, B1 => n21647, B2 => 
                           n21210, ZN => n5861);
   U14393 : OAI22_X1 port map( A1 => n21218, A2 => n15627, B1 => n21650, B2 => 
                           n21210, ZN => n5862);
   U14394 : OAI22_X1 port map( A1 => n21218, A2 => n15626, B1 => n21653, B2 => 
                           n21210, ZN => n5863);
   U14395 : OAI22_X1 port map( A1 => n21218, A2 => n15625, B1 => n21656, B2 => 
                           n21210, ZN => n5864);
   U14396 : OAI22_X1 port map( A1 => n21218, A2 => n15624, B1 => n21659, B2 => 
                           n21210, ZN => n5865);
   U14397 : OAI22_X1 port map( A1 => n21218, A2 => n15623, B1 => n21662, B2 => 
                           n21210, ZN => n5866);
   U14398 : OAI22_X1 port map( A1 => n21218, A2 => n15622, B1 => n21665, B2 => 
                           n21210, ZN => n5867);
   U14399 : OAI22_X1 port map( A1 => n21218, A2 => n15621, B1 => n21668, B2 => 
                           n21210, ZN => n5868);
   U14400 : OAI22_X1 port map( A1 => n21218, A2 => n15620, B1 => n21671, B2 => 
                           n21211, ZN => n5869);
   U14401 : OAI22_X1 port map( A1 => n21218, A2 => n15619, B1 => n21674, B2 => 
                           n21211, ZN => n5870);
   U14402 : OAI22_X1 port map( A1 => n21218, A2 => n15618, B1 => n21677, B2 => 
                           n21211, ZN => n5871);
   U14403 : OAI22_X1 port map( A1 => n21219, A2 => n15617, B1 => n21680, B2 => 
                           n21211, ZN => n5872);
   U14404 : OAI22_X1 port map( A1 => n21219, A2 => n15616, B1 => n21683, B2 => 
                           n21211, ZN => n5873);
   U14405 : OAI22_X1 port map( A1 => n21219, A2 => n15615, B1 => n21686, B2 => 
                           n21211, ZN => n5874);
   U14406 : OAI22_X1 port map( A1 => n21219, A2 => n15614, B1 => n21689, B2 => 
                           n21211, ZN => n5875);
   U14407 : OAI22_X1 port map( A1 => n21219, A2 => n15613, B1 => n21692, B2 => 
                           n21211, ZN => n5876);
   U14408 : OAI22_X1 port map( A1 => n21219, A2 => n15612, B1 => n21695, B2 => 
                           n21211, ZN => n5877);
   U14409 : OAI22_X1 port map( A1 => n21219, A2 => n15611, B1 => n21698, B2 => 
                           n21211, ZN => n5878);
   U14410 : OAI22_X1 port map( A1 => n21219, A2 => n15610, B1 => n21701, B2 => 
                           n21211, ZN => n5879);
   U14411 : OAI22_X1 port map( A1 => n21219, A2 => n15609, B1 => n21704, B2 => 
                           n21211, ZN => n5880);
   U14412 : OAI22_X1 port map( A1 => n21254, A2 => n15469, B1 => n21527, B2 => 
                           n21246, ZN => n6013);
   U14413 : OAI22_X1 port map( A1 => n21254, A2 => n15468, B1 => n21530, B2 => 
                           n21246, ZN => n6014);
   U14414 : OAI22_X1 port map( A1 => n21254, A2 => n15467, B1 => n21533, B2 => 
                           n21246, ZN => n6015);
   U14415 : OAI22_X1 port map( A1 => n21254, A2 => n15466, B1 => n21536, B2 => 
                           n21246, ZN => n6016);
   U14416 : OAI22_X1 port map( A1 => n21254, A2 => n15465, B1 => n21539, B2 => 
                           n21246, ZN => n6017);
   U14417 : OAI22_X1 port map( A1 => n21254, A2 => n15464, B1 => n21542, B2 => 
                           n21246, ZN => n6018);
   U14418 : OAI22_X1 port map( A1 => n21254, A2 => n15463, B1 => n21545, B2 => 
                           n21246, ZN => n6019);
   U14419 : OAI22_X1 port map( A1 => n21254, A2 => n15462, B1 => n21548, B2 => 
                           n21246, ZN => n6020);
   U14420 : OAI22_X1 port map( A1 => n21254, A2 => n15461, B1 => n21551, B2 => 
                           n21246, ZN => n6021);
   U14421 : OAI22_X1 port map( A1 => n21254, A2 => n15460, B1 => n21554, B2 => 
                           n21246, ZN => n6022);
   U14422 : OAI22_X1 port map( A1 => n21254, A2 => n15459, B1 => n21557, B2 => 
                           n21246, ZN => n6023);
   U14423 : OAI22_X1 port map( A1 => n21254, A2 => n15458, B1 => n21560, B2 => 
                           n21246, ZN => n6024);
   U14424 : OAI22_X1 port map( A1 => n21255, A2 => n15457, B1 => n21563, B2 => 
                           n21247, ZN => n6025);
   U14425 : OAI22_X1 port map( A1 => n21255, A2 => n15456, B1 => n21566, B2 => 
                           n21247, ZN => n6026);
   U14426 : OAI22_X1 port map( A1 => n21255, A2 => n15455, B1 => n21569, B2 => 
                           n21247, ZN => n6027);
   U14427 : OAI22_X1 port map( A1 => n21255, A2 => n15454, B1 => n21572, B2 => 
                           n21247, ZN => n6028);
   U14428 : OAI22_X1 port map( A1 => n21255, A2 => n15453, B1 => n21575, B2 => 
                           n21247, ZN => n6029);
   U14429 : OAI22_X1 port map( A1 => n21255, A2 => n15452, B1 => n21578, B2 => 
                           n21247, ZN => n6030);
   U14430 : OAI22_X1 port map( A1 => n21255, A2 => n15451, B1 => n21581, B2 => 
                           n21247, ZN => n6031);
   U14431 : OAI22_X1 port map( A1 => n21255, A2 => n15450, B1 => n21584, B2 => 
                           n21247, ZN => n6032);
   U14432 : OAI22_X1 port map( A1 => n21255, A2 => n15449, B1 => n21587, B2 => 
                           n21247, ZN => n6033);
   U14433 : OAI22_X1 port map( A1 => n21255, A2 => n15448, B1 => n21590, B2 => 
                           n21247, ZN => n6034);
   U14434 : OAI22_X1 port map( A1 => n21255, A2 => n15447, B1 => n21593, B2 => 
                           n21247, ZN => n6035);
   U14435 : OAI22_X1 port map( A1 => n21255, A2 => n15446, B1 => n21596, B2 => 
                           n21247, ZN => n6036);
   U14436 : OAI22_X1 port map( A1 => n21255, A2 => n15445, B1 => n21599, B2 => 
                           n21248, ZN => n6037);
   U14437 : OAI22_X1 port map( A1 => n21256, A2 => n15444, B1 => n21602, B2 => 
                           n21248, ZN => n6038);
   U14438 : OAI22_X1 port map( A1 => n21256, A2 => n15443, B1 => n21605, B2 => 
                           n21248, ZN => n6039);
   U14439 : OAI22_X1 port map( A1 => n21256, A2 => n15442, B1 => n21608, B2 => 
                           n21248, ZN => n6040);
   U14440 : OAI22_X1 port map( A1 => n21256, A2 => n15441, B1 => n21611, B2 => 
                           n21248, ZN => n6041);
   U14441 : OAI22_X1 port map( A1 => n21256, A2 => n15440, B1 => n21614, B2 => 
                           n21248, ZN => n6042);
   U14442 : OAI22_X1 port map( A1 => n21256, A2 => n15439, B1 => n21617, B2 => 
                           n21248, ZN => n6043);
   U14443 : OAI22_X1 port map( A1 => n21256, A2 => n15438, B1 => n21620, B2 => 
                           n21248, ZN => n6044);
   U14444 : OAI22_X1 port map( A1 => n21256, A2 => n15437, B1 => n21623, B2 => 
                           n21248, ZN => n6045);
   U14445 : OAI22_X1 port map( A1 => n21256, A2 => n15436, B1 => n21626, B2 => 
                           n21248, ZN => n6046);
   U14446 : OAI22_X1 port map( A1 => n21256, A2 => n15435, B1 => n21629, B2 => 
                           n21248, ZN => n6047);
   U14447 : OAI22_X1 port map( A1 => n21256, A2 => n15434, B1 => n21632, B2 => 
                           n21248, ZN => n6048);
   U14448 : OAI22_X1 port map( A1 => n21256, A2 => n15433, B1 => n21635, B2 => 
                           n21249, ZN => n6049);
   U14449 : OAI22_X1 port map( A1 => n21256, A2 => n15432, B1 => n21638, B2 => 
                           n21249, ZN => n6050);
   U14450 : OAI22_X1 port map( A1 => n21257, A2 => n15431, B1 => n21641, B2 => 
                           n21249, ZN => n6051);
   U14451 : OAI22_X1 port map( A1 => n21257, A2 => n15430, B1 => n21644, B2 => 
                           n21249, ZN => n6052);
   U14452 : OAI22_X1 port map( A1 => n21257, A2 => n15429, B1 => n21647, B2 => 
                           n21249, ZN => n6053);
   U14453 : OAI22_X1 port map( A1 => n21257, A2 => n15428, B1 => n21650, B2 => 
                           n21249, ZN => n6054);
   U14454 : OAI22_X1 port map( A1 => n21257, A2 => n15427, B1 => n21653, B2 => 
                           n21249, ZN => n6055);
   U14455 : OAI22_X1 port map( A1 => n21257, A2 => n15426, B1 => n21656, B2 => 
                           n21249, ZN => n6056);
   U14456 : OAI22_X1 port map( A1 => n21257, A2 => n15425, B1 => n21659, B2 => 
                           n21249, ZN => n6057);
   U14457 : OAI22_X1 port map( A1 => n21257, A2 => n15424, B1 => n21662, B2 => 
                           n21249, ZN => n6058);
   U14458 : OAI22_X1 port map( A1 => n21257, A2 => n15423, B1 => n21665, B2 => 
                           n21249, ZN => n6059);
   U14459 : OAI22_X1 port map( A1 => n21257, A2 => n15422, B1 => n21668, B2 => 
                           n21249, ZN => n6060);
   U14460 : OAI22_X1 port map( A1 => n21257, A2 => n15421, B1 => n21671, B2 => 
                           n21250, ZN => n6061);
   U14461 : OAI22_X1 port map( A1 => n21257, A2 => n15420, B1 => n21674, B2 => 
                           n21250, ZN => n6062);
   U14462 : OAI22_X1 port map( A1 => n21257, A2 => n15419, B1 => n21677, B2 => 
                           n21250, ZN => n6063);
   U14463 : OAI22_X1 port map( A1 => n21258, A2 => n15418, B1 => n21680, B2 => 
                           n21250, ZN => n6064);
   U14464 : OAI22_X1 port map( A1 => n21258, A2 => n15417, B1 => n21683, B2 => 
                           n21250, ZN => n6065);
   U14465 : OAI22_X1 port map( A1 => n21258, A2 => n15416, B1 => n21686, B2 => 
                           n21250, ZN => n6066);
   U14466 : OAI22_X1 port map( A1 => n21258, A2 => n15415, B1 => n21689, B2 => 
                           n21250, ZN => n6067);
   U14467 : OAI22_X1 port map( A1 => n21258, A2 => n15414, B1 => n21692, B2 => 
                           n21250, ZN => n6068);
   U14468 : OAI22_X1 port map( A1 => n21258, A2 => n15413, B1 => n21695, B2 => 
                           n21250, ZN => n6069);
   U14469 : OAI22_X1 port map( A1 => n21258, A2 => n15412, B1 => n21698, B2 => 
                           n21250, ZN => n6070);
   U14470 : OAI22_X1 port map( A1 => n21258, A2 => n15411, B1 => n21701, B2 => 
                           n21250, ZN => n6071);
   U14471 : OAI22_X1 port map( A1 => n21258, A2 => n15410, B1 => n21704, B2 => 
                           n21250, ZN => n6072);
   U14472 : OAI22_X1 port map( A1 => n21280, A2 => n15337, B1 => n21527, B2 => 
                           n21272, ZN => n6141);
   U14473 : OAI22_X1 port map( A1 => n21280, A2 => n15336, B1 => n21530, B2 => 
                           n21272, ZN => n6142);
   U14474 : OAI22_X1 port map( A1 => n21280, A2 => n15335, B1 => n21533, B2 => 
                           n21272, ZN => n6143);
   U14475 : OAI22_X1 port map( A1 => n21280, A2 => n15334, B1 => n21536, B2 => 
                           n21272, ZN => n6144);
   U14476 : OAI22_X1 port map( A1 => n21280, A2 => n15333, B1 => n21539, B2 => 
                           n21272, ZN => n6145);
   U14477 : OAI22_X1 port map( A1 => n21280, A2 => n15332, B1 => n21542, B2 => 
                           n21272, ZN => n6146);
   U14478 : OAI22_X1 port map( A1 => n21280, A2 => n15331, B1 => n21545, B2 => 
                           n21272, ZN => n6147);
   U14479 : OAI22_X1 port map( A1 => n21280, A2 => n15330, B1 => n21548, B2 => 
                           n21272, ZN => n6148);
   U14480 : OAI22_X1 port map( A1 => n21280, A2 => n15329, B1 => n21551, B2 => 
                           n21272, ZN => n6149);
   U14481 : OAI22_X1 port map( A1 => n21280, A2 => n15328, B1 => n21554, B2 => 
                           n21272, ZN => n6150);
   U14482 : OAI22_X1 port map( A1 => n21280, A2 => n15327, B1 => n21557, B2 => 
                           n21272, ZN => n6151);
   U14483 : OAI22_X1 port map( A1 => n21280, A2 => n15326, B1 => n21560, B2 => 
                           n21272, ZN => n6152);
   U14484 : OAI22_X1 port map( A1 => n21281, A2 => n15325, B1 => n21563, B2 => 
                           n21273, ZN => n6153);
   U14485 : OAI22_X1 port map( A1 => n21281, A2 => n15324, B1 => n21566, B2 => 
                           n21273, ZN => n6154);
   U14486 : OAI22_X1 port map( A1 => n21281, A2 => n15323, B1 => n21569, B2 => 
                           n21273, ZN => n6155);
   U14487 : OAI22_X1 port map( A1 => n21281, A2 => n15322, B1 => n21572, B2 => 
                           n21273, ZN => n6156);
   U14488 : OAI22_X1 port map( A1 => n21281, A2 => n15321, B1 => n21575, B2 => 
                           n21273, ZN => n6157);
   U14489 : OAI22_X1 port map( A1 => n21281, A2 => n15320, B1 => n21578, B2 => 
                           n21273, ZN => n6158);
   U14490 : OAI22_X1 port map( A1 => n21281, A2 => n15319, B1 => n21581, B2 => 
                           n21273, ZN => n6159);
   U14491 : OAI22_X1 port map( A1 => n21281, A2 => n15318, B1 => n21584, B2 => 
                           n21273, ZN => n6160);
   U14492 : OAI22_X1 port map( A1 => n21281, A2 => n15317, B1 => n21587, B2 => 
                           n21273, ZN => n6161);
   U14493 : OAI22_X1 port map( A1 => n21281, A2 => n15316, B1 => n21590, B2 => 
                           n21273, ZN => n6162);
   U14494 : OAI22_X1 port map( A1 => n21281, A2 => n15315, B1 => n21593, B2 => 
                           n21273, ZN => n6163);
   U14495 : OAI22_X1 port map( A1 => n21281, A2 => n15314, B1 => n21596, B2 => 
                           n21273, ZN => n6164);
   U14496 : OAI22_X1 port map( A1 => n21281, A2 => n15313, B1 => n21599, B2 => 
                           n21274, ZN => n6165);
   U14497 : OAI22_X1 port map( A1 => n21282, A2 => n15312, B1 => n21602, B2 => 
                           n21274, ZN => n6166);
   U14498 : OAI22_X1 port map( A1 => n21282, A2 => n15311, B1 => n21605, B2 => 
                           n21274, ZN => n6167);
   U14499 : OAI22_X1 port map( A1 => n21282, A2 => n15310, B1 => n21608, B2 => 
                           n21274, ZN => n6168);
   U14500 : OAI22_X1 port map( A1 => n21282, A2 => n15309, B1 => n21611, B2 => 
                           n21274, ZN => n6169);
   U14501 : OAI22_X1 port map( A1 => n21282, A2 => n15308, B1 => n21614, B2 => 
                           n21274, ZN => n6170);
   U14502 : OAI22_X1 port map( A1 => n21282, A2 => n15307, B1 => n21617, B2 => 
                           n21274, ZN => n6171);
   U14503 : OAI22_X1 port map( A1 => n21282, A2 => n15306, B1 => n21620, B2 => 
                           n21274, ZN => n6172);
   U14504 : OAI22_X1 port map( A1 => n21282, A2 => n15305, B1 => n21623, B2 => 
                           n21274, ZN => n6173);
   U14505 : OAI22_X1 port map( A1 => n21282, A2 => n15304, B1 => n21626, B2 => 
                           n21274, ZN => n6174);
   U14506 : OAI22_X1 port map( A1 => n21282, A2 => n15303, B1 => n21629, B2 => 
                           n21274, ZN => n6175);
   U14507 : OAI22_X1 port map( A1 => n21282, A2 => n15302, B1 => n21632, B2 => 
                           n21274, ZN => n6176);
   U14508 : OAI22_X1 port map( A1 => n21282, A2 => n15301, B1 => n21635, B2 => 
                           n21275, ZN => n6177);
   U14509 : OAI22_X1 port map( A1 => n21282, A2 => n15300, B1 => n21638, B2 => 
                           n21275, ZN => n6178);
   U14510 : OAI22_X1 port map( A1 => n21283, A2 => n15299, B1 => n21641, B2 => 
                           n21275, ZN => n6179);
   U14511 : OAI22_X1 port map( A1 => n21283, A2 => n15298, B1 => n21644, B2 => 
                           n21275, ZN => n6180);
   U14512 : OAI22_X1 port map( A1 => n21283, A2 => n15297, B1 => n21647, B2 => 
                           n21275, ZN => n6181);
   U14513 : OAI22_X1 port map( A1 => n21283, A2 => n15296, B1 => n21650, B2 => 
                           n21275, ZN => n6182);
   U14514 : OAI22_X1 port map( A1 => n21283, A2 => n15295, B1 => n21653, B2 => 
                           n21275, ZN => n6183);
   U14515 : OAI22_X1 port map( A1 => n21283, A2 => n15294, B1 => n21656, B2 => 
                           n21275, ZN => n6184);
   U14516 : OAI22_X1 port map( A1 => n21283, A2 => n15293, B1 => n21659, B2 => 
                           n21275, ZN => n6185);
   U14517 : OAI22_X1 port map( A1 => n21283, A2 => n15292, B1 => n21662, B2 => 
                           n21275, ZN => n6186);
   U14518 : OAI22_X1 port map( A1 => n21283, A2 => n15291, B1 => n21665, B2 => 
                           n21275, ZN => n6187);
   U14519 : OAI22_X1 port map( A1 => n21283, A2 => n15290, B1 => n21668, B2 => 
                           n21275, ZN => n6188);
   U14520 : OAI22_X1 port map( A1 => n21283, A2 => n15289, B1 => n21671, B2 => 
                           n21276, ZN => n6189);
   U14521 : OAI22_X1 port map( A1 => n21283, A2 => n15288, B1 => n21674, B2 => 
                           n21276, ZN => n6190);
   U14522 : OAI22_X1 port map( A1 => n21283, A2 => n15287, B1 => n21677, B2 => 
                           n21276, ZN => n6191);
   U14523 : OAI22_X1 port map( A1 => n21284, A2 => n15286, B1 => n21680, B2 => 
                           n21276, ZN => n6192);
   U14524 : OAI22_X1 port map( A1 => n21284, A2 => n15285, B1 => n21683, B2 => 
                           n21276, ZN => n6193);
   U14525 : OAI22_X1 port map( A1 => n21284, A2 => n15284, B1 => n21686, B2 => 
                           n21276, ZN => n6194);
   U14526 : OAI22_X1 port map( A1 => n21284, A2 => n15283, B1 => n21689, B2 => 
                           n21276, ZN => n6195);
   U14527 : OAI22_X1 port map( A1 => n21284, A2 => n15282, B1 => n21692, B2 => 
                           n21276, ZN => n6196);
   U14528 : OAI22_X1 port map( A1 => n21284, A2 => n15281, B1 => n21695, B2 => 
                           n21276, ZN => n6197);
   U14529 : OAI22_X1 port map( A1 => n21284, A2 => n15280, B1 => n21698, B2 => 
                           n21276, ZN => n6198);
   U14530 : OAI22_X1 port map( A1 => n21284, A2 => n15279, B1 => n21701, B2 => 
                           n21276, ZN => n6199);
   U14531 : OAI22_X1 port map( A1 => n21284, A2 => n15278, B1 => n21704, B2 => 
                           n21276, ZN => n6200);
   U14532 : OAI22_X1 port map( A1 => n21332, A2 => n15070, B1 => n21527, B2 => 
                           n21324, ZN => n6397);
   U14533 : OAI22_X1 port map( A1 => n21332, A2 => n15069, B1 => n21530, B2 => 
                           n21324, ZN => n6398);
   U14534 : OAI22_X1 port map( A1 => n21332, A2 => n15068, B1 => n21533, B2 => 
                           n21324, ZN => n6399);
   U14535 : OAI22_X1 port map( A1 => n21332, A2 => n15067, B1 => n21536, B2 => 
                           n21324, ZN => n6400);
   U14536 : OAI22_X1 port map( A1 => n21332, A2 => n15066, B1 => n21539, B2 => 
                           n21324, ZN => n6401);
   U14537 : OAI22_X1 port map( A1 => n21332, A2 => n15065, B1 => n21542, B2 => 
                           n21324, ZN => n6402);
   U14538 : OAI22_X1 port map( A1 => n21332, A2 => n15064, B1 => n21545, B2 => 
                           n21324, ZN => n6403);
   U14539 : OAI22_X1 port map( A1 => n21332, A2 => n15063, B1 => n21548, B2 => 
                           n21324, ZN => n6404);
   U14540 : OAI22_X1 port map( A1 => n21332, A2 => n15062, B1 => n21551, B2 => 
                           n21324, ZN => n6405);
   U14541 : OAI22_X1 port map( A1 => n21332, A2 => n15061, B1 => n21554, B2 => 
                           n21324, ZN => n6406);
   U14542 : OAI22_X1 port map( A1 => n21332, A2 => n15060, B1 => n21557, B2 => 
                           n21324, ZN => n6407);
   U14543 : OAI22_X1 port map( A1 => n21332, A2 => n15059, B1 => n21560, B2 => 
                           n21324, ZN => n6408);
   U14544 : OAI22_X1 port map( A1 => n21333, A2 => n15058, B1 => n21563, B2 => 
                           n21325, ZN => n6409);
   U14545 : OAI22_X1 port map( A1 => n21333, A2 => n15057, B1 => n21566, B2 => 
                           n21325, ZN => n6410);
   U14546 : OAI22_X1 port map( A1 => n21333, A2 => n15056, B1 => n21569, B2 => 
                           n21325, ZN => n6411);
   U14547 : OAI22_X1 port map( A1 => n21333, A2 => n15055, B1 => n21572, B2 => 
                           n21325, ZN => n6412);
   U14548 : OAI22_X1 port map( A1 => n21333, A2 => n15054, B1 => n21575, B2 => 
                           n21325, ZN => n6413);
   U14549 : OAI22_X1 port map( A1 => n21333, A2 => n15053, B1 => n21578, B2 => 
                           n21325, ZN => n6414);
   U14550 : OAI22_X1 port map( A1 => n21333, A2 => n15052, B1 => n21581, B2 => 
                           n21325, ZN => n6415);
   U14551 : OAI22_X1 port map( A1 => n21333, A2 => n15051, B1 => n21584, B2 => 
                           n21325, ZN => n6416);
   U14552 : OAI22_X1 port map( A1 => n21333, A2 => n15050, B1 => n21587, B2 => 
                           n21325, ZN => n6417);
   U14553 : OAI22_X1 port map( A1 => n21333, A2 => n15049, B1 => n21590, B2 => 
                           n21325, ZN => n6418);
   U14554 : OAI22_X1 port map( A1 => n21333, A2 => n15048, B1 => n21593, B2 => 
                           n21325, ZN => n6419);
   U14555 : OAI22_X1 port map( A1 => n21333, A2 => n15047, B1 => n21596, B2 => 
                           n21325, ZN => n6420);
   U14556 : OAI22_X1 port map( A1 => n21333, A2 => n15046, B1 => n21599, B2 => 
                           n21326, ZN => n6421);
   U14557 : OAI22_X1 port map( A1 => n21334, A2 => n15045, B1 => n21602, B2 => 
                           n21326, ZN => n6422);
   U14558 : OAI22_X1 port map( A1 => n21334, A2 => n15044, B1 => n21605, B2 => 
                           n21326, ZN => n6423);
   U14559 : OAI22_X1 port map( A1 => n21334, A2 => n15043, B1 => n21608, B2 => 
                           n21326, ZN => n6424);
   U14560 : OAI22_X1 port map( A1 => n21334, A2 => n15042, B1 => n21611, B2 => 
                           n21326, ZN => n6425);
   U14561 : OAI22_X1 port map( A1 => n21334, A2 => n15041, B1 => n21614, B2 => 
                           n21326, ZN => n6426);
   U14562 : OAI22_X1 port map( A1 => n21334, A2 => n15040, B1 => n21617, B2 => 
                           n21326, ZN => n6427);
   U14563 : OAI22_X1 port map( A1 => n21334, A2 => n15039, B1 => n21620, B2 => 
                           n21326, ZN => n6428);
   U14564 : OAI22_X1 port map( A1 => n21334, A2 => n15038, B1 => n21623, B2 => 
                           n21326, ZN => n6429);
   U14565 : OAI22_X1 port map( A1 => n21334, A2 => n15037, B1 => n21626, B2 => 
                           n21326, ZN => n6430);
   U14566 : OAI22_X1 port map( A1 => n21334, A2 => n15036, B1 => n21629, B2 => 
                           n21326, ZN => n6431);
   U14567 : OAI22_X1 port map( A1 => n21334, A2 => n15035, B1 => n21632, B2 => 
                           n21326, ZN => n6432);
   U14568 : OAI22_X1 port map( A1 => n21334, A2 => n15034, B1 => n21635, B2 => 
                           n21327, ZN => n6433);
   U14569 : OAI22_X1 port map( A1 => n21334, A2 => n15033, B1 => n21638, B2 => 
                           n21327, ZN => n6434);
   U14570 : OAI22_X1 port map( A1 => n21335, A2 => n15032, B1 => n21641, B2 => 
                           n21327, ZN => n6435);
   U14571 : OAI22_X1 port map( A1 => n21335, A2 => n15031, B1 => n21644, B2 => 
                           n21327, ZN => n6436);
   U14572 : OAI22_X1 port map( A1 => n21335, A2 => n15030, B1 => n21647, B2 => 
                           n21327, ZN => n6437);
   U14573 : OAI22_X1 port map( A1 => n21335, A2 => n15029, B1 => n21650, B2 => 
                           n21327, ZN => n6438);
   U14574 : OAI22_X1 port map( A1 => n21335, A2 => n15028, B1 => n21653, B2 => 
                           n21327, ZN => n6439);
   U14575 : OAI22_X1 port map( A1 => n21335, A2 => n15027, B1 => n21656, B2 => 
                           n21327, ZN => n6440);
   U14576 : OAI22_X1 port map( A1 => n21335, A2 => n15026, B1 => n21659, B2 => 
                           n21327, ZN => n6441);
   U14577 : OAI22_X1 port map( A1 => n21335, A2 => n15025, B1 => n21662, B2 => 
                           n21327, ZN => n6442);
   U14578 : OAI22_X1 port map( A1 => n21335, A2 => n15024, B1 => n21665, B2 => 
                           n21327, ZN => n6443);
   U14579 : OAI22_X1 port map( A1 => n21335, A2 => n15023, B1 => n21668, B2 => 
                           n21327, ZN => n6444);
   U14580 : OAI22_X1 port map( A1 => n21335, A2 => n15022, B1 => n21671, B2 => 
                           n21328, ZN => n6445);
   U14581 : OAI22_X1 port map( A1 => n21335, A2 => n15021, B1 => n21674, B2 => 
                           n21328, ZN => n6446);
   U14582 : OAI22_X1 port map( A1 => n21335, A2 => n15020, B1 => n21677, B2 => 
                           n21328, ZN => n6447);
   U14583 : OAI22_X1 port map( A1 => n21336, A2 => n15019, B1 => n21680, B2 => 
                           n21328, ZN => n6448);
   U14584 : OAI22_X1 port map( A1 => n21336, A2 => n15018, B1 => n21683, B2 => 
                           n21328, ZN => n6449);
   U14585 : OAI22_X1 port map( A1 => n21336, A2 => n15017, B1 => n21686, B2 => 
                           n21328, ZN => n6450);
   U14586 : OAI22_X1 port map( A1 => n21336, A2 => n15016, B1 => n21689, B2 => 
                           n21328, ZN => n6451);
   U14587 : OAI22_X1 port map( A1 => n21336, A2 => n15015, B1 => n21692, B2 => 
                           n21328, ZN => n6452);
   U14588 : OAI22_X1 port map( A1 => n21336, A2 => n15014, B1 => n21695, B2 => 
                           n21328, ZN => n6453);
   U14589 : OAI22_X1 port map( A1 => n21336, A2 => n15013, B1 => n21698, B2 => 
                           n21328, ZN => n6454);
   U14590 : OAI22_X1 port map( A1 => n21336, A2 => n15012, B1 => n21701, B2 => 
                           n21328, ZN => n6455);
   U14591 : OAI22_X1 port map( A1 => n21336, A2 => n15011, B1 => n21704, B2 => 
                           n21328, ZN => n6456);
   U14592 : OAI22_X1 port map( A1 => n21345, A2 => n15004, B1 => n21527, B2 => 
                           n21337, ZN => n6461);
   U14593 : OAI22_X1 port map( A1 => n21345, A2 => n15003, B1 => n21530, B2 => 
                           n21337, ZN => n6462);
   U14594 : OAI22_X1 port map( A1 => n21345, A2 => n15002, B1 => n21533, B2 => 
                           n21337, ZN => n6463);
   U14595 : OAI22_X1 port map( A1 => n21345, A2 => n15001, B1 => n21536, B2 => 
                           n21337, ZN => n6464);
   U14596 : OAI22_X1 port map( A1 => n21345, A2 => n15000, B1 => n21539, B2 => 
                           n21337, ZN => n6465);
   U14597 : OAI22_X1 port map( A1 => n21345, A2 => n14999, B1 => n21542, B2 => 
                           n21337, ZN => n6466);
   U14598 : OAI22_X1 port map( A1 => n21345, A2 => n14998, B1 => n21545, B2 => 
                           n21337, ZN => n6467);
   U14599 : OAI22_X1 port map( A1 => n21345, A2 => n14997, B1 => n21548, B2 => 
                           n21337, ZN => n6468);
   U14600 : OAI22_X1 port map( A1 => n21345, A2 => n14996, B1 => n21551, B2 => 
                           n21337, ZN => n6469);
   U14601 : OAI22_X1 port map( A1 => n21345, A2 => n14995, B1 => n21554, B2 => 
                           n21337, ZN => n6470);
   U14602 : OAI22_X1 port map( A1 => n21345, A2 => n14994, B1 => n21557, B2 => 
                           n21337, ZN => n6471);
   U14603 : OAI22_X1 port map( A1 => n21345, A2 => n14993, B1 => n21560, B2 => 
                           n21337, ZN => n6472);
   U14604 : OAI22_X1 port map( A1 => n21346, A2 => n14992, B1 => n21563, B2 => 
                           n21338, ZN => n6473);
   U14605 : OAI22_X1 port map( A1 => n21346, A2 => n14991, B1 => n21566, B2 => 
                           n21338, ZN => n6474);
   U14606 : OAI22_X1 port map( A1 => n21346, A2 => n14990, B1 => n21569, B2 => 
                           n21338, ZN => n6475);
   U14607 : OAI22_X1 port map( A1 => n21346, A2 => n14989, B1 => n21572, B2 => 
                           n21338, ZN => n6476);
   U14608 : OAI22_X1 port map( A1 => n21346, A2 => n14988, B1 => n21575, B2 => 
                           n21338, ZN => n6477);
   U14609 : OAI22_X1 port map( A1 => n21346, A2 => n14987, B1 => n21578, B2 => 
                           n21338, ZN => n6478);
   U14610 : OAI22_X1 port map( A1 => n21346, A2 => n14986, B1 => n21581, B2 => 
                           n21338, ZN => n6479);
   U14611 : OAI22_X1 port map( A1 => n21346, A2 => n14985, B1 => n21584, B2 => 
                           n21338, ZN => n6480);
   U14612 : OAI22_X1 port map( A1 => n21346, A2 => n14984, B1 => n21587, B2 => 
                           n21338, ZN => n6481);
   U14613 : OAI22_X1 port map( A1 => n21346, A2 => n14983, B1 => n21590, B2 => 
                           n21338, ZN => n6482);
   U14614 : OAI22_X1 port map( A1 => n21346, A2 => n14982, B1 => n21593, B2 => 
                           n21338, ZN => n6483);
   U14615 : OAI22_X1 port map( A1 => n21346, A2 => n14981, B1 => n21596, B2 => 
                           n21338, ZN => n6484);
   U14616 : OAI22_X1 port map( A1 => n21346, A2 => n14980, B1 => n21599, B2 => 
                           n21339, ZN => n6485);
   U14617 : OAI22_X1 port map( A1 => n21347, A2 => n14979, B1 => n21602, B2 => 
                           n21339, ZN => n6486);
   U14618 : OAI22_X1 port map( A1 => n21347, A2 => n14978, B1 => n21605, B2 => 
                           n21339, ZN => n6487);
   U14619 : OAI22_X1 port map( A1 => n21347, A2 => n14977, B1 => n21608, B2 => 
                           n21339, ZN => n6488);
   U14620 : OAI22_X1 port map( A1 => n21347, A2 => n14976, B1 => n21611, B2 => 
                           n21339, ZN => n6489);
   U14621 : OAI22_X1 port map( A1 => n21347, A2 => n14975, B1 => n21614, B2 => 
                           n21339, ZN => n6490);
   U14622 : OAI22_X1 port map( A1 => n21347, A2 => n14974, B1 => n21617, B2 => 
                           n21339, ZN => n6491);
   U14623 : OAI22_X1 port map( A1 => n21347, A2 => n14973, B1 => n21620, B2 => 
                           n21339, ZN => n6492);
   U14624 : OAI22_X1 port map( A1 => n21347, A2 => n14972, B1 => n21623, B2 => 
                           n21339, ZN => n6493);
   U14625 : OAI22_X1 port map( A1 => n21347, A2 => n14971, B1 => n21626, B2 => 
                           n21339, ZN => n6494);
   U14626 : OAI22_X1 port map( A1 => n21347, A2 => n14970, B1 => n21629, B2 => 
                           n21339, ZN => n6495);
   U14627 : OAI22_X1 port map( A1 => n21347, A2 => n14969, B1 => n21632, B2 => 
                           n21339, ZN => n6496);
   U14628 : OAI22_X1 port map( A1 => n21347, A2 => n14968, B1 => n21635, B2 => 
                           n21340, ZN => n6497);
   U14629 : OAI22_X1 port map( A1 => n21347, A2 => n14967, B1 => n21638, B2 => 
                           n21340, ZN => n6498);
   U14630 : OAI22_X1 port map( A1 => n21348, A2 => n14966, B1 => n21641, B2 => 
                           n21340, ZN => n6499);
   U14631 : OAI22_X1 port map( A1 => n21348, A2 => n14965, B1 => n21644, B2 => 
                           n21340, ZN => n6500);
   U14632 : OAI22_X1 port map( A1 => n21348, A2 => n14964, B1 => n21647, B2 => 
                           n21340, ZN => n6501);
   U14633 : OAI22_X1 port map( A1 => n21348, A2 => n14963, B1 => n21650, B2 => 
                           n21340, ZN => n6502);
   U14634 : OAI22_X1 port map( A1 => n21348, A2 => n14962, B1 => n21653, B2 => 
                           n21340, ZN => n6503);
   U14635 : OAI22_X1 port map( A1 => n21348, A2 => n14961, B1 => n21656, B2 => 
                           n21340, ZN => n6504);
   U14636 : OAI22_X1 port map( A1 => n21348, A2 => n14960, B1 => n21659, B2 => 
                           n21340, ZN => n6505);
   U14637 : OAI22_X1 port map( A1 => n21348, A2 => n14959, B1 => n21662, B2 => 
                           n21340, ZN => n6506);
   U14638 : OAI22_X1 port map( A1 => n21348, A2 => n14958, B1 => n21665, B2 => 
                           n21340, ZN => n6507);
   U14639 : OAI22_X1 port map( A1 => n21348, A2 => n14957, B1 => n21668, B2 => 
                           n21340, ZN => n6508);
   U14640 : OAI22_X1 port map( A1 => n21348, A2 => n14956, B1 => n21671, B2 => 
                           n21341, ZN => n6509);
   U14641 : OAI22_X1 port map( A1 => n21348, A2 => n14955, B1 => n21674, B2 => 
                           n21341, ZN => n6510);
   U14642 : OAI22_X1 port map( A1 => n21348, A2 => n14954, B1 => n21677, B2 => 
                           n21341, ZN => n6511);
   U14643 : OAI22_X1 port map( A1 => n21349, A2 => n14953, B1 => n21680, B2 => 
                           n21341, ZN => n6512);
   U14644 : OAI22_X1 port map( A1 => n21349, A2 => n14952, B1 => n21683, B2 => 
                           n21341, ZN => n6513);
   U14645 : OAI22_X1 port map( A1 => n21349, A2 => n14951, B1 => n21686, B2 => 
                           n21341, ZN => n6514);
   U14646 : OAI22_X1 port map( A1 => n21349, A2 => n14950, B1 => n21689, B2 => 
                           n21341, ZN => n6515);
   U14647 : OAI22_X1 port map( A1 => n21349, A2 => n14949, B1 => n21692, B2 => 
                           n21341, ZN => n6516);
   U14648 : OAI22_X1 port map( A1 => n21349, A2 => n14948, B1 => n21695, B2 => 
                           n21341, ZN => n6517);
   U14649 : OAI22_X1 port map( A1 => n21349, A2 => n14947, B1 => n21698, B2 => 
                           n21341, ZN => n6518);
   U14650 : OAI22_X1 port map( A1 => n21349, A2 => n14946, B1 => n21701, B2 => 
                           n21341, ZN => n6519);
   U14651 : OAI22_X1 port map( A1 => n21349, A2 => n14945, B1 => n21704, B2 => 
                           n21341, ZN => n6520);
   U14652 : OAI22_X1 port map( A1 => n21358, A2 => n14938, B1 => n21527, B2 => 
                           n21350, ZN => n6525);
   U14653 : OAI22_X1 port map( A1 => n21358, A2 => n14937, B1 => n21530, B2 => 
                           n21350, ZN => n6526);
   U14654 : OAI22_X1 port map( A1 => n21358, A2 => n14936, B1 => n21533, B2 => 
                           n21350, ZN => n6527);
   U14655 : OAI22_X1 port map( A1 => n21358, A2 => n14935, B1 => n21536, B2 => 
                           n21350, ZN => n6528);
   U14656 : OAI22_X1 port map( A1 => n21358, A2 => n14934, B1 => n21539, B2 => 
                           n21350, ZN => n6529);
   U14657 : OAI22_X1 port map( A1 => n21358, A2 => n14933, B1 => n21542, B2 => 
                           n21350, ZN => n6530);
   U14658 : OAI22_X1 port map( A1 => n21358, A2 => n14932, B1 => n21545, B2 => 
                           n21350, ZN => n6531);
   U14659 : OAI22_X1 port map( A1 => n21358, A2 => n14931, B1 => n21548, B2 => 
                           n21350, ZN => n6532);
   U14660 : OAI22_X1 port map( A1 => n21358, A2 => n14930, B1 => n21551, B2 => 
                           n21350, ZN => n6533);
   U14661 : OAI22_X1 port map( A1 => n21358, A2 => n14929, B1 => n21554, B2 => 
                           n21350, ZN => n6534);
   U14662 : OAI22_X1 port map( A1 => n21358, A2 => n14928, B1 => n21557, B2 => 
                           n21350, ZN => n6535);
   U14663 : OAI22_X1 port map( A1 => n21358, A2 => n14927, B1 => n21560, B2 => 
                           n21350, ZN => n6536);
   U14664 : OAI22_X1 port map( A1 => n21359, A2 => n14926, B1 => n21563, B2 => 
                           n21351, ZN => n6537);
   U14665 : OAI22_X1 port map( A1 => n21359, A2 => n14925, B1 => n21566, B2 => 
                           n21351, ZN => n6538);
   U14666 : OAI22_X1 port map( A1 => n21359, A2 => n14924, B1 => n21569, B2 => 
                           n21351, ZN => n6539);
   U14667 : OAI22_X1 port map( A1 => n21359, A2 => n14923, B1 => n21572, B2 => 
                           n21351, ZN => n6540);
   U14668 : OAI22_X1 port map( A1 => n21359, A2 => n14922, B1 => n21575, B2 => 
                           n21351, ZN => n6541);
   U14669 : OAI22_X1 port map( A1 => n21359, A2 => n14921, B1 => n21578, B2 => 
                           n21351, ZN => n6542);
   U14670 : OAI22_X1 port map( A1 => n21359, A2 => n14920, B1 => n21581, B2 => 
                           n21351, ZN => n6543);
   U14671 : OAI22_X1 port map( A1 => n21359, A2 => n14919, B1 => n21584, B2 => 
                           n21351, ZN => n6544);
   U14672 : OAI22_X1 port map( A1 => n21359, A2 => n14918, B1 => n21587, B2 => 
                           n21351, ZN => n6545);
   U14673 : OAI22_X1 port map( A1 => n21359, A2 => n14917, B1 => n21590, B2 => 
                           n21351, ZN => n6546);
   U14674 : OAI22_X1 port map( A1 => n21359, A2 => n14916, B1 => n21593, B2 => 
                           n21351, ZN => n6547);
   U14675 : OAI22_X1 port map( A1 => n21359, A2 => n14915, B1 => n21596, B2 => 
                           n21351, ZN => n6548);
   U14676 : OAI22_X1 port map( A1 => n21359, A2 => n14914, B1 => n21599, B2 => 
                           n21352, ZN => n6549);
   U14677 : OAI22_X1 port map( A1 => n21360, A2 => n14913, B1 => n21602, B2 => 
                           n21352, ZN => n6550);
   U14678 : OAI22_X1 port map( A1 => n21360, A2 => n14912, B1 => n21605, B2 => 
                           n21352, ZN => n6551);
   U14679 : OAI22_X1 port map( A1 => n21360, A2 => n14911, B1 => n21608, B2 => 
                           n21352, ZN => n6552);
   U14680 : OAI22_X1 port map( A1 => n21360, A2 => n14910, B1 => n21611, B2 => 
                           n21352, ZN => n6553);
   U14681 : OAI22_X1 port map( A1 => n21360, A2 => n14909, B1 => n21614, B2 => 
                           n21352, ZN => n6554);
   U14682 : OAI22_X1 port map( A1 => n21360, A2 => n14908, B1 => n21617, B2 => 
                           n21352, ZN => n6555);
   U14683 : OAI22_X1 port map( A1 => n21360, A2 => n14907, B1 => n21620, B2 => 
                           n21352, ZN => n6556);
   U14684 : OAI22_X1 port map( A1 => n21360, A2 => n14906, B1 => n21623, B2 => 
                           n21352, ZN => n6557);
   U14685 : OAI22_X1 port map( A1 => n21360, A2 => n14905, B1 => n21626, B2 => 
                           n21352, ZN => n6558);
   U14686 : OAI22_X1 port map( A1 => n21360, A2 => n14904, B1 => n21629, B2 => 
                           n21352, ZN => n6559);
   U14687 : OAI22_X1 port map( A1 => n21360, A2 => n14903, B1 => n21632, B2 => 
                           n21352, ZN => n6560);
   U14688 : OAI22_X1 port map( A1 => n21360, A2 => n14902, B1 => n21635, B2 => 
                           n21353, ZN => n6561);
   U14689 : OAI22_X1 port map( A1 => n21360, A2 => n14901, B1 => n21638, B2 => 
                           n21353, ZN => n6562);
   U14690 : OAI22_X1 port map( A1 => n21361, A2 => n14900, B1 => n21641, B2 => 
                           n21353, ZN => n6563);
   U14691 : OAI22_X1 port map( A1 => n21361, A2 => n14899, B1 => n21644, B2 => 
                           n21353, ZN => n6564);
   U14692 : OAI22_X1 port map( A1 => n21361, A2 => n14898, B1 => n21647, B2 => 
                           n21353, ZN => n6565);
   U14693 : OAI22_X1 port map( A1 => n21361, A2 => n14897, B1 => n21650, B2 => 
                           n21353, ZN => n6566);
   U14694 : OAI22_X1 port map( A1 => n21361, A2 => n14896, B1 => n21653, B2 => 
                           n21353, ZN => n6567);
   U14695 : OAI22_X1 port map( A1 => n21361, A2 => n14895, B1 => n21656, B2 => 
                           n21353, ZN => n6568);
   U14696 : OAI22_X1 port map( A1 => n21361, A2 => n14894, B1 => n21659, B2 => 
                           n21353, ZN => n6569);
   U14697 : OAI22_X1 port map( A1 => n21361, A2 => n14893, B1 => n21662, B2 => 
                           n21353, ZN => n6570);
   U14698 : OAI22_X1 port map( A1 => n21361, A2 => n14892, B1 => n21665, B2 => 
                           n21353, ZN => n6571);
   U14699 : OAI22_X1 port map( A1 => n21361, A2 => n14891, B1 => n21668, B2 => 
                           n21353, ZN => n6572);
   U14700 : OAI22_X1 port map( A1 => n21361, A2 => n14890, B1 => n21671, B2 => 
                           n21354, ZN => n6573);
   U14701 : OAI22_X1 port map( A1 => n21361, A2 => n14889, B1 => n21674, B2 => 
                           n21354, ZN => n6574);
   U14702 : OAI22_X1 port map( A1 => n21361, A2 => n14888, B1 => n21677, B2 => 
                           n21354, ZN => n6575);
   U14703 : OAI22_X1 port map( A1 => n21362, A2 => n14887, B1 => n21680, B2 => 
                           n21354, ZN => n6576);
   U14704 : OAI22_X1 port map( A1 => n21362, A2 => n14886, B1 => n21683, B2 => 
                           n21354, ZN => n6577);
   U14705 : OAI22_X1 port map( A1 => n21362, A2 => n14885, B1 => n21686, B2 => 
                           n21354, ZN => n6578);
   U14706 : OAI22_X1 port map( A1 => n21362, A2 => n14884, B1 => n21689, B2 => 
                           n21354, ZN => n6579);
   U14707 : OAI22_X1 port map( A1 => n21362, A2 => n14883, B1 => n21692, B2 => 
                           n21354, ZN => n6580);
   U14708 : OAI22_X1 port map( A1 => n21362, A2 => n14882, B1 => n21695, B2 => 
                           n21354, ZN => n6581);
   U14709 : OAI22_X1 port map( A1 => n21362, A2 => n14881, B1 => n21698, B2 => 
                           n21354, ZN => n6582);
   U14710 : OAI22_X1 port map( A1 => n21362, A2 => n14880, B1 => n21701, B2 => 
                           n21354, ZN => n6583);
   U14711 : OAI22_X1 port map( A1 => n21362, A2 => n14879, B1 => n21704, B2 => 
                           n21354, ZN => n6584);
   U14712 : OAI22_X1 port map( A1 => n21371, A2 => n14872, B1 => n21527, B2 => 
                           n21363, ZN => n6589);
   U14713 : OAI22_X1 port map( A1 => n21371, A2 => n14871, B1 => n21530, B2 => 
                           n21363, ZN => n6590);
   U14714 : OAI22_X1 port map( A1 => n21371, A2 => n14870, B1 => n21533, B2 => 
                           n21363, ZN => n6591);
   U14715 : OAI22_X1 port map( A1 => n21371, A2 => n14869, B1 => n21536, B2 => 
                           n21363, ZN => n6592);
   U14716 : OAI22_X1 port map( A1 => n21371, A2 => n14868, B1 => n21539, B2 => 
                           n21363, ZN => n6593);
   U14717 : OAI22_X1 port map( A1 => n21371, A2 => n14867, B1 => n21542, B2 => 
                           n21363, ZN => n6594);
   U14718 : OAI22_X1 port map( A1 => n21371, A2 => n14866, B1 => n21545, B2 => 
                           n21363, ZN => n6595);
   U14719 : OAI22_X1 port map( A1 => n21371, A2 => n14865, B1 => n21548, B2 => 
                           n21363, ZN => n6596);
   U14720 : OAI22_X1 port map( A1 => n21371, A2 => n14864, B1 => n21551, B2 => 
                           n21363, ZN => n6597);
   U14721 : OAI22_X1 port map( A1 => n21371, A2 => n14863, B1 => n21554, B2 => 
                           n21363, ZN => n6598);
   U14722 : OAI22_X1 port map( A1 => n21371, A2 => n14862, B1 => n21557, B2 => 
                           n21363, ZN => n6599);
   U14723 : OAI22_X1 port map( A1 => n21371, A2 => n14861, B1 => n21560, B2 => 
                           n21363, ZN => n6600);
   U14724 : OAI22_X1 port map( A1 => n21372, A2 => n14860, B1 => n21563, B2 => 
                           n21364, ZN => n6601);
   U14725 : OAI22_X1 port map( A1 => n21372, A2 => n14859, B1 => n21566, B2 => 
                           n21364, ZN => n6602);
   U14726 : OAI22_X1 port map( A1 => n21372, A2 => n14858, B1 => n21569, B2 => 
                           n21364, ZN => n6603);
   U14727 : OAI22_X1 port map( A1 => n21372, A2 => n14857, B1 => n21572, B2 => 
                           n21364, ZN => n6604);
   U14728 : OAI22_X1 port map( A1 => n21372, A2 => n14856, B1 => n21575, B2 => 
                           n21364, ZN => n6605);
   U14729 : OAI22_X1 port map( A1 => n21372, A2 => n14855, B1 => n21578, B2 => 
                           n21364, ZN => n6606);
   U14730 : OAI22_X1 port map( A1 => n21372, A2 => n14854, B1 => n21581, B2 => 
                           n21364, ZN => n6607);
   U14731 : OAI22_X1 port map( A1 => n21372, A2 => n14853, B1 => n21584, B2 => 
                           n21364, ZN => n6608);
   U14732 : OAI22_X1 port map( A1 => n21372, A2 => n14852, B1 => n21587, B2 => 
                           n21364, ZN => n6609);
   U14733 : OAI22_X1 port map( A1 => n21372, A2 => n14851, B1 => n21590, B2 => 
                           n21364, ZN => n6610);
   U14734 : OAI22_X1 port map( A1 => n21372, A2 => n14850, B1 => n21593, B2 => 
                           n21364, ZN => n6611);
   U14735 : OAI22_X1 port map( A1 => n21372, A2 => n14849, B1 => n21596, B2 => 
                           n21364, ZN => n6612);
   U14736 : OAI22_X1 port map( A1 => n21372, A2 => n14848, B1 => n21599, B2 => 
                           n21365, ZN => n6613);
   U14737 : OAI22_X1 port map( A1 => n21373, A2 => n14847, B1 => n21602, B2 => 
                           n21365, ZN => n6614);
   U14738 : OAI22_X1 port map( A1 => n21373, A2 => n14846, B1 => n21605, B2 => 
                           n21365, ZN => n6615);
   U14739 : OAI22_X1 port map( A1 => n21373, A2 => n14845, B1 => n21608, B2 => 
                           n21365, ZN => n6616);
   U14740 : OAI22_X1 port map( A1 => n21373, A2 => n14844, B1 => n21611, B2 => 
                           n21365, ZN => n6617);
   U14741 : OAI22_X1 port map( A1 => n21373, A2 => n14843, B1 => n21614, B2 => 
                           n21365, ZN => n6618);
   U14742 : OAI22_X1 port map( A1 => n21373, A2 => n14842, B1 => n21617, B2 => 
                           n21365, ZN => n6619);
   U14743 : OAI22_X1 port map( A1 => n21373, A2 => n14841, B1 => n21620, B2 => 
                           n21365, ZN => n6620);
   U14744 : OAI22_X1 port map( A1 => n21373, A2 => n14840, B1 => n21623, B2 => 
                           n21365, ZN => n6621);
   U14745 : OAI22_X1 port map( A1 => n21373, A2 => n14839, B1 => n21626, B2 => 
                           n21365, ZN => n6622);
   U14746 : OAI22_X1 port map( A1 => n21373, A2 => n14838, B1 => n21629, B2 => 
                           n21365, ZN => n6623);
   U14747 : OAI22_X1 port map( A1 => n21373, A2 => n14837, B1 => n21632, B2 => 
                           n21365, ZN => n6624);
   U14748 : OAI22_X1 port map( A1 => n21373, A2 => n14836, B1 => n21635, B2 => 
                           n21366, ZN => n6625);
   U14749 : OAI22_X1 port map( A1 => n21373, A2 => n14835, B1 => n21638, B2 => 
                           n21366, ZN => n6626);
   U14750 : OAI22_X1 port map( A1 => n21374, A2 => n14834, B1 => n21641, B2 => 
                           n21366, ZN => n6627);
   U14751 : OAI22_X1 port map( A1 => n21374, A2 => n14833, B1 => n21644, B2 => 
                           n21366, ZN => n6628);
   U14752 : OAI22_X1 port map( A1 => n21374, A2 => n14832, B1 => n21647, B2 => 
                           n21366, ZN => n6629);
   U14753 : OAI22_X1 port map( A1 => n21374, A2 => n14831, B1 => n21650, B2 => 
                           n21366, ZN => n6630);
   U14754 : OAI22_X1 port map( A1 => n21374, A2 => n14830, B1 => n21653, B2 => 
                           n21366, ZN => n6631);
   U14755 : OAI22_X1 port map( A1 => n21374, A2 => n14829, B1 => n21656, B2 => 
                           n21366, ZN => n6632);
   U14756 : OAI22_X1 port map( A1 => n21374, A2 => n14828, B1 => n21659, B2 => 
                           n21366, ZN => n6633);
   U14757 : OAI22_X1 port map( A1 => n21374, A2 => n14827, B1 => n21662, B2 => 
                           n21366, ZN => n6634);
   U14758 : OAI22_X1 port map( A1 => n21374, A2 => n14826, B1 => n21665, B2 => 
                           n21366, ZN => n6635);
   U14759 : OAI22_X1 port map( A1 => n21374, A2 => n14825, B1 => n21668, B2 => 
                           n21366, ZN => n6636);
   U14760 : OAI22_X1 port map( A1 => n21374, A2 => n14824, B1 => n21671, B2 => 
                           n21367, ZN => n6637);
   U14761 : OAI22_X1 port map( A1 => n21374, A2 => n14823, B1 => n21674, B2 => 
                           n21367, ZN => n6638);
   U14762 : OAI22_X1 port map( A1 => n21374, A2 => n14822, B1 => n21677, B2 => 
                           n21367, ZN => n6639);
   U14763 : OAI22_X1 port map( A1 => n21375, A2 => n14821, B1 => n21680, B2 => 
                           n21367, ZN => n6640);
   U14764 : OAI22_X1 port map( A1 => n21375, A2 => n14820, B1 => n21683, B2 => 
                           n21367, ZN => n6641);
   U14765 : OAI22_X1 port map( A1 => n21375, A2 => n14819, B1 => n21686, B2 => 
                           n21367, ZN => n6642);
   U14766 : OAI22_X1 port map( A1 => n21375, A2 => n14818, B1 => n21689, B2 => 
                           n21367, ZN => n6643);
   U14767 : OAI22_X1 port map( A1 => n21375, A2 => n14817, B1 => n21692, B2 => 
                           n21367, ZN => n6644);
   U14768 : OAI22_X1 port map( A1 => n21375, A2 => n14816, B1 => n21695, B2 => 
                           n21367, ZN => n6645);
   U14769 : OAI22_X1 port map( A1 => n21375, A2 => n14815, B1 => n21698, B2 => 
                           n21367, ZN => n6646);
   U14770 : OAI22_X1 port map( A1 => n21375, A2 => n14814, B1 => n21701, B2 => 
                           n21367, ZN => n6647);
   U14771 : OAI22_X1 port map( A1 => n21375, A2 => n14813, B1 => n21704, B2 => 
                           n21367, ZN => n6648);
   U14772 : OAI22_X1 port map( A1 => n21384, A2 => n14806, B1 => n21526, B2 => 
                           n21376, ZN => n6653);
   U14773 : OAI22_X1 port map( A1 => n21384, A2 => n14805, B1 => n21529, B2 => 
                           n21376, ZN => n6654);
   U14774 : OAI22_X1 port map( A1 => n21384, A2 => n14804, B1 => n21532, B2 => 
                           n21376, ZN => n6655);
   U14775 : OAI22_X1 port map( A1 => n21384, A2 => n14803, B1 => n21535, B2 => 
                           n21376, ZN => n6656);
   U14776 : OAI22_X1 port map( A1 => n21384, A2 => n14802, B1 => n21538, B2 => 
                           n21376, ZN => n6657);
   U14777 : OAI22_X1 port map( A1 => n21384, A2 => n14801, B1 => n21541, B2 => 
                           n21376, ZN => n6658);
   U14778 : OAI22_X1 port map( A1 => n21384, A2 => n14800, B1 => n21544, B2 => 
                           n21376, ZN => n6659);
   U14779 : OAI22_X1 port map( A1 => n21384, A2 => n14799, B1 => n21547, B2 => 
                           n21376, ZN => n6660);
   U14780 : OAI22_X1 port map( A1 => n21384, A2 => n14798, B1 => n21550, B2 => 
                           n21376, ZN => n6661);
   U14781 : OAI22_X1 port map( A1 => n21384, A2 => n14797, B1 => n21553, B2 => 
                           n21376, ZN => n6662);
   U14782 : OAI22_X1 port map( A1 => n21384, A2 => n14796, B1 => n21556, B2 => 
                           n21376, ZN => n6663);
   U14783 : OAI22_X1 port map( A1 => n21384, A2 => n14795, B1 => n21559, B2 => 
                           n21376, ZN => n6664);
   U14784 : OAI22_X1 port map( A1 => n21385, A2 => n14794, B1 => n21562, B2 => 
                           n21377, ZN => n6665);
   U14785 : OAI22_X1 port map( A1 => n21385, A2 => n14793, B1 => n21565, B2 => 
                           n21377, ZN => n6666);
   U14786 : OAI22_X1 port map( A1 => n21385, A2 => n14792, B1 => n21568, B2 => 
                           n21377, ZN => n6667);
   U14787 : OAI22_X1 port map( A1 => n21385, A2 => n14791, B1 => n21571, B2 => 
                           n21377, ZN => n6668);
   U14788 : OAI22_X1 port map( A1 => n21385, A2 => n14790, B1 => n21574, B2 => 
                           n21377, ZN => n6669);
   U14789 : OAI22_X1 port map( A1 => n21385, A2 => n14789, B1 => n21577, B2 => 
                           n21377, ZN => n6670);
   U14790 : OAI22_X1 port map( A1 => n21385, A2 => n14788, B1 => n21580, B2 => 
                           n21377, ZN => n6671);
   U14791 : OAI22_X1 port map( A1 => n21385, A2 => n14787, B1 => n21583, B2 => 
                           n21377, ZN => n6672);
   U14792 : OAI22_X1 port map( A1 => n21385, A2 => n14786, B1 => n21586, B2 => 
                           n21377, ZN => n6673);
   U14793 : OAI22_X1 port map( A1 => n21385, A2 => n14785, B1 => n21589, B2 => 
                           n21377, ZN => n6674);
   U14794 : OAI22_X1 port map( A1 => n21385, A2 => n14784, B1 => n21592, B2 => 
                           n21377, ZN => n6675);
   U14795 : OAI22_X1 port map( A1 => n21385, A2 => n14783, B1 => n21595, B2 => 
                           n21377, ZN => n6676);
   U14796 : OAI22_X1 port map( A1 => n21385, A2 => n14782, B1 => n21598, B2 => 
                           n21378, ZN => n6677);
   U14797 : OAI22_X1 port map( A1 => n21386, A2 => n14781, B1 => n21601, B2 => 
                           n21378, ZN => n6678);
   U14798 : OAI22_X1 port map( A1 => n21386, A2 => n14780, B1 => n21604, B2 => 
                           n21378, ZN => n6679);
   U14799 : OAI22_X1 port map( A1 => n21386, A2 => n14779, B1 => n21607, B2 => 
                           n21378, ZN => n6680);
   U14800 : OAI22_X1 port map( A1 => n21386, A2 => n14778, B1 => n21610, B2 => 
                           n21378, ZN => n6681);
   U14801 : OAI22_X1 port map( A1 => n21386, A2 => n14777, B1 => n21613, B2 => 
                           n21378, ZN => n6682);
   U14802 : OAI22_X1 port map( A1 => n21386, A2 => n14776, B1 => n21616, B2 => 
                           n21378, ZN => n6683);
   U14803 : OAI22_X1 port map( A1 => n21386, A2 => n14775, B1 => n21619, B2 => 
                           n21378, ZN => n6684);
   U14804 : OAI22_X1 port map( A1 => n21386, A2 => n14774, B1 => n21622, B2 => 
                           n21378, ZN => n6685);
   U14805 : OAI22_X1 port map( A1 => n21386, A2 => n14773, B1 => n21625, B2 => 
                           n21378, ZN => n6686);
   U14806 : OAI22_X1 port map( A1 => n21386, A2 => n14772, B1 => n21628, B2 => 
                           n21378, ZN => n6687);
   U14807 : OAI22_X1 port map( A1 => n21386, A2 => n14771, B1 => n21631, B2 => 
                           n21378, ZN => n6688);
   U14808 : OAI22_X1 port map( A1 => n21386, A2 => n14770, B1 => n21634, B2 => 
                           n21379, ZN => n6689);
   U14809 : OAI22_X1 port map( A1 => n21386, A2 => n14769, B1 => n21637, B2 => 
                           n21379, ZN => n6690);
   U14810 : OAI22_X1 port map( A1 => n21387, A2 => n14768, B1 => n21640, B2 => 
                           n21379, ZN => n6691);
   U14811 : OAI22_X1 port map( A1 => n21387, A2 => n14767, B1 => n21643, B2 => 
                           n21379, ZN => n6692);
   U14812 : OAI22_X1 port map( A1 => n21387, A2 => n14766, B1 => n21646, B2 => 
                           n21379, ZN => n6693);
   U14813 : OAI22_X1 port map( A1 => n21387, A2 => n14765, B1 => n21649, B2 => 
                           n21379, ZN => n6694);
   U14814 : OAI22_X1 port map( A1 => n21387, A2 => n14764, B1 => n21652, B2 => 
                           n21379, ZN => n6695);
   U14815 : OAI22_X1 port map( A1 => n21387, A2 => n14763, B1 => n21655, B2 => 
                           n21379, ZN => n6696);
   U14816 : OAI22_X1 port map( A1 => n21387, A2 => n14762, B1 => n21658, B2 => 
                           n21379, ZN => n6697);
   U14817 : OAI22_X1 port map( A1 => n21387, A2 => n14761, B1 => n21661, B2 => 
                           n21379, ZN => n6698);
   U14818 : OAI22_X1 port map( A1 => n21387, A2 => n14760, B1 => n21664, B2 => 
                           n21379, ZN => n6699);
   U14819 : OAI22_X1 port map( A1 => n21387, A2 => n14759, B1 => n21667, B2 => 
                           n21379, ZN => n6700);
   U14820 : OAI22_X1 port map( A1 => n21387, A2 => n14758, B1 => n21670, B2 => 
                           n21380, ZN => n6701);
   U14821 : OAI22_X1 port map( A1 => n21387, A2 => n14757, B1 => n21673, B2 => 
                           n21380, ZN => n6702);
   U14822 : OAI22_X1 port map( A1 => n21387, A2 => n14756, B1 => n21676, B2 => 
                           n21380, ZN => n6703);
   U14823 : OAI22_X1 port map( A1 => n21388, A2 => n14755, B1 => n21679, B2 => 
                           n21380, ZN => n6704);
   U14824 : OAI22_X1 port map( A1 => n21388, A2 => n14754, B1 => n21682, B2 => 
                           n21380, ZN => n6705);
   U14825 : OAI22_X1 port map( A1 => n21388, A2 => n14753, B1 => n21685, B2 => 
                           n21380, ZN => n6706);
   U14826 : OAI22_X1 port map( A1 => n21388, A2 => n14752, B1 => n21688, B2 => 
                           n21380, ZN => n6707);
   U14827 : OAI22_X1 port map( A1 => n21388, A2 => n14751, B1 => n21691, B2 => 
                           n21380, ZN => n6708);
   U14828 : OAI22_X1 port map( A1 => n21388, A2 => n14750, B1 => n21694, B2 => 
                           n21380, ZN => n6709);
   U14829 : OAI22_X1 port map( A1 => n21388, A2 => n14749, B1 => n21697, B2 => 
                           n21380, ZN => n6710);
   U14830 : OAI22_X1 port map( A1 => n21388, A2 => n14748, B1 => n21700, B2 => 
                           n21380, ZN => n6711);
   U14831 : OAI22_X1 port map( A1 => n21388, A2 => n14747, B1 => n21703, B2 => 
                           n21380, ZN => n6712);
   U14832 : OAI22_X1 port map( A1 => n21423, A2 => n14606, B1 => n21526, B2 => 
                           n21415, ZN => n6845);
   U14833 : OAI22_X1 port map( A1 => n21423, A2 => n14605, B1 => n21529, B2 => 
                           n21415, ZN => n6846);
   U14834 : OAI22_X1 port map( A1 => n21423, A2 => n14604, B1 => n21532, B2 => 
                           n21415, ZN => n6847);
   U14835 : OAI22_X1 port map( A1 => n21423, A2 => n14603, B1 => n21535, B2 => 
                           n21415, ZN => n6848);
   U14836 : OAI22_X1 port map( A1 => n21423, A2 => n14602, B1 => n21538, B2 => 
                           n21415, ZN => n6849);
   U14837 : OAI22_X1 port map( A1 => n21423, A2 => n14601, B1 => n21541, B2 => 
                           n21415, ZN => n6850);
   U14838 : OAI22_X1 port map( A1 => n21423, A2 => n14600, B1 => n21544, B2 => 
                           n21415, ZN => n6851);
   U14839 : OAI22_X1 port map( A1 => n21423, A2 => n14599, B1 => n21547, B2 => 
                           n21415, ZN => n6852);
   U14840 : OAI22_X1 port map( A1 => n21423, A2 => n14598, B1 => n21550, B2 => 
                           n21415, ZN => n6853);
   U14841 : OAI22_X1 port map( A1 => n21423, A2 => n14597, B1 => n21553, B2 => 
                           n21415, ZN => n6854);
   U14842 : OAI22_X1 port map( A1 => n21423, A2 => n14596, B1 => n21556, B2 => 
                           n21415, ZN => n6855);
   U14843 : OAI22_X1 port map( A1 => n21423, A2 => n14595, B1 => n21559, B2 => 
                           n21415, ZN => n6856);
   U14844 : OAI22_X1 port map( A1 => n21424, A2 => n14594, B1 => n21562, B2 => 
                           n21416, ZN => n6857);
   U14845 : OAI22_X1 port map( A1 => n21424, A2 => n14593, B1 => n21565, B2 => 
                           n21416, ZN => n6858);
   U14846 : OAI22_X1 port map( A1 => n21424, A2 => n14592, B1 => n21568, B2 => 
                           n21416, ZN => n6859);
   U14847 : OAI22_X1 port map( A1 => n21424, A2 => n14591, B1 => n21571, B2 => 
                           n21416, ZN => n6860);
   U14848 : OAI22_X1 port map( A1 => n21424, A2 => n14590, B1 => n21574, B2 => 
                           n21416, ZN => n6861);
   U14849 : OAI22_X1 port map( A1 => n21424, A2 => n14589, B1 => n21577, B2 => 
                           n21416, ZN => n6862);
   U14850 : OAI22_X1 port map( A1 => n21424, A2 => n14588, B1 => n21580, B2 => 
                           n21416, ZN => n6863);
   U14851 : OAI22_X1 port map( A1 => n21424, A2 => n14587, B1 => n21583, B2 => 
                           n21416, ZN => n6864);
   U14852 : OAI22_X1 port map( A1 => n21424, A2 => n14586, B1 => n21586, B2 => 
                           n21416, ZN => n6865);
   U14853 : OAI22_X1 port map( A1 => n21424, A2 => n14585, B1 => n21589, B2 => 
                           n21416, ZN => n6866);
   U14854 : OAI22_X1 port map( A1 => n21424, A2 => n14584, B1 => n21592, B2 => 
                           n21416, ZN => n6867);
   U14855 : OAI22_X1 port map( A1 => n21424, A2 => n14583, B1 => n21595, B2 => 
                           n21416, ZN => n6868);
   U14856 : OAI22_X1 port map( A1 => n21424, A2 => n14582, B1 => n21598, B2 => 
                           n21417, ZN => n6869);
   U14857 : OAI22_X1 port map( A1 => n21425, A2 => n14581, B1 => n21601, B2 => 
                           n21417, ZN => n6870);
   U14858 : OAI22_X1 port map( A1 => n21425, A2 => n14580, B1 => n21604, B2 => 
                           n21417, ZN => n6871);
   U14859 : OAI22_X1 port map( A1 => n21425, A2 => n14579, B1 => n21607, B2 => 
                           n21417, ZN => n6872);
   U14860 : OAI22_X1 port map( A1 => n21425, A2 => n14578, B1 => n21610, B2 => 
                           n21417, ZN => n6873);
   U14861 : OAI22_X1 port map( A1 => n21425, A2 => n14577, B1 => n21613, B2 => 
                           n21417, ZN => n6874);
   U14862 : OAI22_X1 port map( A1 => n21425, A2 => n14576, B1 => n21616, B2 => 
                           n21417, ZN => n6875);
   U14863 : OAI22_X1 port map( A1 => n21425, A2 => n14575, B1 => n21619, B2 => 
                           n21417, ZN => n6876);
   U14864 : OAI22_X1 port map( A1 => n21425, A2 => n14574, B1 => n21622, B2 => 
                           n21417, ZN => n6877);
   U14865 : OAI22_X1 port map( A1 => n21425, A2 => n14573, B1 => n21625, B2 => 
                           n21417, ZN => n6878);
   U14866 : OAI22_X1 port map( A1 => n21425, A2 => n14572, B1 => n21628, B2 => 
                           n21417, ZN => n6879);
   U14867 : OAI22_X1 port map( A1 => n21425, A2 => n14571, B1 => n21631, B2 => 
                           n21417, ZN => n6880);
   U14868 : OAI22_X1 port map( A1 => n21425, A2 => n14570, B1 => n21634, B2 => 
                           n21418, ZN => n6881);
   U14869 : OAI22_X1 port map( A1 => n21425, A2 => n14569, B1 => n21637, B2 => 
                           n21418, ZN => n6882);
   U14870 : OAI22_X1 port map( A1 => n21426, A2 => n14568, B1 => n21640, B2 => 
                           n21418, ZN => n6883);
   U14871 : OAI22_X1 port map( A1 => n21426, A2 => n14567, B1 => n21643, B2 => 
                           n21418, ZN => n6884);
   U14872 : OAI22_X1 port map( A1 => n21426, A2 => n14566, B1 => n21646, B2 => 
                           n21418, ZN => n6885);
   U14873 : OAI22_X1 port map( A1 => n21426, A2 => n14565, B1 => n21649, B2 => 
                           n21418, ZN => n6886);
   U14874 : OAI22_X1 port map( A1 => n21426, A2 => n14564, B1 => n21652, B2 => 
                           n21418, ZN => n6887);
   U14875 : OAI22_X1 port map( A1 => n21426, A2 => n14563, B1 => n21655, B2 => 
                           n21418, ZN => n6888);
   U14876 : OAI22_X1 port map( A1 => n21426, A2 => n14562, B1 => n21658, B2 => 
                           n21418, ZN => n6889);
   U14877 : OAI22_X1 port map( A1 => n21426, A2 => n14561, B1 => n21661, B2 => 
                           n21418, ZN => n6890);
   U14878 : OAI22_X1 port map( A1 => n21426, A2 => n14560, B1 => n21664, B2 => 
                           n21418, ZN => n6891);
   U14879 : OAI22_X1 port map( A1 => n21426, A2 => n14559, B1 => n21667, B2 => 
                           n21418, ZN => n6892);
   U14880 : OAI22_X1 port map( A1 => n21426, A2 => n14558, B1 => n21670, B2 => 
                           n21419, ZN => n6893);
   U14881 : OAI22_X1 port map( A1 => n21426, A2 => n14557, B1 => n21673, B2 => 
                           n21419, ZN => n6894);
   U14882 : OAI22_X1 port map( A1 => n21426, A2 => n14556, B1 => n21676, B2 => 
                           n21419, ZN => n6895);
   U14883 : OAI22_X1 port map( A1 => n21427, A2 => n14555, B1 => n21679, B2 => 
                           n21419, ZN => n6896);
   U14884 : OAI22_X1 port map( A1 => n21427, A2 => n14554, B1 => n21682, B2 => 
                           n21419, ZN => n6897);
   U14885 : OAI22_X1 port map( A1 => n21427, A2 => n14553, B1 => n21685, B2 => 
                           n21419, ZN => n6898);
   U14886 : OAI22_X1 port map( A1 => n21427, A2 => n14552, B1 => n21688, B2 => 
                           n21419, ZN => n6899);
   U14887 : OAI22_X1 port map( A1 => n21427, A2 => n14551, B1 => n21691, B2 => 
                           n21419, ZN => n6900);
   U14888 : OAI22_X1 port map( A1 => n21427, A2 => n14550, B1 => n21694, B2 => 
                           n21419, ZN => n6901);
   U14889 : OAI22_X1 port map( A1 => n21427, A2 => n14549, B1 => n21697, B2 => 
                           n21419, ZN => n6902);
   U14890 : OAI22_X1 port map( A1 => n21427, A2 => n14548, B1 => n21700, B2 => 
                           n21419, ZN => n6903);
   U14891 : OAI22_X1 port map( A1 => n21427, A2 => n14547, B1 => n21703, B2 => 
                           n21419, ZN => n6904);
   U14892 : OAI22_X1 port map( A1 => n21436, A2 => n14540, B1 => n21526, B2 => 
                           n21428, ZN => n6909);
   U14893 : OAI22_X1 port map( A1 => n21436, A2 => n14539, B1 => n21529, B2 => 
                           n21428, ZN => n6910);
   U14894 : OAI22_X1 port map( A1 => n21436, A2 => n14538, B1 => n21532, B2 => 
                           n21428, ZN => n6911);
   U14895 : OAI22_X1 port map( A1 => n21436, A2 => n14537, B1 => n21535, B2 => 
                           n21428, ZN => n6912);
   U14896 : OAI22_X1 port map( A1 => n21436, A2 => n14536, B1 => n21538, B2 => 
                           n21428, ZN => n6913);
   U14897 : OAI22_X1 port map( A1 => n21436, A2 => n14535, B1 => n21541, B2 => 
                           n21428, ZN => n6914);
   U14898 : OAI22_X1 port map( A1 => n21436, A2 => n14534, B1 => n21544, B2 => 
                           n21428, ZN => n6915);
   U14899 : OAI22_X1 port map( A1 => n21436, A2 => n14533, B1 => n21547, B2 => 
                           n21428, ZN => n6916);
   U14900 : OAI22_X1 port map( A1 => n21436, A2 => n14532, B1 => n21550, B2 => 
                           n21428, ZN => n6917);
   U14901 : OAI22_X1 port map( A1 => n21436, A2 => n14531, B1 => n21553, B2 => 
                           n21428, ZN => n6918);
   U14902 : OAI22_X1 port map( A1 => n21436, A2 => n14530, B1 => n21556, B2 => 
                           n21428, ZN => n6919);
   U14903 : OAI22_X1 port map( A1 => n21436, A2 => n14529, B1 => n21559, B2 => 
                           n21428, ZN => n6920);
   U14904 : OAI22_X1 port map( A1 => n21437, A2 => n14528, B1 => n21562, B2 => 
                           n21429, ZN => n6921);
   U14905 : OAI22_X1 port map( A1 => n21437, A2 => n14527, B1 => n21565, B2 => 
                           n21429, ZN => n6922);
   U14906 : OAI22_X1 port map( A1 => n21437, A2 => n14526, B1 => n21568, B2 => 
                           n21429, ZN => n6923);
   U14907 : OAI22_X1 port map( A1 => n21437, A2 => n14525, B1 => n21571, B2 => 
                           n21429, ZN => n6924);
   U14908 : OAI22_X1 port map( A1 => n21437, A2 => n14524, B1 => n21574, B2 => 
                           n21429, ZN => n6925);
   U14909 : OAI22_X1 port map( A1 => n21437, A2 => n14523, B1 => n21577, B2 => 
                           n21429, ZN => n6926);
   U14910 : OAI22_X1 port map( A1 => n21437, A2 => n14522, B1 => n21580, B2 => 
                           n21429, ZN => n6927);
   U14911 : OAI22_X1 port map( A1 => n21437, A2 => n14521, B1 => n21583, B2 => 
                           n21429, ZN => n6928);
   U14912 : OAI22_X1 port map( A1 => n21437, A2 => n14520, B1 => n21586, B2 => 
                           n21429, ZN => n6929);
   U14913 : OAI22_X1 port map( A1 => n21437, A2 => n14519, B1 => n21589, B2 => 
                           n21429, ZN => n6930);
   U14914 : OAI22_X1 port map( A1 => n21437, A2 => n14518, B1 => n21592, B2 => 
                           n21429, ZN => n6931);
   U14915 : OAI22_X1 port map( A1 => n21437, A2 => n14517, B1 => n21595, B2 => 
                           n21429, ZN => n6932);
   U14916 : OAI22_X1 port map( A1 => n21437, A2 => n14516, B1 => n21598, B2 => 
                           n21430, ZN => n6933);
   U14917 : OAI22_X1 port map( A1 => n21438, A2 => n14515, B1 => n21601, B2 => 
                           n21430, ZN => n6934);
   U14918 : OAI22_X1 port map( A1 => n21438, A2 => n14514, B1 => n21604, B2 => 
                           n21430, ZN => n6935);
   U14919 : OAI22_X1 port map( A1 => n21438, A2 => n14513, B1 => n21607, B2 => 
                           n21430, ZN => n6936);
   U14920 : OAI22_X1 port map( A1 => n21438, A2 => n14512, B1 => n21610, B2 => 
                           n21430, ZN => n6937);
   U14921 : OAI22_X1 port map( A1 => n21438, A2 => n14511, B1 => n21613, B2 => 
                           n21430, ZN => n6938);
   U14922 : OAI22_X1 port map( A1 => n21438, A2 => n14510, B1 => n21616, B2 => 
                           n21430, ZN => n6939);
   U14923 : OAI22_X1 port map( A1 => n21438, A2 => n14509, B1 => n21619, B2 => 
                           n21430, ZN => n6940);
   U14924 : OAI22_X1 port map( A1 => n21438, A2 => n14508, B1 => n21622, B2 => 
                           n21430, ZN => n6941);
   U14925 : OAI22_X1 port map( A1 => n21438, A2 => n14507, B1 => n21625, B2 => 
                           n21430, ZN => n6942);
   U14926 : OAI22_X1 port map( A1 => n21438, A2 => n14506, B1 => n21628, B2 => 
                           n21430, ZN => n6943);
   U14927 : OAI22_X1 port map( A1 => n21438, A2 => n14505, B1 => n21631, B2 => 
                           n21430, ZN => n6944);
   U14928 : OAI22_X1 port map( A1 => n21438, A2 => n14504, B1 => n21634, B2 => 
                           n21431, ZN => n6945);
   U14929 : OAI22_X1 port map( A1 => n21438, A2 => n14503, B1 => n21637, B2 => 
                           n21431, ZN => n6946);
   U14930 : OAI22_X1 port map( A1 => n21439, A2 => n14502, B1 => n21640, B2 => 
                           n21431, ZN => n6947);
   U14931 : OAI22_X1 port map( A1 => n21439, A2 => n14501, B1 => n21643, B2 => 
                           n21431, ZN => n6948);
   U14932 : OAI22_X1 port map( A1 => n21439, A2 => n14500, B1 => n21646, B2 => 
                           n21431, ZN => n6949);
   U14933 : OAI22_X1 port map( A1 => n21439, A2 => n14499, B1 => n21649, B2 => 
                           n21431, ZN => n6950);
   U14934 : OAI22_X1 port map( A1 => n21439, A2 => n14498, B1 => n21652, B2 => 
                           n21431, ZN => n6951);
   U14935 : OAI22_X1 port map( A1 => n21439, A2 => n14497, B1 => n21655, B2 => 
                           n21431, ZN => n6952);
   U14936 : OAI22_X1 port map( A1 => n21439, A2 => n14496, B1 => n21658, B2 => 
                           n21431, ZN => n6953);
   U14937 : OAI22_X1 port map( A1 => n21439, A2 => n14495, B1 => n21661, B2 => 
                           n21431, ZN => n6954);
   U14938 : OAI22_X1 port map( A1 => n21439, A2 => n14494, B1 => n21664, B2 => 
                           n21431, ZN => n6955);
   U14939 : OAI22_X1 port map( A1 => n21439, A2 => n14493, B1 => n21667, B2 => 
                           n21431, ZN => n6956);
   U14940 : OAI22_X1 port map( A1 => n21439, A2 => n14492, B1 => n21670, B2 => 
                           n21432, ZN => n6957);
   U14941 : OAI22_X1 port map( A1 => n21439, A2 => n14491, B1 => n21673, B2 => 
                           n21432, ZN => n6958);
   U14942 : OAI22_X1 port map( A1 => n21439, A2 => n14490, B1 => n21676, B2 => 
                           n21432, ZN => n6959);
   U14943 : OAI22_X1 port map( A1 => n21440, A2 => n14489, B1 => n21679, B2 => 
                           n21432, ZN => n6960);
   U14944 : OAI22_X1 port map( A1 => n21440, A2 => n14488, B1 => n21682, B2 => 
                           n21432, ZN => n6961);
   U14945 : OAI22_X1 port map( A1 => n21440, A2 => n14487, B1 => n21685, B2 => 
                           n21432, ZN => n6962);
   U14946 : OAI22_X1 port map( A1 => n21440, A2 => n14486, B1 => n21688, B2 => 
                           n21432, ZN => n6963);
   U14947 : OAI22_X1 port map( A1 => n21440, A2 => n14485, B1 => n21691, B2 => 
                           n21432, ZN => n6964);
   U14948 : OAI22_X1 port map( A1 => n21440, A2 => n14484, B1 => n21694, B2 => 
                           n21432, ZN => n6965);
   U14949 : OAI22_X1 port map( A1 => n21440, A2 => n14483, B1 => n21697, B2 => 
                           n21432, ZN => n6966);
   U14950 : OAI22_X1 port map( A1 => n21440, A2 => n14482, B1 => n21700, B2 => 
                           n21432, ZN => n6967);
   U14951 : OAI22_X1 port map( A1 => n21440, A2 => n14481, B1 => n21703, B2 => 
                           n21432, ZN => n6968);
   U14952 : OAI22_X1 port map( A1 => n21462, A2 => n14404, B1 => n21526, B2 => 
                           n21454, ZN => n7037);
   U14953 : OAI22_X1 port map( A1 => n21462, A2 => n14403, B1 => n21529, B2 => 
                           n21454, ZN => n7038);
   U14954 : OAI22_X1 port map( A1 => n21462, A2 => n14402, B1 => n21532, B2 => 
                           n21454, ZN => n7039);
   U14955 : OAI22_X1 port map( A1 => n21462, A2 => n14401, B1 => n21535, B2 => 
                           n21454, ZN => n7040);
   U14956 : OAI22_X1 port map( A1 => n21462, A2 => n14400, B1 => n21538, B2 => 
                           n21454, ZN => n7041);
   U14957 : OAI22_X1 port map( A1 => n21462, A2 => n14399, B1 => n21541, B2 => 
                           n21454, ZN => n7042);
   U14958 : OAI22_X1 port map( A1 => n21462, A2 => n14398, B1 => n21544, B2 => 
                           n21454, ZN => n7043);
   U14959 : OAI22_X1 port map( A1 => n21462, A2 => n14397, B1 => n21547, B2 => 
                           n21454, ZN => n7044);
   U14960 : OAI22_X1 port map( A1 => n21462, A2 => n14396, B1 => n21550, B2 => 
                           n21454, ZN => n7045);
   U14961 : OAI22_X1 port map( A1 => n21462, A2 => n14395, B1 => n21553, B2 => 
                           n21454, ZN => n7046);
   U14962 : OAI22_X1 port map( A1 => n21462, A2 => n14394, B1 => n21556, B2 => 
                           n21454, ZN => n7047);
   U14963 : OAI22_X1 port map( A1 => n21462, A2 => n14393, B1 => n21559, B2 => 
                           n21454, ZN => n7048);
   U14964 : OAI22_X1 port map( A1 => n21463, A2 => n14392, B1 => n21562, B2 => 
                           n21455, ZN => n7049);
   U14965 : OAI22_X1 port map( A1 => n21463, A2 => n14391, B1 => n21565, B2 => 
                           n21455, ZN => n7050);
   U14966 : OAI22_X1 port map( A1 => n21463, A2 => n14390, B1 => n21568, B2 => 
                           n21455, ZN => n7051);
   U14967 : OAI22_X1 port map( A1 => n21463, A2 => n14389, B1 => n21571, B2 => 
                           n21455, ZN => n7052);
   U14968 : OAI22_X1 port map( A1 => n21463, A2 => n14388, B1 => n21574, B2 => 
                           n21455, ZN => n7053);
   U14969 : OAI22_X1 port map( A1 => n21463, A2 => n14387, B1 => n21577, B2 => 
                           n21455, ZN => n7054);
   U14970 : OAI22_X1 port map( A1 => n21463, A2 => n14386, B1 => n21580, B2 => 
                           n21455, ZN => n7055);
   U14971 : OAI22_X1 port map( A1 => n21463, A2 => n14385, B1 => n21583, B2 => 
                           n21455, ZN => n7056);
   U14972 : OAI22_X1 port map( A1 => n21463, A2 => n14384, B1 => n21586, B2 => 
                           n21455, ZN => n7057);
   U14973 : OAI22_X1 port map( A1 => n21463, A2 => n14383, B1 => n21589, B2 => 
                           n21455, ZN => n7058);
   U14974 : OAI22_X1 port map( A1 => n21463, A2 => n14382, B1 => n21592, B2 => 
                           n21455, ZN => n7059);
   U14975 : OAI22_X1 port map( A1 => n21463, A2 => n14381, B1 => n21595, B2 => 
                           n21455, ZN => n7060);
   U14976 : OAI22_X1 port map( A1 => n21463, A2 => n14380, B1 => n21598, B2 => 
                           n21456, ZN => n7061);
   U14977 : OAI22_X1 port map( A1 => n21464, A2 => n14379, B1 => n21601, B2 => 
                           n21456, ZN => n7062);
   U14978 : OAI22_X1 port map( A1 => n21464, A2 => n14378, B1 => n21604, B2 => 
                           n21456, ZN => n7063);
   U14979 : OAI22_X1 port map( A1 => n21464, A2 => n14377, B1 => n21607, B2 => 
                           n21456, ZN => n7064);
   U14980 : OAI22_X1 port map( A1 => n21464, A2 => n14376, B1 => n21610, B2 => 
                           n21456, ZN => n7065);
   U14981 : OAI22_X1 port map( A1 => n21464, A2 => n14375, B1 => n21613, B2 => 
                           n21456, ZN => n7066);
   U14982 : OAI22_X1 port map( A1 => n21464, A2 => n14374, B1 => n21616, B2 => 
                           n21456, ZN => n7067);
   U14983 : OAI22_X1 port map( A1 => n21464, A2 => n14373, B1 => n21619, B2 => 
                           n21456, ZN => n7068);
   U14984 : OAI22_X1 port map( A1 => n21464, A2 => n14372, B1 => n21622, B2 => 
                           n21456, ZN => n7069);
   U14985 : OAI22_X1 port map( A1 => n21464, A2 => n14371, B1 => n21625, B2 => 
                           n21456, ZN => n7070);
   U14986 : OAI22_X1 port map( A1 => n21464, A2 => n14370, B1 => n21628, B2 => 
                           n21456, ZN => n7071);
   U14987 : OAI22_X1 port map( A1 => n21464, A2 => n14369, B1 => n21631, B2 => 
                           n21456, ZN => n7072);
   U14988 : OAI22_X1 port map( A1 => n21464, A2 => n14368, B1 => n21634, B2 => 
                           n21457, ZN => n7073);
   U14989 : OAI22_X1 port map( A1 => n21464, A2 => n14367, B1 => n21637, B2 => 
                           n21457, ZN => n7074);
   U14990 : OAI22_X1 port map( A1 => n21465, A2 => n14366, B1 => n21640, B2 => 
                           n21457, ZN => n7075);
   U14991 : OAI22_X1 port map( A1 => n21465, A2 => n14365, B1 => n21643, B2 => 
                           n21457, ZN => n7076);
   U14992 : OAI22_X1 port map( A1 => n21465, A2 => n14364, B1 => n21646, B2 => 
                           n21457, ZN => n7077);
   U14993 : OAI22_X1 port map( A1 => n21465, A2 => n14363, B1 => n21649, B2 => 
                           n21457, ZN => n7078);
   U14994 : OAI22_X1 port map( A1 => n21465, A2 => n14362, B1 => n21652, B2 => 
                           n21457, ZN => n7079);
   U14995 : OAI22_X1 port map( A1 => n21465, A2 => n14361, B1 => n21655, B2 => 
                           n21457, ZN => n7080);
   U14996 : OAI22_X1 port map( A1 => n21465, A2 => n14360, B1 => n21658, B2 => 
                           n21457, ZN => n7081);
   U14997 : OAI22_X1 port map( A1 => n21465, A2 => n14359, B1 => n21661, B2 => 
                           n21457, ZN => n7082);
   U14998 : OAI22_X1 port map( A1 => n21465, A2 => n14358, B1 => n21664, B2 => 
                           n21457, ZN => n7083);
   U14999 : OAI22_X1 port map( A1 => n21465, A2 => n14357, B1 => n21667, B2 => 
                           n21457, ZN => n7084);
   U15000 : OAI22_X1 port map( A1 => n21465, A2 => n14356, B1 => n21670, B2 => 
                           n21458, ZN => n7085);
   U15001 : OAI22_X1 port map( A1 => n21465, A2 => n14355, B1 => n21673, B2 => 
                           n21458, ZN => n7086);
   U15002 : OAI22_X1 port map( A1 => n21465, A2 => n14354, B1 => n21676, B2 => 
                           n21458, ZN => n7087);
   U15003 : OAI22_X1 port map( A1 => n21466, A2 => n14353, B1 => n21679, B2 => 
                           n21458, ZN => n7088);
   U15004 : OAI22_X1 port map( A1 => n21466, A2 => n14352, B1 => n21682, B2 => 
                           n21458, ZN => n7089);
   U15005 : OAI22_X1 port map( A1 => n21466, A2 => n14351, B1 => n21685, B2 => 
                           n21458, ZN => n7090);
   U15006 : OAI22_X1 port map( A1 => n21466, A2 => n14350, B1 => n21688, B2 => 
                           n21458, ZN => n7091);
   U15007 : OAI22_X1 port map( A1 => n21466, A2 => n14349, B1 => n21691, B2 => 
                           n21458, ZN => n7092);
   U15008 : OAI22_X1 port map( A1 => n21466, A2 => n14348, B1 => n21694, B2 => 
                           n21458, ZN => n7093);
   U15009 : OAI22_X1 port map( A1 => n21466, A2 => n14347, B1 => n21697, B2 => 
                           n21458, ZN => n7094);
   U15010 : OAI22_X1 port map( A1 => n21466, A2 => n14346, B1 => n21700, B2 => 
                           n21458, ZN => n7095);
   U15011 : OAI22_X1 port map( A1 => n21466, A2 => n14345, B1 => n21703, B2 => 
                           n21458, ZN => n7096);
   U15012 : OAI22_X1 port map( A1 => n21475, A2 => n14337, B1 => n21526, B2 => 
                           n21467, ZN => n7101);
   U15013 : OAI22_X1 port map( A1 => n21475, A2 => n14336, B1 => n21529, B2 => 
                           n21467, ZN => n7102);
   U15014 : OAI22_X1 port map( A1 => n21475, A2 => n14335, B1 => n21532, B2 => 
                           n21467, ZN => n7103);
   U15015 : OAI22_X1 port map( A1 => n21475, A2 => n14334, B1 => n21535, B2 => 
                           n21467, ZN => n7104);
   U15016 : OAI22_X1 port map( A1 => n21475, A2 => n14333, B1 => n21538, B2 => 
                           n21467, ZN => n7105);
   U15017 : OAI22_X1 port map( A1 => n21475, A2 => n14332, B1 => n21541, B2 => 
                           n21467, ZN => n7106);
   U15018 : OAI22_X1 port map( A1 => n21475, A2 => n14331, B1 => n21544, B2 => 
                           n21467, ZN => n7107);
   U15019 : OAI22_X1 port map( A1 => n21475, A2 => n14330, B1 => n21547, B2 => 
                           n21467, ZN => n7108);
   U15020 : OAI22_X1 port map( A1 => n21475, A2 => n14329, B1 => n21550, B2 => 
                           n21467, ZN => n7109);
   U15021 : OAI22_X1 port map( A1 => n21475, A2 => n14328, B1 => n21553, B2 => 
                           n21467, ZN => n7110);
   U15022 : OAI22_X1 port map( A1 => n21475, A2 => n14327, B1 => n21556, B2 => 
                           n21467, ZN => n7111);
   U15023 : OAI22_X1 port map( A1 => n21475, A2 => n14326, B1 => n21559, B2 => 
                           n21467, ZN => n7112);
   U15024 : OAI22_X1 port map( A1 => n21476, A2 => n14325, B1 => n21562, B2 => 
                           n21468, ZN => n7113);
   U15025 : OAI22_X1 port map( A1 => n21476, A2 => n14324, B1 => n21565, B2 => 
                           n21468, ZN => n7114);
   U15026 : OAI22_X1 port map( A1 => n21476, A2 => n14323, B1 => n21568, B2 => 
                           n21468, ZN => n7115);
   U15027 : OAI22_X1 port map( A1 => n21476, A2 => n14322, B1 => n21571, B2 => 
                           n21468, ZN => n7116);
   U15028 : OAI22_X1 port map( A1 => n21476, A2 => n14321, B1 => n21574, B2 => 
                           n21468, ZN => n7117);
   U15029 : OAI22_X1 port map( A1 => n21476, A2 => n14320, B1 => n21577, B2 => 
                           n21468, ZN => n7118);
   U15030 : OAI22_X1 port map( A1 => n21476, A2 => n14319, B1 => n21580, B2 => 
                           n21468, ZN => n7119);
   U15031 : OAI22_X1 port map( A1 => n21476, A2 => n14318, B1 => n21583, B2 => 
                           n21468, ZN => n7120);
   U15032 : OAI22_X1 port map( A1 => n21476, A2 => n14317, B1 => n21586, B2 => 
                           n21468, ZN => n7121);
   U15033 : OAI22_X1 port map( A1 => n21476, A2 => n14316, B1 => n21589, B2 => 
                           n21468, ZN => n7122);
   U15034 : OAI22_X1 port map( A1 => n21476, A2 => n14315, B1 => n21592, B2 => 
                           n21468, ZN => n7123);
   U15035 : OAI22_X1 port map( A1 => n21476, A2 => n14314, B1 => n21595, B2 => 
                           n21468, ZN => n7124);
   U15036 : OAI22_X1 port map( A1 => n21476, A2 => n14313, B1 => n21598, B2 => 
                           n21469, ZN => n7125);
   U15037 : OAI22_X1 port map( A1 => n21477, A2 => n14312, B1 => n21601, B2 => 
                           n21469, ZN => n7126);
   U15038 : OAI22_X1 port map( A1 => n21477, A2 => n14311, B1 => n21604, B2 => 
                           n21469, ZN => n7127);
   U15039 : OAI22_X1 port map( A1 => n21477, A2 => n14310, B1 => n21607, B2 => 
                           n21469, ZN => n7128);
   U15040 : OAI22_X1 port map( A1 => n21477, A2 => n14309, B1 => n21610, B2 => 
                           n21469, ZN => n7129);
   U15041 : OAI22_X1 port map( A1 => n21477, A2 => n14308, B1 => n21613, B2 => 
                           n21469, ZN => n7130);
   U15042 : OAI22_X1 port map( A1 => n21477, A2 => n14307, B1 => n21616, B2 => 
                           n21469, ZN => n7131);
   U15043 : OAI22_X1 port map( A1 => n21477, A2 => n14306, B1 => n21619, B2 => 
                           n21469, ZN => n7132);
   U15044 : OAI22_X1 port map( A1 => n21477, A2 => n14305, B1 => n21622, B2 => 
                           n21469, ZN => n7133);
   U15045 : OAI22_X1 port map( A1 => n21477, A2 => n14304, B1 => n21625, B2 => 
                           n21469, ZN => n7134);
   U15046 : OAI22_X1 port map( A1 => n21477, A2 => n14303, B1 => n21628, B2 => 
                           n21469, ZN => n7135);
   U15047 : OAI22_X1 port map( A1 => n21477, A2 => n14302, B1 => n21631, B2 => 
                           n21469, ZN => n7136);
   U15048 : OAI22_X1 port map( A1 => n21477, A2 => n14301, B1 => n21634, B2 => 
                           n21470, ZN => n7137);
   U15049 : OAI22_X1 port map( A1 => n21477, A2 => n14300, B1 => n21637, B2 => 
                           n21470, ZN => n7138);
   U15050 : OAI22_X1 port map( A1 => n21478, A2 => n14299, B1 => n21640, B2 => 
                           n21470, ZN => n7139);
   U15051 : OAI22_X1 port map( A1 => n21478, A2 => n14298, B1 => n21643, B2 => 
                           n21470, ZN => n7140);
   U15052 : OAI22_X1 port map( A1 => n21478, A2 => n14297, B1 => n21646, B2 => 
                           n21470, ZN => n7141);
   U15053 : OAI22_X1 port map( A1 => n21478, A2 => n14296, B1 => n21649, B2 => 
                           n21470, ZN => n7142);
   U15054 : OAI22_X1 port map( A1 => n21478, A2 => n14295, B1 => n21652, B2 => 
                           n21470, ZN => n7143);
   U15055 : OAI22_X1 port map( A1 => n21478, A2 => n14294, B1 => n21655, B2 => 
                           n21470, ZN => n7144);
   U15056 : OAI22_X1 port map( A1 => n21478, A2 => n14293, B1 => n21658, B2 => 
                           n21470, ZN => n7145);
   U15057 : OAI22_X1 port map( A1 => n21478, A2 => n14292, B1 => n21661, B2 => 
                           n21470, ZN => n7146);
   U15058 : OAI22_X1 port map( A1 => n21478, A2 => n14291, B1 => n21664, B2 => 
                           n21470, ZN => n7147);
   U15059 : OAI22_X1 port map( A1 => n21478, A2 => n14290, B1 => n21667, B2 => 
                           n21470, ZN => n7148);
   U15060 : OAI22_X1 port map( A1 => n21478, A2 => n14289, B1 => n21670, B2 => 
                           n21471, ZN => n7149);
   U15061 : OAI22_X1 port map( A1 => n21478, A2 => n14288, B1 => n21673, B2 => 
                           n21471, ZN => n7150);
   U15062 : OAI22_X1 port map( A1 => n21478, A2 => n14287, B1 => n21676, B2 => 
                           n21471, ZN => n7151);
   U15063 : OAI22_X1 port map( A1 => n21479, A2 => n14286, B1 => n21679, B2 => 
                           n21471, ZN => n7152);
   U15064 : OAI22_X1 port map( A1 => n21479, A2 => n14285, B1 => n21682, B2 => 
                           n21471, ZN => n7153);
   U15065 : OAI22_X1 port map( A1 => n21479, A2 => n14284, B1 => n21685, B2 => 
                           n21471, ZN => n7154);
   U15066 : OAI22_X1 port map( A1 => n21479, A2 => n14283, B1 => n21688, B2 => 
                           n21471, ZN => n7155);
   U15067 : OAI22_X1 port map( A1 => n21479, A2 => n14282, B1 => n21691, B2 => 
                           n21471, ZN => n7156);
   U15068 : OAI22_X1 port map( A1 => n21479, A2 => n14281, B1 => n21694, B2 => 
                           n21471, ZN => n7157);
   U15069 : OAI22_X1 port map( A1 => n21479, A2 => n14280, B1 => n21697, B2 => 
                           n21471, ZN => n7158);
   U15070 : OAI22_X1 port map( A1 => n21479, A2 => n14279, B1 => n21700, B2 => 
                           n21471, ZN => n7159);
   U15071 : OAI22_X1 port map( A1 => n21479, A2 => n14278, B1 => n21703, B2 => 
                           n21471, ZN => n7160);
   U15072 : OAI22_X1 port map( A1 => n21488, A2 => n14271, B1 => n21526, B2 => 
                           n21480, ZN => n7165);
   U15073 : OAI22_X1 port map( A1 => n21488, A2 => n14270, B1 => n21529, B2 => 
                           n21480, ZN => n7166);
   U15074 : OAI22_X1 port map( A1 => n21488, A2 => n14269, B1 => n21532, B2 => 
                           n21480, ZN => n7167);
   U15075 : OAI22_X1 port map( A1 => n21488, A2 => n14268, B1 => n21535, B2 => 
                           n21480, ZN => n7168);
   U15076 : OAI22_X1 port map( A1 => n21488, A2 => n14267, B1 => n21538, B2 => 
                           n21480, ZN => n7169);
   U15077 : OAI22_X1 port map( A1 => n21488, A2 => n14266, B1 => n21541, B2 => 
                           n21480, ZN => n7170);
   U15078 : OAI22_X1 port map( A1 => n21488, A2 => n14265, B1 => n21544, B2 => 
                           n21480, ZN => n7171);
   U15079 : OAI22_X1 port map( A1 => n21488, A2 => n14264, B1 => n21547, B2 => 
                           n21480, ZN => n7172);
   U15080 : OAI22_X1 port map( A1 => n21488, A2 => n14263, B1 => n21550, B2 => 
                           n21480, ZN => n7173);
   U15081 : OAI22_X1 port map( A1 => n21488, A2 => n14262, B1 => n21553, B2 => 
                           n21480, ZN => n7174);
   U15082 : OAI22_X1 port map( A1 => n21488, A2 => n14261, B1 => n21556, B2 => 
                           n21480, ZN => n7175);
   U15083 : OAI22_X1 port map( A1 => n21488, A2 => n14260, B1 => n21559, B2 => 
                           n21480, ZN => n7176);
   U15084 : OAI22_X1 port map( A1 => n21489, A2 => n14259, B1 => n21562, B2 => 
                           n21481, ZN => n7177);
   U15085 : OAI22_X1 port map( A1 => n21489, A2 => n14258, B1 => n21565, B2 => 
                           n21481, ZN => n7178);
   U15086 : OAI22_X1 port map( A1 => n21489, A2 => n14257, B1 => n21568, B2 => 
                           n21481, ZN => n7179);
   U15087 : OAI22_X1 port map( A1 => n21489, A2 => n14256, B1 => n21571, B2 => 
                           n21481, ZN => n7180);
   U15088 : OAI22_X1 port map( A1 => n21489, A2 => n14255, B1 => n21574, B2 => 
                           n21481, ZN => n7181);
   U15089 : OAI22_X1 port map( A1 => n21489, A2 => n14254, B1 => n21577, B2 => 
                           n21481, ZN => n7182);
   U15090 : OAI22_X1 port map( A1 => n21489, A2 => n14253, B1 => n21580, B2 => 
                           n21481, ZN => n7183);
   U15091 : OAI22_X1 port map( A1 => n21489, A2 => n14252, B1 => n21583, B2 => 
                           n21481, ZN => n7184);
   U15092 : OAI22_X1 port map( A1 => n21489, A2 => n14251, B1 => n21586, B2 => 
                           n21481, ZN => n7185);
   U15093 : OAI22_X1 port map( A1 => n21489, A2 => n14250, B1 => n21589, B2 => 
                           n21481, ZN => n7186);
   U15094 : OAI22_X1 port map( A1 => n21489, A2 => n14249, B1 => n21592, B2 => 
                           n21481, ZN => n7187);
   U15095 : OAI22_X1 port map( A1 => n21489, A2 => n14248, B1 => n21595, B2 => 
                           n21481, ZN => n7188);
   U15096 : OAI22_X1 port map( A1 => n21489, A2 => n14247, B1 => n21598, B2 => 
                           n21482, ZN => n7189);
   U15097 : OAI22_X1 port map( A1 => n21490, A2 => n14246, B1 => n21601, B2 => 
                           n21482, ZN => n7190);
   U15098 : OAI22_X1 port map( A1 => n21490, A2 => n14245, B1 => n21604, B2 => 
                           n21482, ZN => n7191);
   U15099 : OAI22_X1 port map( A1 => n21490, A2 => n14244, B1 => n21607, B2 => 
                           n21482, ZN => n7192);
   U15100 : OAI22_X1 port map( A1 => n21490, A2 => n14243, B1 => n21610, B2 => 
                           n21482, ZN => n7193);
   U15101 : OAI22_X1 port map( A1 => n21490, A2 => n14242, B1 => n21613, B2 => 
                           n21482, ZN => n7194);
   U15102 : OAI22_X1 port map( A1 => n21490, A2 => n14241, B1 => n21616, B2 => 
                           n21482, ZN => n7195);
   U15103 : OAI22_X1 port map( A1 => n21490, A2 => n14240, B1 => n21619, B2 => 
                           n21482, ZN => n7196);
   U15104 : OAI22_X1 port map( A1 => n21490, A2 => n14239, B1 => n21622, B2 => 
                           n21482, ZN => n7197);
   U15105 : OAI22_X1 port map( A1 => n21490, A2 => n14238, B1 => n21625, B2 => 
                           n21482, ZN => n7198);
   U15106 : OAI22_X1 port map( A1 => n21490, A2 => n14237, B1 => n21628, B2 => 
                           n21482, ZN => n7199);
   U15107 : OAI22_X1 port map( A1 => n21490, A2 => n14236, B1 => n21631, B2 => 
                           n21482, ZN => n7200);
   U15108 : OAI22_X1 port map( A1 => n21490, A2 => n14235, B1 => n21634, B2 => 
                           n21483, ZN => n7201);
   U15109 : OAI22_X1 port map( A1 => n21490, A2 => n14234, B1 => n21637, B2 => 
                           n21483, ZN => n7202);
   U15110 : OAI22_X1 port map( A1 => n21491, A2 => n14233, B1 => n21640, B2 => 
                           n21483, ZN => n7203);
   U15111 : OAI22_X1 port map( A1 => n21491, A2 => n14232, B1 => n21643, B2 => 
                           n21483, ZN => n7204);
   U15112 : OAI22_X1 port map( A1 => n21491, A2 => n14231, B1 => n21646, B2 => 
                           n21483, ZN => n7205);
   U15113 : OAI22_X1 port map( A1 => n21491, A2 => n14230, B1 => n21649, B2 => 
                           n21483, ZN => n7206);
   U15114 : OAI22_X1 port map( A1 => n21491, A2 => n14229, B1 => n21652, B2 => 
                           n21483, ZN => n7207);
   U15115 : OAI22_X1 port map( A1 => n21491, A2 => n14228, B1 => n21655, B2 => 
                           n21483, ZN => n7208);
   U15116 : OAI22_X1 port map( A1 => n21491, A2 => n14227, B1 => n21658, B2 => 
                           n21483, ZN => n7209);
   U15117 : OAI22_X1 port map( A1 => n21491, A2 => n14226, B1 => n21661, B2 => 
                           n21483, ZN => n7210);
   U15118 : OAI22_X1 port map( A1 => n21491, A2 => n14225, B1 => n21664, B2 => 
                           n21483, ZN => n7211);
   U15119 : OAI22_X1 port map( A1 => n21491, A2 => n14224, B1 => n21667, B2 => 
                           n21483, ZN => n7212);
   U15120 : OAI22_X1 port map( A1 => n21491, A2 => n14223, B1 => n21670, B2 => 
                           n21484, ZN => n7213);
   U15121 : OAI22_X1 port map( A1 => n21491, A2 => n14222, B1 => n21673, B2 => 
                           n21484, ZN => n7214);
   U15122 : OAI22_X1 port map( A1 => n21491, A2 => n14221, B1 => n21676, B2 => 
                           n21484, ZN => n7215);
   U15123 : OAI22_X1 port map( A1 => n21492, A2 => n14220, B1 => n21679, B2 => 
                           n21484, ZN => n7216);
   U15124 : OAI22_X1 port map( A1 => n21492, A2 => n14219, B1 => n21682, B2 => 
                           n21484, ZN => n7217);
   U15125 : OAI22_X1 port map( A1 => n21492, A2 => n14218, B1 => n21685, B2 => 
                           n21484, ZN => n7218);
   U15126 : OAI22_X1 port map( A1 => n21492, A2 => n14217, B1 => n21688, B2 => 
                           n21484, ZN => n7219);
   U15127 : OAI22_X1 port map( A1 => n21492, A2 => n14216, B1 => n21691, B2 => 
                           n21484, ZN => n7220);
   U15128 : OAI22_X1 port map( A1 => n21492, A2 => n14215, B1 => n21694, B2 => 
                           n21484, ZN => n7221);
   U15129 : OAI22_X1 port map( A1 => n21492, A2 => n14214, B1 => n21697, B2 => 
                           n21484, ZN => n7222);
   U15130 : OAI22_X1 port map( A1 => n21492, A2 => n14213, B1 => n21700, B2 => 
                           n21484, ZN => n7223);
   U15131 : OAI22_X1 port map( A1 => n21492, A2 => n14212, B1 => n21703, B2 => 
                           n21484, ZN => n7224);
   U15132 : OAI22_X1 port map( A1 => n21514, A2 => n14137, B1 => n21526, B2 => 
                           n21506, ZN => n7293);
   U15133 : OAI22_X1 port map( A1 => n21514, A2 => n14136, B1 => n21529, B2 => 
                           n21506, ZN => n7294);
   U15134 : OAI22_X1 port map( A1 => n21514, A2 => n14135, B1 => n21532, B2 => 
                           n21506, ZN => n7295);
   U15135 : OAI22_X1 port map( A1 => n21514, A2 => n14134, B1 => n21535, B2 => 
                           n21506, ZN => n7296);
   U15136 : OAI22_X1 port map( A1 => n21514, A2 => n14133, B1 => n21538, B2 => 
                           n21506, ZN => n7297);
   U15137 : OAI22_X1 port map( A1 => n21514, A2 => n14132, B1 => n21541, B2 => 
                           n21506, ZN => n7298);
   U15138 : OAI22_X1 port map( A1 => n21514, A2 => n14131, B1 => n21544, B2 => 
                           n21506, ZN => n7299);
   U15139 : OAI22_X1 port map( A1 => n21514, A2 => n14130, B1 => n21547, B2 => 
                           n21506, ZN => n7300);
   U15140 : OAI22_X1 port map( A1 => n21514, A2 => n14129, B1 => n21550, B2 => 
                           n21506, ZN => n7301);
   U15141 : OAI22_X1 port map( A1 => n21514, A2 => n14128, B1 => n21553, B2 => 
                           n21506, ZN => n7302);
   U15142 : OAI22_X1 port map( A1 => n21514, A2 => n14127, B1 => n21556, B2 => 
                           n21506, ZN => n7303);
   U15143 : OAI22_X1 port map( A1 => n21514, A2 => n14126, B1 => n21559, B2 => 
                           n21506, ZN => n7304);
   U15144 : OAI22_X1 port map( A1 => n21515, A2 => n14125, B1 => n21562, B2 => 
                           n21507, ZN => n7305);
   U15145 : OAI22_X1 port map( A1 => n21515, A2 => n14124, B1 => n21565, B2 => 
                           n21507, ZN => n7306);
   U15146 : OAI22_X1 port map( A1 => n21515, A2 => n14123, B1 => n21568, B2 => 
                           n21507, ZN => n7307);
   U15147 : OAI22_X1 port map( A1 => n21515, A2 => n14122, B1 => n21571, B2 => 
                           n21507, ZN => n7308);
   U15148 : OAI22_X1 port map( A1 => n21515, A2 => n14121, B1 => n21574, B2 => 
                           n21507, ZN => n7309);
   U15149 : OAI22_X1 port map( A1 => n21515, A2 => n14120, B1 => n21577, B2 => 
                           n21507, ZN => n7310);
   U15150 : OAI22_X1 port map( A1 => n21515, A2 => n14119, B1 => n21580, B2 => 
                           n21507, ZN => n7311);
   U15151 : OAI22_X1 port map( A1 => n21515, A2 => n14118, B1 => n21583, B2 => 
                           n21507, ZN => n7312);
   U15152 : OAI22_X1 port map( A1 => n21515, A2 => n14117, B1 => n21586, B2 => 
                           n21507, ZN => n7313);
   U15153 : OAI22_X1 port map( A1 => n21515, A2 => n14116, B1 => n21589, B2 => 
                           n21507, ZN => n7314);
   U15154 : OAI22_X1 port map( A1 => n21515, A2 => n14115, B1 => n21592, B2 => 
                           n21507, ZN => n7315);
   U15155 : OAI22_X1 port map( A1 => n21515, A2 => n14114, B1 => n21595, B2 => 
                           n21507, ZN => n7316);
   U15156 : OAI22_X1 port map( A1 => n21515, A2 => n14113, B1 => n21598, B2 => 
                           n21508, ZN => n7317);
   U15157 : OAI22_X1 port map( A1 => n21516, A2 => n14112, B1 => n21601, B2 => 
                           n21508, ZN => n7318);
   U15158 : OAI22_X1 port map( A1 => n21516, A2 => n14111, B1 => n21604, B2 => 
                           n21508, ZN => n7319);
   U15159 : OAI22_X1 port map( A1 => n21516, A2 => n14110, B1 => n21607, B2 => 
                           n21508, ZN => n7320);
   U15160 : OAI22_X1 port map( A1 => n21516, A2 => n14109, B1 => n21610, B2 => 
                           n21508, ZN => n7321);
   U15161 : OAI22_X1 port map( A1 => n21516, A2 => n14108, B1 => n21613, B2 => 
                           n21508, ZN => n7322);
   U15162 : OAI22_X1 port map( A1 => n21516, A2 => n14107, B1 => n21616, B2 => 
                           n21508, ZN => n7323);
   U15163 : OAI22_X1 port map( A1 => n21516, A2 => n14106, B1 => n21619, B2 => 
                           n21508, ZN => n7324);
   U15164 : OAI22_X1 port map( A1 => n21516, A2 => n14105, B1 => n21622, B2 => 
                           n21508, ZN => n7325);
   U15165 : OAI22_X1 port map( A1 => n21516, A2 => n14104, B1 => n21625, B2 => 
                           n21508, ZN => n7326);
   U15166 : OAI22_X1 port map( A1 => n21516, A2 => n14103, B1 => n21628, B2 => 
                           n21508, ZN => n7327);
   U15167 : OAI22_X1 port map( A1 => n21516, A2 => n14102, B1 => n21631, B2 => 
                           n21508, ZN => n7328);
   U15168 : OAI22_X1 port map( A1 => n21516, A2 => n14101, B1 => n21634, B2 => 
                           n21509, ZN => n7329);
   U15169 : OAI22_X1 port map( A1 => n21516, A2 => n14100, B1 => n21637, B2 => 
                           n21509, ZN => n7330);
   U15170 : OAI22_X1 port map( A1 => n21517, A2 => n14099, B1 => n21640, B2 => 
                           n21509, ZN => n7331);
   U15171 : OAI22_X1 port map( A1 => n21517, A2 => n14098, B1 => n21643, B2 => 
                           n21509, ZN => n7332);
   U15172 : OAI22_X1 port map( A1 => n21517, A2 => n14097, B1 => n21646, B2 => 
                           n21509, ZN => n7333);
   U15173 : OAI22_X1 port map( A1 => n21517, A2 => n14096, B1 => n21649, B2 => 
                           n21509, ZN => n7334);
   U15174 : OAI22_X1 port map( A1 => n21517, A2 => n14095, B1 => n21652, B2 => 
                           n21509, ZN => n7335);
   U15175 : OAI22_X1 port map( A1 => n21517, A2 => n14094, B1 => n21655, B2 => 
                           n21509, ZN => n7336);
   U15176 : OAI22_X1 port map( A1 => n21517, A2 => n14093, B1 => n21658, B2 => 
                           n21509, ZN => n7337);
   U15177 : OAI22_X1 port map( A1 => n21517, A2 => n14092, B1 => n21661, B2 => 
                           n21509, ZN => n7338);
   U15178 : OAI22_X1 port map( A1 => n21517, A2 => n14091, B1 => n21664, B2 => 
                           n21509, ZN => n7339);
   U15179 : OAI22_X1 port map( A1 => n21517, A2 => n14090, B1 => n21667, B2 => 
                           n21509, ZN => n7340);
   U15180 : OAI22_X1 port map( A1 => n21517, A2 => n14089, B1 => n21670, B2 => 
                           n21510, ZN => n7341);
   U15181 : OAI22_X1 port map( A1 => n21517, A2 => n14088, B1 => n21673, B2 => 
                           n21510, ZN => n7342);
   U15182 : OAI22_X1 port map( A1 => n21517, A2 => n14087, B1 => n21676, B2 => 
                           n21510, ZN => n7343);
   U15183 : OAI22_X1 port map( A1 => n21518, A2 => n14086, B1 => n21679, B2 => 
                           n21510, ZN => n7344);
   U15184 : OAI22_X1 port map( A1 => n21518, A2 => n14085, B1 => n21682, B2 => 
                           n21510, ZN => n7345);
   U15185 : OAI22_X1 port map( A1 => n21518, A2 => n14084, B1 => n21685, B2 => 
                           n21510, ZN => n7346);
   U15186 : OAI22_X1 port map( A1 => n21518, A2 => n14083, B1 => n21688, B2 => 
                           n21510, ZN => n7347);
   U15187 : OAI22_X1 port map( A1 => n21518, A2 => n14082, B1 => n21691, B2 => 
                           n21510, ZN => n7348);
   U15188 : OAI22_X1 port map( A1 => n21518, A2 => n14081, B1 => n21694, B2 => 
                           n21510, ZN => n7349);
   U15189 : OAI22_X1 port map( A1 => n21518, A2 => n14080, B1 => n21697, B2 => 
                           n21510, ZN => n7350);
   U15190 : OAI22_X1 port map( A1 => n21518, A2 => n14079, B1 => n21700, B2 => 
                           n21510, ZN => n7351);
   U15191 : OAI22_X1 port map( A1 => n21518, A2 => n14078, B1 => n21703, B2 => 
                           n21510, ZN => n7352);
   U15192 : NAND2_X1 port map( A1 => n17315, A2 => n17320, ZN => n16087);
   U15193 : OAI21_X1 port map( B1 => n14138, B2 => n14471, A => n21523, ZN => 
                           n14475);
   U15194 : OAI21_X1 port map( B1 => n14138, B2 => n14338, A => n21522, ZN => 
                           n14339);
   U15195 : OAI21_X1 port map( B1 => n14138, B2 => n14205, A => n21521, ZN => 
                           n14206);
   U15196 : OAI21_X1 port map( B1 => n14070, B2 => n14471, A => n21522, ZN => 
                           n14405);
   U15197 : OAI21_X1 port map( B1 => n14070, B2 => n14338, A => n21522, ZN => 
                           n14272);
   U15198 : OAI21_X1 port map( B1 => n14070, B2 => n14205, A => n21521, ZN => 
                           n14139);
   U15199 : BUF_X1 port map( A => n14068, Z => n21528);
   U15200 : BUF_X1 port map( A => n14066, Z => n21531);
   U15201 : BUF_X1 port map( A => n14064, Z => n21534);
   U15202 : BUF_X1 port map( A => n14062, Z => n21537);
   U15203 : BUF_X1 port map( A => n14060, Z => n21540);
   U15204 : BUF_X1 port map( A => n14058, Z => n21543);
   U15205 : BUF_X1 port map( A => n14056, Z => n21546);
   U15206 : BUF_X1 port map( A => n14054, Z => n21549);
   U15207 : BUF_X1 port map( A => n14052, Z => n21552);
   U15208 : BUF_X1 port map( A => n14050, Z => n21555);
   U15209 : BUF_X1 port map( A => n14048, Z => n21558);
   U15210 : BUF_X1 port map( A => n14046, Z => n21561);
   U15211 : BUF_X1 port map( A => n14044, Z => n21564);
   U15212 : BUF_X1 port map( A => n14042, Z => n21567);
   U15213 : BUF_X1 port map( A => n14040, Z => n21570);
   U15214 : BUF_X1 port map( A => n14038, Z => n21573);
   U15215 : BUF_X1 port map( A => n14036, Z => n21576);
   U15216 : BUF_X1 port map( A => n14034, Z => n21579);
   U15217 : BUF_X1 port map( A => n14032, Z => n21582);
   U15218 : BUF_X1 port map( A => n14030, Z => n21585);
   U15219 : BUF_X1 port map( A => n14028, Z => n21588);
   U15220 : BUF_X1 port map( A => n14026, Z => n21591);
   U15221 : BUF_X1 port map( A => n14024, Z => n21594);
   U15222 : BUF_X1 port map( A => n14022, Z => n21597);
   U15223 : BUF_X1 port map( A => n14020, Z => n21600);
   U15224 : BUF_X1 port map( A => n14018, Z => n21603);
   U15225 : BUF_X1 port map( A => n14016, Z => n21606);
   U15226 : BUF_X1 port map( A => n14014, Z => n21609);
   U15227 : BUF_X1 port map( A => n14012, Z => n21612);
   U15228 : BUF_X1 port map( A => n14010, Z => n21615);
   U15229 : BUF_X1 port map( A => n14008, Z => n21618);
   U15230 : BUF_X1 port map( A => n14006, Z => n21621);
   U15231 : BUF_X1 port map( A => n14004, Z => n21624);
   U15232 : BUF_X1 port map( A => n14002, Z => n21627);
   U15233 : BUF_X1 port map( A => n14000, Z => n21630);
   U15234 : BUF_X1 port map( A => n13998, Z => n21633);
   U15235 : BUF_X1 port map( A => n13996, Z => n21636);
   U15236 : BUF_X1 port map( A => n13994, Z => n21639);
   U15237 : BUF_X1 port map( A => n13992, Z => n21642);
   U15238 : BUF_X1 port map( A => n13990, Z => n21645);
   U15239 : BUF_X1 port map( A => n13988, Z => n21648);
   U15240 : BUF_X1 port map( A => n13986, Z => n21651);
   U15241 : BUF_X1 port map( A => n13984, Z => n21654);
   U15242 : BUF_X1 port map( A => n13982, Z => n21657);
   U15243 : BUF_X1 port map( A => n13980, Z => n21660);
   U15244 : BUF_X1 port map( A => n13978, Z => n21663);
   U15245 : BUF_X1 port map( A => n13976, Z => n21666);
   U15246 : BUF_X1 port map( A => n13974, Z => n21669);
   U15247 : BUF_X1 port map( A => n13972, Z => n21672);
   U15248 : BUF_X1 port map( A => n13970, Z => n21675);
   U15249 : BUF_X1 port map( A => n13968, Z => n21678);
   U15250 : BUF_X1 port map( A => n13966, Z => n21681);
   U15251 : BUF_X1 port map( A => n13964, Z => n21684);
   U15252 : BUF_X1 port map( A => n13962, Z => n21687);
   U15253 : BUF_X1 port map( A => n13960, Z => n21690);
   U15254 : BUF_X1 port map( A => n13958, Z => n21693);
   U15255 : BUF_X1 port map( A => n13956, Z => n21696);
   U15256 : BUF_X1 port map( A => n13954, Z => n21699);
   U15257 : BUF_X1 port map( A => n13952, Z => n21702);
   U15258 : BUF_X1 port map( A => n13950, Z => n21705);
   U15259 : BUF_X1 port map( A => n13948, Z => n21708);
   U15260 : BUF_X1 port map( A => n13946, Z => n21711);
   U15261 : BUF_X1 port map( A => n13944, Z => n21714);
   U15262 : BUF_X1 port map( A => n13942, Z => n21717);
   U15263 : OAI21_X1 port map( B1 => n14471, B2 => n15736, A => n21521, ZN => 
                           n16069);
   U15264 : OAI21_X1 port map( B1 => n14471, B2 => n15669, A => n21521, ZN => 
                           n16003);
   U15265 : OAI21_X1 port map( B1 => n14338, B2 => n15736, A => n21521, ZN => 
                           n15937);
   U15266 : OAI21_X1 port map( B1 => n14338, B2 => n15669, A => n21521, ZN => 
                           n15871);
   U15267 : OAI21_X1 port map( B1 => n14205, B2 => n15736, A => n21521, ZN => 
                           n15805);
   U15268 : OAI21_X1 port map( B1 => n14205, B2 => n15669, A => n21521, ZN => 
                           n15739);
   U15269 : OAI21_X1 port map( B1 => n14071, B2 => n15736, A => n21521, ZN => 
                           n15670);
   U15270 : OAI21_X1 port map( B1 => n14071, B2 => n15669, A => n21521, ZN => 
                           n15603);
   U15271 : OAI21_X1 port map( B1 => n14471, B2 => n15205, A => n21522, ZN => 
                           n15537);
   U15272 : OAI21_X1 port map( B1 => n14471, B2 => n15138, A => n21522, ZN => 
                           n15470);
   U15273 : OAI21_X1 port map( B1 => n14338, B2 => n15205, A => n21522, ZN => 
                           n15404);
   U15274 : OAI21_X1 port map( B1 => n14338, B2 => n15138, A => n21522, ZN => 
                           n15338);
   U15275 : OAI21_X1 port map( B1 => n14205, B2 => n15205, A => n21522, ZN => 
                           n15272);
   U15276 : OAI21_X1 port map( B1 => n14205, B2 => n15138, A => n21522, ZN => 
                           n15206);
   U15277 : OAI21_X1 port map( B1 => n14071, B2 => n15205, A => n21522, ZN => 
                           n15139);
   U15278 : OAI21_X1 port map( B1 => n14471, B2 => n14607, A => n21523, ZN => 
                           n14939);
   U15279 : OAI21_X1 port map( B1 => n14338, B2 => n14607, A => n21523, ZN => 
                           n14807);
   U15280 : OAI21_X1 port map( B1 => n14205, B2 => n14607, A => n21523, ZN => 
                           n14675);
   U15281 : OAI21_X1 port map( B1 => n14071, B2 => n14607, A => n21523, ZN => 
                           n14541);
   U15282 : OAI21_X1 port map( B1 => n14471, B2 => n14674, A => n21523, ZN => 
                           n15005);
   U15283 : OAI21_X1 port map( B1 => n14338, B2 => n14674, A => n21522, ZN => 
                           n14873);
   U15284 : OAI21_X1 port map( B1 => n14205, B2 => n14674, A => n21523, ZN => 
                           n14741);
   U15285 : OAI21_X1 port map( B1 => n14071, B2 => n14674, A => n21522, ZN => 
                           n14608);
   U15286 : OAI21_X1 port map( B1 => n14071, B2 => n14138, A => n21521, ZN => 
                           n14072);
   U15287 : AND2_X1 port map( A1 => n18514, A2 => n18513, ZN => n17363);
   U15288 : AND2_X1 port map( A1 => n18514, A2 => n18515, ZN => n17348);
   U15289 : AND2_X1 port map( A1 => n17313, A2 => n17312, ZN => n16097);
   U15290 : AND2_X1 port map( A1 => n17313, A2 => n17314, ZN => n16081);
   U15291 : AND2_X1 port map( A1 => n18512, A2 => n18513, ZN => n17349);
   U15292 : AND2_X1 port map( A1 => n18512, A2 => n18524, ZN => n17377);
   U15293 : AND2_X1 port map( A1 => n17311, A2 => n17312, ZN => n16082);
   U15294 : AND2_X1 port map( A1 => n17311, A2 => n17323, ZN => n16112);
   U15295 : AND2_X1 port map( A1 => n17320, A2 => n17314, ZN => n16098);
   U15296 : AND2_X1 port map( A1 => n18531, A2 => n18513, ZN => n17373);
   U15297 : AND2_X1 port map( A1 => n18531, A2 => n18516, ZN => n17378);
   U15298 : AND2_X1 port map( A1 => n18531, A2 => n18521, ZN => n17388);
   U15299 : AND2_X1 port map( A1 => n18531, A2 => n18515, ZN => n17387);
   U15300 : AND2_X1 port map( A1 => n17330, A2 => n17312, ZN => n16107);
   U15301 : AND2_X1 port map( A1 => n17330, A2 => n17315, ZN => n16113);
   U15302 : AND2_X1 port map( A1 => n17330, A2 => n17318, ZN => n16123);
   U15303 : AND2_X1 port map( A1 => n17330, A2 => n17314, ZN => n16122);
   U15304 : AND2_X1 port map( A1 => n18520, A2 => n18515, ZN => n17364);
   U15305 : AND2_X1 port map( A1 => n18519, A2 => n18514, ZN => n17354);
   U15306 : AND2_X1 port map( A1 => n18521, A2 => n18512, ZN => n17383);
   U15307 : AND2_X1 port map( A1 => n17318, A2 => n17311, ZN => n16118);
   U15308 : AND2_X1 port map( A1 => n17312, A2 => n17320, ZN => n16099);
   U15309 : AND2_X1 port map( A1 => n17318, A2 => n17320, ZN => n16093);
   U15310 : AND2_X1 port map( A1 => n17319, A2 => n17320, ZN => n16092);
   U15311 : AND2_X1 port map( A1 => n17323, A2 => n17320, ZN => n16117);
   U15312 : AND2_X1 port map( A1 => n18513, A2 => n18520, ZN => n17365);
   U15313 : AND2_X1 port map( A1 => n18521, A2 => n18520, ZN => n17359);
   U15314 : AND2_X1 port map( A1 => n18519, A2 => n18520, ZN => n17358);
   U15315 : AND2_X1 port map( A1 => n18516, A2 => n18520, ZN => n17353);
   U15316 : AND2_X1 port map( A1 => n18524, A2 => n18520, ZN => n17382);
   U15317 : NAND2_X1 port map( A1 => n15071, A2 => n21521, ZN => n16108);
   U15318 : BUF_X1 port map( A => n14069, Z => n21519);
   U15319 : NAND2_X1 port map( A1 => n16163, A2 => n16164, ZN => n5429);
   U15320 : NOR4_X1 port map( A1 => n16173, A2 => n16174, A3 => n16175, A4 => 
                           n16176, ZN => n16163);
   U15321 : NOR4_X1 port map( A1 => n16165, A2 => n16166, A3 => n16167, A4 => 
                           n16168, ZN => n16164);
   U15322 : OAI221_X1 port map( B1 => n14480, B2 => n20933, C1 => n15876, C2 =>
                           n20927, A => n16180, ZN => n16173);
   U15323 : NAND2_X1 port map( A1 => n16144, A2 => n16145, ZN => n5431);
   U15324 : NOR4_X1 port map( A1 => n16154, A2 => n16155, A3 => n16156, A4 => 
                           n16157, ZN => n16144);
   U15325 : NOR4_X1 port map( A1 => n16146, A2 => n16147, A3 => n16148, A4 => 
                           n16149, ZN => n16145);
   U15326 : OAI221_X1 port map( B1 => n14479, B2 => n20933, C1 => n15875, C2 =>
                           n20927, A => n16161, ZN => n16154);
   U15327 : NAND2_X1 port map( A1 => n16125, A2 => n16126, ZN => n5433);
   U15328 : NOR4_X1 port map( A1 => n16135, A2 => n16136, A3 => n16137, A4 => 
                           n16138, ZN => n16125);
   U15329 : NOR4_X1 port map( A1 => n16127, A2 => n16128, A3 => n16129, A4 => 
                           n16130, ZN => n16126);
   U15330 : OAI221_X1 port map( B1 => n14478, B2 => n20933, C1 => n15874, C2 =>
                           n20927, A => n16142, ZN => n16135);
   U15331 : NAND2_X1 port map( A1 => n16072, A2 => n16073, ZN => n5435);
   U15332 : NOR4_X1 port map( A1 => n16100, A2 => n16101, A3 => n16102, A4 => 
                           n16103, ZN => n16072);
   U15333 : NOR4_X1 port map( A1 => n16074, A2 => n16075, A3 => n16076, A4 => 
                           n16077, ZN => n16073);
   U15334 : OAI221_X1 port map( B1 => n14476, B2 => n20933, C1 => n15872, C2 =>
                           n20927, A => n16121, ZN => n16100);
   U15335 : NAND2_X1 port map( A1 => n18505, A2 => n18506, ZN => n5245);
   U15336 : NOR4_X1 port map( A1 => n18526, A2 => n18527, A3 => n18528, A4 => 
                           n18529, ZN => n18505);
   U15337 : NOR4_X1 port map( A1 => n18507, A2 => n18508, A3 => n18509, A4 => 
                           n18510, ZN => n18506);
   U15338 : OAI221_X1 port map( B1 => n14540, B2 => n20736, C1 => n15936, C2 =>
                           n20730, A => n18537, ZN => n18526);
   U15339 : NAND2_X1 port map( A1 => n18487, A2 => n18488, ZN => n5246);
   U15340 : NOR4_X1 port map( A1 => n18497, A2 => n18498, A3 => n18499, A4 => 
                           n18500, ZN => n18487);
   U15341 : NOR4_X1 port map( A1 => n18489, A2 => n18490, A3 => n18491, A4 => 
                           n18492, ZN => n18488);
   U15342 : OAI221_X1 port map( B1 => n14539, B2 => n20736, C1 => n15935, C2 =>
                           n20730, A => n18504, ZN => n18497);
   U15343 : NAND2_X1 port map( A1 => n18469, A2 => n18470, ZN => n5247);
   U15344 : NOR4_X1 port map( A1 => n18479, A2 => n18480, A3 => n18481, A4 => 
                           n18482, ZN => n18469);
   U15345 : NOR4_X1 port map( A1 => n18471, A2 => n18472, A3 => n18473, A4 => 
                           n18474, ZN => n18470);
   U15346 : OAI221_X1 port map( B1 => n14538, B2 => n20736, C1 => n15934, C2 =>
                           n20730, A => n18486, ZN => n18479);
   U15347 : NAND2_X1 port map( A1 => n18451, A2 => n18452, ZN => n5248);
   U15348 : NOR4_X1 port map( A1 => n18461, A2 => n18462, A3 => n18463, A4 => 
                           n18464, ZN => n18451);
   U15349 : NOR4_X1 port map( A1 => n18453, A2 => n18454, A3 => n18455, A4 => 
                           n18456, ZN => n18452);
   U15350 : OAI221_X1 port map( B1 => n14537, B2 => n20736, C1 => n15933, C2 =>
                           n20730, A => n18468, ZN => n18461);
   U15351 : NAND2_X1 port map( A1 => n18433, A2 => n18434, ZN => n5249);
   U15352 : NOR4_X1 port map( A1 => n18443, A2 => n18444, A3 => n18445, A4 => 
                           n18446, ZN => n18433);
   U15353 : NOR4_X1 port map( A1 => n18435, A2 => n18436, A3 => n18437, A4 => 
                           n18438, ZN => n18434);
   U15354 : OAI221_X1 port map( B1 => n14536, B2 => n20736, C1 => n15932, C2 =>
                           n20730, A => n18450, ZN => n18443);
   U15355 : NAND2_X1 port map( A1 => n18415, A2 => n18416, ZN => n5250);
   U15356 : NOR4_X1 port map( A1 => n18425, A2 => n18426, A3 => n18427, A4 => 
                           n18428, ZN => n18415);
   U15357 : NOR4_X1 port map( A1 => n18417, A2 => n18418, A3 => n18419, A4 => 
                           n18420, ZN => n18416);
   U15358 : OAI221_X1 port map( B1 => n14535, B2 => n20736, C1 => n15931, C2 =>
                           n20730, A => n18432, ZN => n18425);
   U15359 : NAND2_X1 port map( A1 => n18397, A2 => n18398, ZN => n5251);
   U15360 : NOR4_X1 port map( A1 => n18407, A2 => n18408, A3 => n18409, A4 => 
                           n18410, ZN => n18397);
   U15361 : NOR4_X1 port map( A1 => n18399, A2 => n18400, A3 => n18401, A4 => 
                           n18402, ZN => n18398);
   U15362 : OAI221_X1 port map( B1 => n14534, B2 => n20736, C1 => n15930, C2 =>
                           n20730, A => n18414, ZN => n18407);
   U15363 : NAND2_X1 port map( A1 => n18379, A2 => n18380, ZN => n5252);
   U15364 : NOR4_X1 port map( A1 => n18389, A2 => n18390, A3 => n18391, A4 => 
                           n18392, ZN => n18379);
   U15365 : NOR4_X1 port map( A1 => n18381, A2 => n18382, A3 => n18383, A4 => 
                           n18384, ZN => n18380);
   U15366 : OAI221_X1 port map( B1 => n14533, B2 => n20736, C1 => n15929, C2 =>
                           n20730, A => n18396, ZN => n18389);
   U15367 : NAND2_X1 port map( A1 => n18361, A2 => n18362, ZN => n5253);
   U15368 : NOR4_X1 port map( A1 => n18371, A2 => n18372, A3 => n18373, A4 => 
                           n18374, ZN => n18361);
   U15369 : NOR4_X1 port map( A1 => n18363, A2 => n18364, A3 => n18365, A4 => 
                           n18366, ZN => n18362);
   U15370 : OAI221_X1 port map( B1 => n14532, B2 => n20736, C1 => n15928, C2 =>
                           n20730, A => n18378, ZN => n18371);
   U15371 : NAND2_X1 port map( A1 => n18343, A2 => n18344, ZN => n5254);
   U15372 : NOR4_X1 port map( A1 => n18353, A2 => n18354, A3 => n18355, A4 => 
                           n18356, ZN => n18343);
   U15373 : NOR4_X1 port map( A1 => n18345, A2 => n18346, A3 => n18347, A4 => 
                           n18348, ZN => n18344);
   U15374 : OAI221_X1 port map( B1 => n14531, B2 => n20736, C1 => n15927, C2 =>
                           n20730, A => n18360, ZN => n18353);
   U15375 : NAND2_X1 port map( A1 => n18325, A2 => n18326, ZN => n5255);
   U15376 : NOR4_X1 port map( A1 => n18335, A2 => n18336, A3 => n18337, A4 => 
                           n18338, ZN => n18325);
   U15377 : NOR4_X1 port map( A1 => n18327, A2 => n18328, A3 => n18329, A4 => 
                           n18330, ZN => n18326);
   U15378 : OAI221_X1 port map( B1 => n14530, B2 => n20736, C1 => n15926, C2 =>
                           n20730, A => n18342, ZN => n18335);
   U15379 : NAND2_X1 port map( A1 => n18307, A2 => n18308, ZN => n5256);
   U15380 : NOR4_X1 port map( A1 => n18317, A2 => n18318, A3 => n18319, A4 => 
                           n18320, ZN => n18307);
   U15381 : NOR4_X1 port map( A1 => n18309, A2 => n18310, A3 => n18311, A4 => 
                           n18312, ZN => n18308);
   U15382 : OAI221_X1 port map( B1 => n14529, B2 => n20736, C1 => n15925, C2 =>
                           n20730, A => n18324, ZN => n18317);
   U15383 : NAND2_X1 port map( A1 => n18289, A2 => n18290, ZN => n5257);
   U15384 : NOR4_X1 port map( A1 => n18299, A2 => n18300, A3 => n18301, A4 => 
                           n18302, ZN => n18289);
   U15385 : NOR4_X1 port map( A1 => n18291, A2 => n18292, A3 => n18293, A4 => 
                           n18294, ZN => n18290);
   U15386 : OAI221_X1 port map( B1 => n14528, B2 => n20737, C1 => n15924, C2 =>
                           n20731, A => n18306, ZN => n18299);
   U15387 : NAND2_X1 port map( A1 => n18271, A2 => n18272, ZN => n5258);
   U15388 : NOR4_X1 port map( A1 => n18281, A2 => n18282, A3 => n18283, A4 => 
                           n18284, ZN => n18271);
   U15389 : NOR4_X1 port map( A1 => n18273, A2 => n18274, A3 => n18275, A4 => 
                           n18276, ZN => n18272);
   U15390 : OAI221_X1 port map( B1 => n14527, B2 => n20737, C1 => n15923, C2 =>
                           n20731, A => n18288, ZN => n18281);
   U15391 : NAND2_X1 port map( A1 => n18253, A2 => n18254, ZN => n5259);
   U15392 : NOR4_X1 port map( A1 => n18263, A2 => n18264, A3 => n18265, A4 => 
                           n18266, ZN => n18253);
   U15393 : NOR4_X1 port map( A1 => n18255, A2 => n18256, A3 => n18257, A4 => 
                           n18258, ZN => n18254);
   U15394 : OAI221_X1 port map( B1 => n14526, B2 => n20737, C1 => n15922, C2 =>
                           n20731, A => n18270, ZN => n18263);
   U15395 : NAND2_X1 port map( A1 => n18235, A2 => n18236, ZN => n5260);
   U15396 : NOR4_X1 port map( A1 => n18245, A2 => n18246, A3 => n18247, A4 => 
                           n18248, ZN => n18235);
   U15397 : NOR4_X1 port map( A1 => n18237, A2 => n18238, A3 => n18239, A4 => 
                           n18240, ZN => n18236);
   U15398 : OAI221_X1 port map( B1 => n14525, B2 => n20737, C1 => n15921, C2 =>
                           n20731, A => n18252, ZN => n18245);
   U15399 : NAND2_X1 port map( A1 => n18217, A2 => n18218, ZN => n5261);
   U15400 : NOR4_X1 port map( A1 => n18227, A2 => n18228, A3 => n18229, A4 => 
                           n18230, ZN => n18217);
   U15401 : NOR4_X1 port map( A1 => n18219, A2 => n18220, A3 => n18221, A4 => 
                           n18222, ZN => n18218);
   U15402 : OAI221_X1 port map( B1 => n14524, B2 => n20737, C1 => n15920, C2 =>
                           n20731, A => n18234, ZN => n18227);
   U15403 : NAND2_X1 port map( A1 => n18199, A2 => n18200, ZN => n5262);
   U15404 : NOR4_X1 port map( A1 => n18209, A2 => n18210, A3 => n18211, A4 => 
                           n18212, ZN => n18199);
   U15405 : NOR4_X1 port map( A1 => n18201, A2 => n18202, A3 => n18203, A4 => 
                           n18204, ZN => n18200);
   U15406 : OAI221_X1 port map( B1 => n14523, B2 => n20737, C1 => n15919, C2 =>
                           n20731, A => n18216, ZN => n18209);
   U15407 : NAND2_X1 port map( A1 => n18181, A2 => n18182, ZN => n5263);
   U15408 : NOR4_X1 port map( A1 => n18191, A2 => n18192, A3 => n18193, A4 => 
                           n18194, ZN => n18181);
   U15409 : NOR4_X1 port map( A1 => n18183, A2 => n18184, A3 => n18185, A4 => 
                           n18186, ZN => n18182);
   U15410 : OAI221_X1 port map( B1 => n14522, B2 => n20737, C1 => n15918, C2 =>
                           n20731, A => n18198, ZN => n18191);
   U15411 : NAND2_X1 port map( A1 => n18163, A2 => n18164, ZN => n5264);
   U15412 : NOR4_X1 port map( A1 => n18173, A2 => n18174, A3 => n18175, A4 => 
                           n18176, ZN => n18163);
   U15413 : NOR4_X1 port map( A1 => n18165, A2 => n18166, A3 => n18167, A4 => 
                           n18168, ZN => n18164);
   U15414 : OAI221_X1 port map( B1 => n14521, B2 => n20737, C1 => n15917, C2 =>
                           n20731, A => n18180, ZN => n18173);
   U15415 : NAND2_X1 port map( A1 => n18145, A2 => n18146, ZN => n5265);
   U15416 : NOR4_X1 port map( A1 => n18155, A2 => n18156, A3 => n18157, A4 => 
                           n18158, ZN => n18145);
   U15417 : NOR4_X1 port map( A1 => n18147, A2 => n18148, A3 => n18149, A4 => 
                           n18150, ZN => n18146);
   U15418 : OAI221_X1 port map( B1 => n14520, B2 => n20737, C1 => n15916, C2 =>
                           n20731, A => n18162, ZN => n18155);
   U15419 : NAND2_X1 port map( A1 => n18127, A2 => n18128, ZN => n5266);
   U15420 : NOR4_X1 port map( A1 => n18137, A2 => n18138, A3 => n18139, A4 => 
                           n18140, ZN => n18127);
   U15421 : NOR4_X1 port map( A1 => n18129, A2 => n18130, A3 => n18131, A4 => 
                           n18132, ZN => n18128);
   U15422 : OAI221_X1 port map( B1 => n14519, B2 => n20737, C1 => n15915, C2 =>
                           n20731, A => n18144, ZN => n18137);
   U15423 : NAND2_X1 port map( A1 => n18109, A2 => n18110, ZN => n5267);
   U15424 : NOR4_X1 port map( A1 => n18119, A2 => n18120, A3 => n18121, A4 => 
                           n18122, ZN => n18109);
   U15425 : NOR4_X1 port map( A1 => n18111, A2 => n18112, A3 => n18113, A4 => 
                           n18114, ZN => n18110);
   U15426 : OAI221_X1 port map( B1 => n14518, B2 => n20737, C1 => n15914, C2 =>
                           n20731, A => n18126, ZN => n18119);
   U15427 : NAND2_X1 port map( A1 => n18091, A2 => n18092, ZN => n5268);
   U15428 : NOR4_X1 port map( A1 => n18101, A2 => n18102, A3 => n18103, A4 => 
                           n18104, ZN => n18091);
   U15429 : NOR4_X1 port map( A1 => n18093, A2 => n18094, A3 => n18095, A4 => 
                           n18096, ZN => n18092);
   U15430 : OAI221_X1 port map( B1 => n14517, B2 => n20737, C1 => n15913, C2 =>
                           n20731, A => n18108, ZN => n18101);
   U15431 : NAND2_X1 port map( A1 => n18073, A2 => n18074, ZN => n5269);
   U15432 : NOR4_X1 port map( A1 => n18083, A2 => n18084, A3 => n18085, A4 => 
                           n18086, ZN => n18073);
   U15433 : NOR4_X1 port map( A1 => n18075, A2 => n18076, A3 => n18077, A4 => 
                           n18078, ZN => n18074);
   U15434 : OAI221_X1 port map( B1 => n14516, B2 => n20738, C1 => n15912, C2 =>
                           n20732, A => n18090, ZN => n18083);
   U15435 : NAND2_X1 port map( A1 => n18055, A2 => n18056, ZN => n5270);
   U15436 : NOR4_X1 port map( A1 => n18065, A2 => n18066, A3 => n18067, A4 => 
                           n18068, ZN => n18055);
   U15437 : NOR4_X1 port map( A1 => n18057, A2 => n18058, A3 => n18059, A4 => 
                           n18060, ZN => n18056);
   U15438 : OAI221_X1 port map( B1 => n14515, B2 => n20738, C1 => n15911, C2 =>
                           n20732, A => n18072, ZN => n18065);
   U15439 : NAND2_X1 port map( A1 => n18037, A2 => n18038, ZN => n5271);
   U15440 : NOR4_X1 port map( A1 => n18047, A2 => n18048, A3 => n18049, A4 => 
                           n18050, ZN => n18037);
   U15441 : NOR4_X1 port map( A1 => n18039, A2 => n18040, A3 => n18041, A4 => 
                           n18042, ZN => n18038);
   U15442 : OAI221_X1 port map( B1 => n14514, B2 => n20738, C1 => n15910, C2 =>
                           n20732, A => n18054, ZN => n18047);
   U15443 : NAND2_X1 port map( A1 => n18019, A2 => n18020, ZN => n5272);
   U15444 : NOR4_X1 port map( A1 => n18029, A2 => n18030, A3 => n18031, A4 => 
                           n18032, ZN => n18019);
   U15445 : NOR4_X1 port map( A1 => n18021, A2 => n18022, A3 => n18023, A4 => 
                           n18024, ZN => n18020);
   U15446 : OAI221_X1 port map( B1 => n14513, B2 => n20738, C1 => n15909, C2 =>
                           n20732, A => n18036, ZN => n18029);
   U15447 : NAND2_X1 port map( A1 => n18001, A2 => n18002, ZN => n5273);
   U15448 : NOR4_X1 port map( A1 => n18011, A2 => n18012, A3 => n18013, A4 => 
                           n18014, ZN => n18001);
   U15449 : NOR4_X1 port map( A1 => n18003, A2 => n18004, A3 => n18005, A4 => 
                           n18006, ZN => n18002);
   U15450 : OAI221_X1 port map( B1 => n14512, B2 => n20738, C1 => n15908, C2 =>
                           n20732, A => n18018, ZN => n18011);
   U15451 : NAND2_X1 port map( A1 => n17983, A2 => n17984, ZN => n5274);
   U15452 : NOR4_X1 port map( A1 => n17993, A2 => n17994, A3 => n17995, A4 => 
                           n17996, ZN => n17983);
   U15453 : NOR4_X1 port map( A1 => n17985, A2 => n17986, A3 => n17987, A4 => 
                           n17988, ZN => n17984);
   U15454 : OAI221_X1 port map( B1 => n14511, B2 => n20738, C1 => n15907, C2 =>
                           n20732, A => n18000, ZN => n17993);
   U15455 : NAND2_X1 port map( A1 => n17965, A2 => n17966, ZN => n5275);
   U15456 : NOR4_X1 port map( A1 => n17975, A2 => n17976, A3 => n17977, A4 => 
                           n17978, ZN => n17965);
   U15457 : NOR4_X1 port map( A1 => n17967, A2 => n17968, A3 => n17969, A4 => 
                           n17970, ZN => n17966);
   U15458 : OAI221_X1 port map( B1 => n14510, B2 => n20738, C1 => n15906, C2 =>
                           n20732, A => n17982, ZN => n17975);
   U15459 : NAND2_X1 port map( A1 => n17947, A2 => n17948, ZN => n5276);
   U15460 : NOR4_X1 port map( A1 => n17957, A2 => n17958, A3 => n17959, A4 => 
                           n17960, ZN => n17947);
   U15461 : NOR4_X1 port map( A1 => n17949, A2 => n17950, A3 => n17951, A4 => 
                           n17952, ZN => n17948);
   U15462 : OAI221_X1 port map( B1 => n14509, B2 => n20738, C1 => n15905, C2 =>
                           n20732, A => n17964, ZN => n17957);
   U15463 : NAND2_X1 port map( A1 => n17929, A2 => n17930, ZN => n5277);
   U15464 : NOR4_X1 port map( A1 => n17939, A2 => n17940, A3 => n17941, A4 => 
                           n17942, ZN => n17929);
   U15465 : NOR4_X1 port map( A1 => n17931, A2 => n17932, A3 => n17933, A4 => 
                           n17934, ZN => n17930);
   U15466 : OAI221_X1 port map( B1 => n14508, B2 => n20738, C1 => n15904, C2 =>
                           n20732, A => n17946, ZN => n17939);
   U15467 : NAND2_X1 port map( A1 => n17911, A2 => n17912, ZN => n5278);
   U15468 : NOR4_X1 port map( A1 => n17921, A2 => n17922, A3 => n17923, A4 => 
                           n17924, ZN => n17911);
   U15469 : NOR4_X1 port map( A1 => n17913, A2 => n17914, A3 => n17915, A4 => 
                           n17916, ZN => n17912);
   U15470 : OAI221_X1 port map( B1 => n14507, B2 => n20738, C1 => n15903, C2 =>
                           n20732, A => n17928, ZN => n17921);
   U15471 : NAND2_X1 port map( A1 => n17893, A2 => n17894, ZN => n5279);
   U15472 : NOR4_X1 port map( A1 => n17903, A2 => n17904, A3 => n17905, A4 => 
                           n17906, ZN => n17893);
   U15473 : NOR4_X1 port map( A1 => n17895, A2 => n17896, A3 => n17897, A4 => 
                           n17898, ZN => n17894);
   U15474 : OAI221_X1 port map( B1 => n14506, B2 => n20738, C1 => n15902, C2 =>
                           n20732, A => n17910, ZN => n17903);
   U15475 : NAND2_X1 port map( A1 => n17875, A2 => n17876, ZN => n5280);
   U15476 : NOR4_X1 port map( A1 => n17885, A2 => n17886, A3 => n17887, A4 => 
                           n17888, ZN => n17875);
   U15477 : NOR4_X1 port map( A1 => n17877, A2 => n17878, A3 => n17879, A4 => 
                           n17880, ZN => n17876);
   U15478 : OAI221_X1 port map( B1 => n14505, B2 => n20738, C1 => n15901, C2 =>
                           n20732, A => n17892, ZN => n17885);
   U15479 : NAND2_X1 port map( A1 => n17857, A2 => n17858, ZN => n5281);
   U15480 : NOR4_X1 port map( A1 => n17867, A2 => n17868, A3 => n17869, A4 => 
                           n17870, ZN => n17857);
   U15481 : NOR4_X1 port map( A1 => n17859, A2 => n17860, A3 => n17861, A4 => 
                           n17862, ZN => n17858);
   U15482 : OAI221_X1 port map( B1 => n14504, B2 => n20739, C1 => n15900, C2 =>
                           n20733, A => n17874, ZN => n17867);
   U15483 : NAND2_X1 port map( A1 => n17839, A2 => n17840, ZN => n5282);
   U15484 : NOR4_X1 port map( A1 => n17849, A2 => n17850, A3 => n17851, A4 => 
                           n17852, ZN => n17839);
   U15485 : NOR4_X1 port map( A1 => n17841, A2 => n17842, A3 => n17843, A4 => 
                           n17844, ZN => n17840);
   U15486 : OAI221_X1 port map( B1 => n14503, B2 => n20739, C1 => n15899, C2 =>
                           n20733, A => n17856, ZN => n17849);
   U15487 : NAND2_X1 port map( A1 => n17821, A2 => n17822, ZN => n5283);
   U15488 : NOR4_X1 port map( A1 => n17831, A2 => n17832, A3 => n17833, A4 => 
                           n17834, ZN => n17821);
   U15489 : NOR4_X1 port map( A1 => n17823, A2 => n17824, A3 => n17825, A4 => 
                           n17826, ZN => n17822);
   U15490 : OAI221_X1 port map( B1 => n14502, B2 => n20739, C1 => n15898, C2 =>
                           n20733, A => n17838, ZN => n17831);
   U15491 : NAND2_X1 port map( A1 => n17803, A2 => n17804, ZN => n5284);
   U15492 : NOR4_X1 port map( A1 => n17813, A2 => n17814, A3 => n17815, A4 => 
                           n17816, ZN => n17803);
   U15493 : NOR4_X1 port map( A1 => n17805, A2 => n17806, A3 => n17807, A4 => 
                           n17808, ZN => n17804);
   U15494 : OAI221_X1 port map( B1 => n14501, B2 => n20739, C1 => n15897, C2 =>
                           n20733, A => n17820, ZN => n17813);
   U15495 : NAND2_X1 port map( A1 => n17785, A2 => n17786, ZN => n5285);
   U15496 : NOR4_X1 port map( A1 => n17795, A2 => n17796, A3 => n17797, A4 => 
                           n17798, ZN => n17785);
   U15497 : NOR4_X1 port map( A1 => n17787, A2 => n17788, A3 => n17789, A4 => 
                           n17790, ZN => n17786);
   U15498 : OAI221_X1 port map( B1 => n14500, B2 => n20739, C1 => n15896, C2 =>
                           n20733, A => n17802, ZN => n17795);
   U15499 : NAND2_X1 port map( A1 => n17767, A2 => n17768, ZN => n5286);
   U15500 : NOR4_X1 port map( A1 => n17777, A2 => n17778, A3 => n17779, A4 => 
                           n17780, ZN => n17767);
   U15501 : NOR4_X1 port map( A1 => n17769, A2 => n17770, A3 => n17771, A4 => 
                           n17772, ZN => n17768);
   U15502 : OAI221_X1 port map( B1 => n14499, B2 => n20739, C1 => n15895, C2 =>
                           n20733, A => n17784, ZN => n17777);
   U15503 : NAND2_X1 port map( A1 => n17749, A2 => n17750, ZN => n5287);
   U15504 : NOR4_X1 port map( A1 => n17759, A2 => n17760, A3 => n17761, A4 => 
                           n17762, ZN => n17749);
   U15505 : NOR4_X1 port map( A1 => n17751, A2 => n17752, A3 => n17753, A4 => 
                           n17754, ZN => n17750);
   U15506 : OAI221_X1 port map( B1 => n14498, B2 => n20739, C1 => n15894, C2 =>
                           n20733, A => n17766, ZN => n17759);
   U15507 : NAND2_X1 port map( A1 => n17731, A2 => n17732, ZN => n5288);
   U15508 : NOR4_X1 port map( A1 => n17741, A2 => n17742, A3 => n17743, A4 => 
                           n17744, ZN => n17731);
   U15509 : NOR4_X1 port map( A1 => n17733, A2 => n17734, A3 => n17735, A4 => 
                           n17736, ZN => n17732);
   U15510 : OAI221_X1 port map( B1 => n14497, B2 => n20739, C1 => n15893, C2 =>
                           n20733, A => n17748, ZN => n17741);
   U15511 : NAND2_X1 port map( A1 => n17713, A2 => n17714, ZN => n5289);
   U15512 : NOR4_X1 port map( A1 => n17723, A2 => n17724, A3 => n17725, A4 => 
                           n17726, ZN => n17713);
   U15513 : NOR4_X1 port map( A1 => n17715, A2 => n17716, A3 => n17717, A4 => 
                           n17718, ZN => n17714);
   U15514 : OAI221_X1 port map( B1 => n14496, B2 => n20739, C1 => n15892, C2 =>
                           n20733, A => n17730, ZN => n17723);
   U15515 : NAND2_X1 port map( A1 => n17695, A2 => n17696, ZN => n5290);
   U15516 : NOR4_X1 port map( A1 => n17705, A2 => n17706, A3 => n17707, A4 => 
                           n17708, ZN => n17695);
   U15517 : NOR4_X1 port map( A1 => n17697, A2 => n17698, A3 => n17699, A4 => 
                           n17700, ZN => n17696);
   U15518 : OAI221_X1 port map( B1 => n14495, B2 => n20739, C1 => n15891, C2 =>
                           n20733, A => n17712, ZN => n17705);
   U15519 : NAND2_X1 port map( A1 => n17677, A2 => n17678, ZN => n5291);
   U15520 : NOR4_X1 port map( A1 => n17687, A2 => n17688, A3 => n17689, A4 => 
                           n17690, ZN => n17677);
   U15521 : NOR4_X1 port map( A1 => n17679, A2 => n17680, A3 => n17681, A4 => 
                           n17682, ZN => n17678);
   U15522 : OAI221_X1 port map( B1 => n14494, B2 => n20739, C1 => n15890, C2 =>
                           n20733, A => n17694, ZN => n17687);
   U15523 : NAND2_X1 port map( A1 => n17659, A2 => n17660, ZN => n5292);
   U15524 : NOR4_X1 port map( A1 => n17669, A2 => n17670, A3 => n17671, A4 => 
                           n17672, ZN => n17659);
   U15525 : NOR4_X1 port map( A1 => n17661, A2 => n17662, A3 => n17663, A4 => 
                           n17664, ZN => n17660);
   U15526 : OAI221_X1 port map( B1 => n14493, B2 => n20739, C1 => n15889, C2 =>
                           n20733, A => n17676, ZN => n17669);
   U15527 : NAND2_X1 port map( A1 => n17641, A2 => n17642, ZN => n5293);
   U15528 : NOR4_X1 port map( A1 => n17651, A2 => n17652, A3 => n17653, A4 => 
                           n17654, ZN => n17641);
   U15529 : NOR4_X1 port map( A1 => n17643, A2 => n17644, A3 => n17645, A4 => 
                           n17646, ZN => n17642);
   U15530 : OAI221_X1 port map( B1 => n14492, B2 => n20740, C1 => n15888, C2 =>
                           n20734, A => n17658, ZN => n17651);
   U15531 : NAND2_X1 port map( A1 => n17623, A2 => n17624, ZN => n5294);
   U15532 : NOR4_X1 port map( A1 => n17633, A2 => n17634, A3 => n17635, A4 => 
                           n17636, ZN => n17623);
   U15533 : NOR4_X1 port map( A1 => n17625, A2 => n17626, A3 => n17627, A4 => 
                           n17628, ZN => n17624);
   U15534 : OAI221_X1 port map( B1 => n14491, B2 => n20740, C1 => n15887, C2 =>
                           n20734, A => n17640, ZN => n17633);
   U15535 : NAND2_X1 port map( A1 => n17605, A2 => n17606, ZN => n5295);
   U15536 : NOR4_X1 port map( A1 => n17615, A2 => n17616, A3 => n17617, A4 => 
                           n17618, ZN => n17605);
   U15537 : NOR4_X1 port map( A1 => n17607, A2 => n17608, A3 => n17609, A4 => 
                           n17610, ZN => n17606);
   U15538 : OAI221_X1 port map( B1 => n14490, B2 => n20740, C1 => n15886, C2 =>
                           n20734, A => n17622, ZN => n17615);
   U15539 : NAND2_X1 port map( A1 => n17587, A2 => n17588, ZN => n5296);
   U15540 : NOR4_X1 port map( A1 => n17597, A2 => n17598, A3 => n17599, A4 => 
                           n17600, ZN => n17587);
   U15541 : NOR4_X1 port map( A1 => n17589, A2 => n17590, A3 => n17591, A4 => 
                           n17592, ZN => n17588);
   U15542 : OAI221_X1 port map( B1 => n14489, B2 => n20740, C1 => n15885, C2 =>
                           n20734, A => n17604, ZN => n17597);
   U15543 : NAND2_X1 port map( A1 => n17569, A2 => n17570, ZN => n5297);
   U15544 : NOR4_X1 port map( A1 => n17579, A2 => n17580, A3 => n17581, A4 => 
                           n17582, ZN => n17569);
   U15545 : NOR4_X1 port map( A1 => n17571, A2 => n17572, A3 => n17573, A4 => 
                           n17574, ZN => n17570);
   U15546 : OAI221_X1 port map( B1 => n14488, B2 => n20740, C1 => n15884, C2 =>
                           n20734, A => n17586, ZN => n17579);
   U15547 : NAND2_X1 port map( A1 => n17551, A2 => n17552, ZN => n5298);
   U15548 : NOR4_X1 port map( A1 => n17561, A2 => n17562, A3 => n17563, A4 => 
                           n17564, ZN => n17551);
   U15549 : NOR4_X1 port map( A1 => n17553, A2 => n17554, A3 => n17555, A4 => 
                           n17556, ZN => n17552);
   U15550 : OAI221_X1 port map( B1 => n14487, B2 => n20740, C1 => n15883, C2 =>
                           n20734, A => n17568, ZN => n17561);
   U15551 : NAND2_X1 port map( A1 => n17533, A2 => n17534, ZN => n5299);
   U15552 : NOR4_X1 port map( A1 => n17543, A2 => n17544, A3 => n17545, A4 => 
                           n17546, ZN => n17533);
   U15553 : NOR4_X1 port map( A1 => n17535, A2 => n17536, A3 => n17537, A4 => 
                           n17538, ZN => n17534);
   U15554 : OAI221_X1 port map( B1 => n14486, B2 => n20740, C1 => n15882, C2 =>
                           n20734, A => n17550, ZN => n17543);
   U15555 : NAND2_X1 port map( A1 => n17515, A2 => n17516, ZN => n5300);
   U15556 : NOR4_X1 port map( A1 => n17525, A2 => n17526, A3 => n17527, A4 => 
                           n17528, ZN => n17515);
   U15557 : NOR4_X1 port map( A1 => n17517, A2 => n17518, A3 => n17519, A4 => 
                           n17520, ZN => n17516);
   U15558 : OAI221_X1 port map( B1 => n14485, B2 => n20740, C1 => n15881, C2 =>
                           n20734, A => n17532, ZN => n17525);
   U15559 : NAND2_X1 port map( A1 => n17497, A2 => n17498, ZN => n5301);
   U15560 : NOR4_X1 port map( A1 => n17507, A2 => n17508, A3 => n17509, A4 => 
                           n17510, ZN => n17497);
   U15561 : NOR4_X1 port map( A1 => n17499, A2 => n17500, A3 => n17501, A4 => 
                           n17502, ZN => n17498);
   U15562 : OAI221_X1 port map( B1 => n14484, B2 => n20740, C1 => n15880, C2 =>
                           n20734, A => n17514, ZN => n17507);
   U15563 : NAND2_X1 port map( A1 => n17479, A2 => n17480, ZN => n5302);
   U15564 : NOR4_X1 port map( A1 => n17489, A2 => n17490, A3 => n17491, A4 => 
                           n17492, ZN => n17479);
   U15565 : NOR4_X1 port map( A1 => n17481, A2 => n17482, A3 => n17483, A4 => 
                           n17484, ZN => n17480);
   U15566 : OAI221_X1 port map( B1 => n14483, B2 => n20740, C1 => n15879, C2 =>
                           n20734, A => n17496, ZN => n17489);
   U15567 : NAND2_X1 port map( A1 => n17461, A2 => n17462, ZN => n5303);
   U15568 : NOR4_X1 port map( A1 => n17471, A2 => n17472, A3 => n17473, A4 => 
                           n17474, ZN => n17461);
   U15569 : NOR4_X1 port map( A1 => n17463, A2 => n17464, A3 => n17465, A4 => 
                           n17466, ZN => n17462);
   U15570 : OAI221_X1 port map( B1 => n14482, B2 => n20740, C1 => n15878, C2 =>
                           n20734, A => n17478, ZN => n17471);
   U15571 : NAND2_X1 port map( A1 => n17443, A2 => n17444, ZN => n5304);
   U15572 : NOR4_X1 port map( A1 => n17453, A2 => n17454, A3 => n17455, A4 => 
                           n17456, ZN => n17443);
   U15573 : NOR4_X1 port map( A1 => n17445, A2 => n17446, A3 => n17447, A4 => 
                           n17448, ZN => n17444);
   U15574 : OAI221_X1 port map( B1 => n14481, B2 => n20740, C1 => n15877, C2 =>
                           n20734, A => n17460, ZN => n17453);
   U15575 : NAND2_X1 port map( A1 => n17304, A2 => n17305, ZN => n5309);
   U15576 : NOR4_X1 port map( A1 => n17325, A2 => n17326, A3 => n17327, A4 => 
                           n17328, ZN => n17304);
   U15577 : NOR4_X1 port map( A1 => n17306, A2 => n17307, A3 => n17308, A4 => 
                           n17309, ZN => n17305);
   U15578 : OAI221_X1 port map( B1 => n14540, B2 => n20928, C1 => n15936, C2 =>
                           n20922, A => n17336, ZN => n17325);
   U15579 : NAND2_X1 port map( A1 => n17284, A2 => n17285, ZN => n5311);
   U15580 : NOR4_X1 port map( A1 => n17294, A2 => n17295, A3 => n17296, A4 => 
                           n17297, ZN => n17284);
   U15581 : NOR4_X1 port map( A1 => n17286, A2 => n17287, A3 => n17288, A4 => 
                           n17289, ZN => n17285);
   U15582 : OAI221_X1 port map( B1 => n14539, B2 => n20928, C1 => n15935, C2 =>
                           n20922, A => n17301, ZN => n17294);
   U15583 : NAND2_X1 port map( A1 => n17265, A2 => n17266, ZN => n5313);
   U15584 : NOR4_X1 port map( A1 => n17275, A2 => n17276, A3 => n17277, A4 => 
                           n17278, ZN => n17265);
   U15585 : NOR4_X1 port map( A1 => n17267, A2 => n17268, A3 => n17269, A4 => 
                           n17270, ZN => n17266);
   U15586 : OAI221_X1 port map( B1 => n14538, B2 => n20928, C1 => n15934, C2 =>
                           n20922, A => n17282, ZN => n17275);
   U15587 : NAND2_X1 port map( A1 => n17246, A2 => n17247, ZN => n5315);
   U15588 : NOR4_X1 port map( A1 => n17256, A2 => n17257, A3 => n17258, A4 => 
                           n17259, ZN => n17246);
   U15589 : NOR4_X1 port map( A1 => n17248, A2 => n17249, A3 => n17250, A4 => 
                           n17251, ZN => n17247);
   U15590 : OAI221_X1 port map( B1 => n14537, B2 => n20928, C1 => n15933, C2 =>
                           n20922, A => n17263, ZN => n17256);
   U15591 : NAND2_X1 port map( A1 => n17227, A2 => n17228, ZN => n5317);
   U15592 : NOR4_X1 port map( A1 => n17237, A2 => n17238, A3 => n17239, A4 => 
                           n17240, ZN => n17227);
   U15593 : NOR4_X1 port map( A1 => n17229, A2 => n17230, A3 => n17231, A4 => 
                           n17232, ZN => n17228);
   U15594 : OAI221_X1 port map( B1 => n14536, B2 => n20928, C1 => n15932, C2 =>
                           n20922, A => n17244, ZN => n17237);
   U15595 : NAND2_X1 port map( A1 => n17208, A2 => n17209, ZN => n5319);
   U15596 : NOR4_X1 port map( A1 => n17218, A2 => n17219, A3 => n17220, A4 => 
                           n17221, ZN => n17208);
   U15597 : NOR4_X1 port map( A1 => n17210, A2 => n17211, A3 => n17212, A4 => 
                           n17213, ZN => n17209);
   U15598 : OAI221_X1 port map( B1 => n14535, B2 => n20928, C1 => n15931, C2 =>
                           n20922, A => n17225, ZN => n17218);
   U15599 : NAND2_X1 port map( A1 => n17189, A2 => n17190, ZN => n5321);
   U15600 : NOR4_X1 port map( A1 => n17199, A2 => n17200, A3 => n17201, A4 => 
                           n17202, ZN => n17189);
   U15601 : NOR4_X1 port map( A1 => n17191, A2 => n17192, A3 => n17193, A4 => 
                           n17194, ZN => n17190);
   U15602 : OAI221_X1 port map( B1 => n14534, B2 => n20928, C1 => n15930, C2 =>
                           n20922, A => n17206, ZN => n17199);
   U15603 : NAND2_X1 port map( A1 => n17170, A2 => n17171, ZN => n5323);
   U15604 : NOR4_X1 port map( A1 => n17180, A2 => n17181, A3 => n17182, A4 => 
                           n17183, ZN => n17170);
   U15605 : NOR4_X1 port map( A1 => n17172, A2 => n17173, A3 => n17174, A4 => 
                           n17175, ZN => n17171);
   U15606 : OAI221_X1 port map( B1 => n14533, B2 => n20928, C1 => n15929, C2 =>
                           n20922, A => n17187, ZN => n17180);
   U15607 : NAND2_X1 port map( A1 => n17151, A2 => n17152, ZN => n5325);
   U15608 : NOR4_X1 port map( A1 => n17161, A2 => n17162, A3 => n17163, A4 => 
                           n17164, ZN => n17151);
   U15609 : NOR4_X1 port map( A1 => n17153, A2 => n17154, A3 => n17155, A4 => 
                           n17156, ZN => n17152);
   U15610 : OAI221_X1 port map( B1 => n14532, B2 => n20928, C1 => n15928, C2 =>
                           n20922, A => n17168, ZN => n17161);
   U15611 : NAND2_X1 port map( A1 => n17132, A2 => n17133, ZN => n5327);
   U15612 : NOR4_X1 port map( A1 => n17142, A2 => n17143, A3 => n17144, A4 => 
                           n17145, ZN => n17132);
   U15613 : NOR4_X1 port map( A1 => n17134, A2 => n17135, A3 => n17136, A4 => 
                           n17137, ZN => n17133);
   U15614 : OAI221_X1 port map( B1 => n14531, B2 => n20928, C1 => n15927, C2 =>
                           n20922, A => n17149, ZN => n17142);
   U15615 : NAND2_X1 port map( A1 => n17113, A2 => n17114, ZN => n5329);
   U15616 : NOR4_X1 port map( A1 => n17123, A2 => n17124, A3 => n17125, A4 => 
                           n17126, ZN => n17113);
   U15617 : NOR4_X1 port map( A1 => n17115, A2 => n17116, A3 => n17117, A4 => 
                           n17118, ZN => n17114);
   U15618 : OAI221_X1 port map( B1 => n14530, B2 => n20928, C1 => n15926, C2 =>
                           n20922, A => n17130, ZN => n17123);
   U15619 : NAND2_X1 port map( A1 => n17094, A2 => n17095, ZN => n5331);
   U15620 : NOR4_X1 port map( A1 => n17104, A2 => n17105, A3 => n17106, A4 => 
                           n17107, ZN => n17094);
   U15621 : NOR4_X1 port map( A1 => n17096, A2 => n17097, A3 => n17098, A4 => 
                           n17099, ZN => n17095);
   U15622 : OAI221_X1 port map( B1 => n14529, B2 => n20928, C1 => n15925, C2 =>
                           n20922, A => n17111, ZN => n17104);
   U15623 : NAND2_X1 port map( A1 => n16866, A2 => n16867, ZN => n5355);
   U15624 : NOR4_X1 port map( A1 => n16876, A2 => n16877, A3 => n16878, A4 => 
                           n16879, ZN => n16866);
   U15625 : NOR4_X1 port map( A1 => n16868, A2 => n16869, A3 => n16870, A4 => 
                           n16871, ZN => n16867);
   U15626 : OAI221_X1 port map( B1 => n14517, B2 => n20929, C1 => n15913, C2 =>
                           n20923, A => n16883, ZN => n16876);
   U15627 : NAND2_X1 port map( A1 => n16847, A2 => n16848, ZN => n5357);
   U15628 : NOR4_X1 port map( A1 => n16857, A2 => n16858, A3 => n16859, A4 => 
                           n16860, ZN => n16847);
   U15629 : NOR4_X1 port map( A1 => n16849, A2 => n16850, A3 => n16851, A4 => 
                           n16852, ZN => n16848);
   U15630 : OAI221_X1 port map( B1 => n14516, B2 => n20930, C1 => n15912, C2 =>
                           n20924, A => n16864, ZN => n16857);
   U15631 : NAND2_X1 port map( A1 => n16828, A2 => n16829, ZN => n5359);
   U15632 : NOR4_X1 port map( A1 => n16838, A2 => n16839, A3 => n16840, A4 => 
                           n16841, ZN => n16828);
   U15633 : NOR4_X1 port map( A1 => n16830, A2 => n16831, A3 => n16832, A4 => 
                           n16833, ZN => n16829);
   U15634 : OAI221_X1 port map( B1 => n14515, B2 => n20930, C1 => n15911, C2 =>
                           n20924, A => n16845, ZN => n16838);
   U15635 : NAND2_X1 port map( A1 => n16809, A2 => n16810, ZN => n5361);
   U15636 : NOR4_X1 port map( A1 => n16819, A2 => n16820, A3 => n16821, A4 => 
                           n16822, ZN => n16809);
   U15637 : NOR4_X1 port map( A1 => n16811, A2 => n16812, A3 => n16813, A4 => 
                           n16814, ZN => n16810);
   U15638 : OAI221_X1 port map( B1 => n14514, B2 => n20930, C1 => n15910, C2 =>
                           n20924, A => n16826, ZN => n16819);
   U15639 : NAND2_X1 port map( A1 => n16790, A2 => n16791, ZN => n5363);
   U15640 : NOR4_X1 port map( A1 => n16800, A2 => n16801, A3 => n16802, A4 => 
                           n16803, ZN => n16790);
   U15641 : NOR4_X1 port map( A1 => n16792, A2 => n16793, A3 => n16794, A4 => 
                           n16795, ZN => n16791);
   U15642 : OAI221_X1 port map( B1 => n14513, B2 => n20930, C1 => n15909, C2 =>
                           n20924, A => n16807, ZN => n16800);
   U15643 : NAND2_X1 port map( A1 => n16771, A2 => n16772, ZN => n5365);
   U15644 : NOR4_X1 port map( A1 => n16781, A2 => n16782, A3 => n16783, A4 => 
                           n16784, ZN => n16771);
   U15645 : NOR4_X1 port map( A1 => n16773, A2 => n16774, A3 => n16775, A4 => 
                           n16776, ZN => n16772);
   U15646 : OAI221_X1 port map( B1 => n14512, B2 => n20930, C1 => n15908, C2 =>
                           n20924, A => n16788, ZN => n16781);
   U15647 : NAND2_X1 port map( A1 => n16752, A2 => n16753, ZN => n5367);
   U15648 : NOR4_X1 port map( A1 => n16762, A2 => n16763, A3 => n16764, A4 => 
                           n16765, ZN => n16752);
   U15649 : NOR4_X1 port map( A1 => n16754, A2 => n16755, A3 => n16756, A4 => 
                           n16757, ZN => n16753);
   U15650 : OAI221_X1 port map( B1 => n14511, B2 => n20930, C1 => n15907, C2 =>
                           n20924, A => n16769, ZN => n16762);
   U15651 : NAND2_X1 port map( A1 => n16733, A2 => n16734, ZN => n5369);
   U15652 : NOR4_X1 port map( A1 => n16743, A2 => n16744, A3 => n16745, A4 => 
                           n16746, ZN => n16733);
   U15653 : NOR4_X1 port map( A1 => n16735, A2 => n16736, A3 => n16737, A4 => 
                           n16738, ZN => n16734);
   U15654 : OAI221_X1 port map( B1 => n14510, B2 => n20930, C1 => n15906, C2 =>
                           n20924, A => n16750, ZN => n16743);
   U15655 : NAND2_X1 port map( A1 => n16714, A2 => n16715, ZN => n5371);
   U15656 : NOR4_X1 port map( A1 => n16724, A2 => n16725, A3 => n16726, A4 => 
                           n16727, ZN => n16714);
   U15657 : NOR4_X1 port map( A1 => n16716, A2 => n16717, A3 => n16718, A4 => 
                           n16719, ZN => n16715);
   U15658 : OAI221_X1 port map( B1 => n14509, B2 => n20930, C1 => n15905, C2 =>
                           n20924, A => n16731, ZN => n16724);
   U15659 : NAND2_X1 port map( A1 => n16695, A2 => n16696, ZN => n5373);
   U15660 : NOR4_X1 port map( A1 => n16705, A2 => n16706, A3 => n16707, A4 => 
                           n16708, ZN => n16695);
   U15661 : NOR4_X1 port map( A1 => n16697, A2 => n16698, A3 => n16699, A4 => 
                           n16700, ZN => n16696);
   U15662 : OAI221_X1 port map( B1 => n14508, B2 => n20930, C1 => n15904, C2 =>
                           n20924, A => n16712, ZN => n16705);
   U15663 : NAND2_X1 port map( A1 => n16676, A2 => n16677, ZN => n5375);
   U15664 : NOR4_X1 port map( A1 => n16686, A2 => n16687, A3 => n16688, A4 => 
                           n16689, ZN => n16676);
   U15665 : NOR4_X1 port map( A1 => n16678, A2 => n16679, A3 => n16680, A4 => 
                           n16681, ZN => n16677);
   U15666 : OAI221_X1 port map( B1 => n14507, B2 => n20930, C1 => n15903, C2 =>
                           n20924, A => n16693, ZN => n16686);
   U15667 : NAND2_X1 port map( A1 => n16657, A2 => n16658, ZN => n5377);
   U15668 : NOR4_X1 port map( A1 => n16667, A2 => n16668, A3 => n16669, A4 => 
                           n16670, ZN => n16657);
   U15669 : NOR4_X1 port map( A1 => n16659, A2 => n16660, A3 => n16661, A4 => 
                           n16662, ZN => n16658);
   U15670 : OAI221_X1 port map( B1 => n14506, B2 => n20930, C1 => n15902, C2 =>
                           n20924, A => n16674, ZN => n16667);
   U15671 : NAND2_X1 port map( A1 => n16638, A2 => n16639, ZN => n5379);
   U15672 : NOR4_X1 port map( A1 => n16648, A2 => n16649, A3 => n16650, A4 => 
                           n16651, ZN => n16638);
   U15673 : NOR4_X1 port map( A1 => n16640, A2 => n16641, A3 => n16642, A4 => 
                           n16643, ZN => n16639);
   U15674 : OAI221_X1 port map( B1 => n14505, B2 => n20930, C1 => n15901, C2 =>
                           n20924, A => n16655, ZN => n16648);
   U15675 : NAND2_X1 port map( A1 => n16619, A2 => n16620, ZN => n5381);
   U15676 : NOR4_X1 port map( A1 => n16629, A2 => n16630, A3 => n16631, A4 => 
                           n16632, ZN => n16619);
   U15677 : NOR4_X1 port map( A1 => n16621, A2 => n16622, A3 => n16623, A4 => 
                           n16624, ZN => n16620);
   U15678 : OAI221_X1 port map( B1 => n14504, B2 => n20931, C1 => n15900, C2 =>
                           n20925, A => n16636, ZN => n16629);
   U15679 : NAND2_X1 port map( A1 => n16600, A2 => n16601, ZN => n5383);
   U15680 : NOR4_X1 port map( A1 => n16610, A2 => n16611, A3 => n16612, A4 => 
                           n16613, ZN => n16600);
   U15681 : NOR4_X1 port map( A1 => n16602, A2 => n16603, A3 => n16604, A4 => 
                           n16605, ZN => n16601);
   U15682 : OAI221_X1 port map( B1 => n14503, B2 => n20931, C1 => n15899, C2 =>
                           n20925, A => n16617, ZN => n16610);
   U15683 : NAND2_X1 port map( A1 => n16581, A2 => n16582, ZN => n5385);
   U15684 : NOR4_X1 port map( A1 => n16591, A2 => n16592, A3 => n16593, A4 => 
                           n16594, ZN => n16581);
   U15685 : NOR4_X1 port map( A1 => n16583, A2 => n16584, A3 => n16585, A4 => 
                           n16586, ZN => n16582);
   U15686 : OAI221_X1 port map( B1 => n14502, B2 => n20931, C1 => n15898, C2 =>
                           n20925, A => n16598, ZN => n16591);
   U15687 : NAND2_X1 port map( A1 => n16562, A2 => n16563, ZN => n5387);
   U15688 : NOR4_X1 port map( A1 => n16572, A2 => n16573, A3 => n16574, A4 => 
                           n16575, ZN => n16562);
   U15689 : NOR4_X1 port map( A1 => n16564, A2 => n16565, A3 => n16566, A4 => 
                           n16567, ZN => n16563);
   U15690 : OAI221_X1 port map( B1 => n14501, B2 => n20931, C1 => n15897, C2 =>
                           n20925, A => n16579, ZN => n16572);
   U15691 : NAND2_X1 port map( A1 => n16543, A2 => n16544, ZN => n5389);
   U15692 : NOR4_X1 port map( A1 => n16553, A2 => n16554, A3 => n16555, A4 => 
                           n16556, ZN => n16543);
   U15693 : NOR4_X1 port map( A1 => n16545, A2 => n16546, A3 => n16547, A4 => 
                           n16548, ZN => n16544);
   U15694 : OAI221_X1 port map( B1 => n14500, B2 => n20931, C1 => n15896, C2 =>
                           n20925, A => n16560, ZN => n16553);
   U15695 : NAND2_X1 port map( A1 => n16524, A2 => n16525, ZN => n5391);
   U15696 : NOR4_X1 port map( A1 => n16534, A2 => n16535, A3 => n16536, A4 => 
                           n16537, ZN => n16524);
   U15697 : NOR4_X1 port map( A1 => n16526, A2 => n16527, A3 => n16528, A4 => 
                           n16529, ZN => n16525);
   U15698 : OAI221_X1 port map( B1 => n14499, B2 => n20931, C1 => n15895, C2 =>
                           n20925, A => n16541, ZN => n16534);
   U15699 : NAND2_X1 port map( A1 => n16505, A2 => n16506, ZN => n5393);
   U15700 : NOR4_X1 port map( A1 => n16515, A2 => n16516, A3 => n16517, A4 => 
                           n16518, ZN => n16505);
   U15701 : NOR4_X1 port map( A1 => n16507, A2 => n16508, A3 => n16509, A4 => 
                           n16510, ZN => n16506);
   U15702 : OAI221_X1 port map( B1 => n14498, B2 => n20931, C1 => n15894, C2 =>
                           n20925, A => n16522, ZN => n16515);
   U15703 : NAND2_X1 port map( A1 => n16486, A2 => n16487, ZN => n5395);
   U15704 : NOR4_X1 port map( A1 => n16496, A2 => n16497, A3 => n16498, A4 => 
                           n16499, ZN => n16486);
   U15705 : NOR4_X1 port map( A1 => n16488, A2 => n16489, A3 => n16490, A4 => 
                           n16491, ZN => n16487);
   U15706 : OAI221_X1 port map( B1 => n14497, B2 => n20931, C1 => n15893, C2 =>
                           n20925, A => n16503, ZN => n16496);
   U15707 : NAND2_X1 port map( A1 => n16467, A2 => n16468, ZN => n5397);
   U15708 : NOR4_X1 port map( A1 => n16477, A2 => n16478, A3 => n16479, A4 => 
                           n16480, ZN => n16467);
   U15709 : NOR4_X1 port map( A1 => n16469, A2 => n16470, A3 => n16471, A4 => 
                           n16472, ZN => n16468);
   U15710 : OAI221_X1 port map( B1 => n14496, B2 => n20931, C1 => n15892, C2 =>
                           n20925, A => n16484, ZN => n16477);
   U15711 : NAND2_X1 port map( A1 => n16448, A2 => n16449, ZN => n5399);
   U15712 : NOR4_X1 port map( A1 => n16458, A2 => n16459, A3 => n16460, A4 => 
                           n16461, ZN => n16448);
   U15713 : NOR4_X1 port map( A1 => n16450, A2 => n16451, A3 => n16452, A4 => 
                           n16453, ZN => n16449);
   U15714 : OAI221_X1 port map( B1 => n14495, B2 => n20931, C1 => n15891, C2 =>
                           n20925, A => n16465, ZN => n16458);
   U15715 : NAND2_X1 port map( A1 => n16429, A2 => n16430, ZN => n5401);
   U15716 : NOR4_X1 port map( A1 => n16439, A2 => n16440, A3 => n16441, A4 => 
                           n16442, ZN => n16429);
   U15717 : NOR4_X1 port map( A1 => n16431, A2 => n16432, A3 => n16433, A4 => 
                           n16434, ZN => n16430);
   U15718 : OAI221_X1 port map( B1 => n14494, B2 => n20931, C1 => n15890, C2 =>
                           n20925, A => n16446, ZN => n16439);
   U15719 : NAND2_X1 port map( A1 => n16410, A2 => n16411, ZN => n5403);
   U15720 : NOR4_X1 port map( A1 => n16420, A2 => n16421, A3 => n16422, A4 => 
                           n16423, ZN => n16410);
   U15721 : NOR4_X1 port map( A1 => n16412, A2 => n16413, A3 => n16414, A4 => 
                           n16415, ZN => n16411);
   U15722 : OAI221_X1 port map( B1 => n14493, B2 => n20931, C1 => n15889, C2 =>
                           n20925, A => n16427, ZN => n16420);
   U15723 : NAND2_X1 port map( A1 => n16391, A2 => n16392, ZN => n5405);
   U15724 : NOR4_X1 port map( A1 => n16401, A2 => n16402, A3 => n16403, A4 => 
                           n16404, ZN => n16391);
   U15725 : NOR4_X1 port map( A1 => n16393, A2 => n16394, A3 => n16395, A4 => 
                           n16396, ZN => n16392);
   U15726 : OAI221_X1 port map( B1 => n14492, B2 => n20932, C1 => n15888, C2 =>
                           n20926, A => n16408, ZN => n16401);
   U15727 : NAND2_X1 port map( A1 => n16372, A2 => n16373, ZN => n5407);
   U15728 : NOR4_X1 port map( A1 => n16382, A2 => n16383, A3 => n16384, A4 => 
                           n16385, ZN => n16372);
   U15729 : NOR4_X1 port map( A1 => n16374, A2 => n16375, A3 => n16376, A4 => 
                           n16377, ZN => n16373);
   U15730 : OAI221_X1 port map( B1 => n14491, B2 => n20932, C1 => n15887, C2 =>
                           n20926, A => n16389, ZN => n16382);
   U15731 : NAND2_X1 port map( A1 => n16353, A2 => n16354, ZN => n5409);
   U15732 : NOR4_X1 port map( A1 => n16363, A2 => n16364, A3 => n16365, A4 => 
                           n16366, ZN => n16353);
   U15733 : NOR4_X1 port map( A1 => n16355, A2 => n16356, A3 => n16357, A4 => 
                           n16358, ZN => n16354);
   U15734 : OAI221_X1 port map( B1 => n14490, B2 => n20932, C1 => n15886, C2 =>
                           n20926, A => n16370, ZN => n16363);
   U15735 : NAND2_X1 port map( A1 => n16315, A2 => n16316, ZN => n5413);
   U15736 : NOR4_X1 port map( A1 => n16325, A2 => n16326, A3 => n16327, A4 => 
                           n16328, ZN => n16315);
   U15737 : NOR4_X1 port map( A1 => n16317, A2 => n16318, A3 => n16319, A4 => 
                           n16320, ZN => n16316);
   U15738 : OAI221_X1 port map( B1 => n14488, B2 => n20932, C1 => n15884, C2 =>
                           n20926, A => n16332, ZN => n16325);
   U15739 : NAND2_X1 port map( A1 => n16296, A2 => n16297, ZN => n5415);
   U15740 : NOR4_X1 port map( A1 => n16306, A2 => n16307, A3 => n16308, A4 => 
                           n16309, ZN => n16296);
   U15741 : NOR4_X1 port map( A1 => n16298, A2 => n16299, A3 => n16300, A4 => 
                           n16301, ZN => n16297);
   U15742 : OAI221_X1 port map( B1 => n14487, B2 => n20932, C1 => n15883, C2 =>
                           n20926, A => n16313, ZN => n16306);
   U15743 : NAND2_X1 port map( A1 => n16277, A2 => n16278, ZN => n5417);
   U15744 : NOR4_X1 port map( A1 => n16287, A2 => n16288, A3 => n16289, A4 => 
                           n16290, ZN => n16277);
   U15745 : NOR4_X1 port map( A1 => n16279, A2 => n16280, A3 => n16281, A4 => 
                           n16282, ZN => n16278);
   U15746 : OAI221_X1 port map( B1 => n14486, B2 => n20932, C1 => n15882, C2 =>
                           n20926, A => n16294, ZN => n16287);
   U15747 : NAND2_X1 port map( A1 => n16258, A2 => n16259, ZN => n5419);
   U15748 : NOR4_X1 port map( A1 => n16268, A2 => n16269, A3 => n16270, A4 => 
                           n16271, ZN => n16258);
   U15749 : NOR4_X1 port map( A1 => n16260, A2 => n16261, A3 => n16262, A4 => 
                           n16263, ZN => n16259);
   U15750 : OAI221_X1 port map( B1 => n14485, B2 => n20932, C1 => n15881, C2 =>
                           n20926, A => n16275, ZN => n16268);
   U15751 : NAND2_X1 port map( A1 => n16239, A2 => n16240, ZN => n5421);
   U15752 : NOR4_X1 port map( A1 => n16249, A2 => n16250, A3 => n16251, A4 => 
                           n16252, ZN => n16239);
   U15753 : NOR4_X1 port map( A1 => n16241, A2 => n16242, A3 => n16243, A4 => 
                           n16244, ZN => n16240);
   U15754 : OAI221_X1 port map( B1 => n14484, B2 => n20932, C1 => n15880, C2 =>
                           n20926, A => n16256, ZN => n16249);
   U15755 : NAND2_X1 port map( A1 => n16220, A2 => n16221, ZN => n5423);
   U15756 : NOR4_X1 port map( A1 => n16230, A2 => n16231, A3 => n16232, A4 => 
                           n16233, ZN => n16220);
   U15757 : NOR4_X1 port map( A1 => n16222, A2 => n16223, A3 => n16224, A4 => 
                           n16225, ZN => n16221);
   U15758 : OAI221_X1 port map( B1 => n14483, B2 => n20932, C1 => n15879, C2 =>
                           n20926, A => n16237, ZN => n16230);
   U15759 : NAND2_X1 port map( A1 => n16201, A2 => n16202, ZN => n5425);
   U15760 : NOR4_X1 port map( A1 => n16211, A2 => n16212, A3 => n16213, A4 => 
                           n16214, ZN => n16201);
   U15761 : NOR4_X1 port map( A1 => n16203, A2 => n16204, A3 => n16205, A4 => 
                           n16206, ZN => n16202);
   U15762 : OAI221_X1 port map( B1 => n14482, B2 => n20932, C1 => n15878, C2 =>
                           n20926, A => n16218, ZN => n16211);
   U15763 : NAND2_X1 port map( A1 => n16182, A2 => n16183, ZN => n5427);
   U15764 : NOR4_X1 port map( A1 => n16192, A2 => n16193, A3 => n16194, A4 => 
                           n16195, ZN => n16182);
   U15765 : NOR4_X1 port map( A1 => n16184, A2 => n16185, A3 => n16186, A4 => 
                           n16187, ZN => n16183);
   U15766 : OAI221_X1 port map( B1 => n14481, B2 => n20932, C1 => n15877, C2 =>
                           n20926, A => n16199, ZN => n16192);
   U15767 : AND2_X1 port map( A1 => n17318, A2 => n17313, ZN => n16085);
   U15768 : BUF_X1 port map( A => n14069, Z => n21520);
   U15769 : NOR3_X1 port map( A1 => n18534, A2 => ADD_RD2(0), A3 => n18532, ZN 
                           => n18523);
   U15770 : NOR3_X1 port map( A1 => n17333, A2 => ADD_RD1(0), A3 => n17331, ZN 
                           => n17322);
   U15771 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n18535,
                           ZN => n18517);
   U15772 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n17334,
                           ZN => n17316);
   U15773 : NOR3_X1 port map( A1 => n17334, A2 => ADD_RD1(4), A3 => n17333, ZN 
                           => n17319);
   U15774 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n17333,
                           ZN => n17315);
   U15775 : NOR3_X1 port map( A1 => n18535, A2 => ADD_RD2(3), A3 => n18532, ZN 
                           => n18524);
   U15776 : NOR3_X1 port map( A1 => n17334, A2 => ADD_RD1(3), A3 => n17331, ZN 
                           => n17323);
   U15777 : NOR3_X1 port map( A1 => n18535, A2 => ADD_RD2(4), A3 => n18534, ZN 
                           => n18519);
   U15778 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n18534,
                           ZN => n18516);
   U15779 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n18521);
   U15780 : OAI221_X1 port map( B1 => n14137, B2 => n21037, C1 => n15668, C2 =>
                           n21031, A => n17324, ZN => n17306);
   U15781 : AOI222_X1 port map( A1 => n21025, A2 => n19801, B1 => n21019, B2 =>
                           n9209, C1 => n21013, C2 => n8825, ZN => n17324);
   U15782 : OAI221_X1 port map( B1 => n14136, B2 => n21037, C1 => n15667, C2 =>
                           n21031, A => n17293, ZN => n17286);
   U15783 : AOI222_X1 port map( A1 => n21025, A2 => n19781, B1 => n21019, B2 =>
                           n9205, C1 => n21013, C2 => n8821, ZN => n17293);
   U15784 : OAI221_X1 port map( B1 => n14135, B2 => n21037, C1 => n15666, C2 =>
                           n21031, A => n17274, ZN => n17267);
   U15785 : AOI222_X1 port map( A1 => n21025, A2 => n19761, B1 => n21019, B2 =>
                           n9201, C1 => n21013, C2 => n8817, ZN => n17274);
   U15786 : OAI221_X1 port map( B1 => n14134, B2 => n21037, C1 => n15665, C2 =>
                           n21031, A => n17255, ZN => n17248);
   U15787 : AOI222_X1 port map( A1 => n21025, A2 => n19741, B1 => n21019, B2 =>
                           n9197, C1 => n21013, C2 => n8813, ZN => n17255);
   U15788 : OAI221_X1 port map( B1 => n14133, B2 => n21037, C1 => n15664, C2 =>
                           n21031, A => n17236, ZN => n17229);
   U15789 : AOI222_X1 port map( A1 => n21025, A2 => n19721, B1 => n21019, B2 =>
                           n9193, C1 => n21013, C2 => n8809, ZN => n17236);
   U15790 : OAI221_X1 port map( B1 => n14132, B2 => n21037, C1 => n15663, C2 =>
                           n21031, A => n17217, ZN => n17210);
   U15791 : AOI222_X1 port map( A1 => n21025, A2 => n19701, B1 => n21019, B2 =>
                           n9189, C1 => n21013, C2 => n8805, ZN => n17217);
   U15792 : OAI221_X1 port map( B1 => n14131, B2 => n21037, C1 => n15662, C2 =>
                           n21031, A => n17198, ZN => n17191);
   U15793 : AOI222_X1 port map( A1 => n21025, A2 => n19681, B1 => n21019, B2 =>
                           n9185, C1 => n21013, C2 => n8801, ZN => n17198);
   U15794 : OAI221_X1 port map( B1 => n14130, B2 => n21037, C1 => n15661, C2 =>
                           n21031, A => n17179, ZN => n17172);
   U15795 : AOI222_X1 port map( A1 => n21025, A2 => n19661, B1 => n21019, B2 =>
                           n9181, C1 => n21013, C2 => n8797, ZN => n17179);
   U15796 : OAI221_X1 port map( B1 => n14129, B2 => n21037, C1 => n15660, C2 =>
                           n21031, A => n17160, ZN => n17153);
   U15797 : AOI222_X1 port map( A1 => n21025, A2 => n19641, B1 => n21019, B2 =>
                           n9177, C1 => n21013, C2 => n8793, ZN => n17160);
   U15798 : OAI221_X1 port map( B1 => n14128, B2 => n21037, C1 => n15659, C2 =>
                           n21031, A => n17141, ZN => n17134);
   U15799 : AOI222_X1 port map( A1 => n21025, A2 => n19621, B1 => n21019, B2 =>
                           n9173, C1 => n21013, C2 => n8789, ZN => n17141);
   U15800 : OAI221_X1 port map( B1 => n14127, B2 => n21037, C1 => n15658, C2 =>
                           n21031, A => n17122, ZN => n17115);
   U15801 : AOI222_X1 port map( A1 => n21025, A2 => n19601, B1 => n21019, B2 =>
                           n9169, C1 => n21013, C2 => n8785, ZN => n17122);
   U15802 : OAI221_X1 port map( B1 => n14126, B2 => n21037, C1 => n15657, C2 =>
                           n21031, A => n17103, ZN => n17096);
   U15803 : AOI222_X1 port map( A1 => n21025, A2 => n19581, B1 => n21019, B2 =>
                           n9165, C1 => n21013, C2 => n8781, ZN => n17103);
   U15804 : OAI221_X1 port map( B1 => n14125, B2 => n21038, C1 => n15656, C2 =>
                           n21032, A => n17084, ZN => n17077);
   U15805 : AOI222_X1 port map( A1 => n21026, A2 => n19561, B1 => n21020, B2 =>
                           n9161, C1 => n21014, C2 => n8777, ZN => n17084);
   U15806 : OAI221_X1 port map( B1 => n14124, B2 => n21038, C1 => n15655, C2 =>
                           n21032, A => n17065, ZN => n17058);
   U15807 : AOI222_X1 port map( A1 => n21026, A2 => n19541, B1 => n21020, B2 =>
                           n9157, C1 => n21014, C2 => n8773, ZN => n17065);
   U15808 : OAI221_X1 port map( B1 => n14123, B2 => n21038, C1 => n15654, C2 =>
                           n21032, A => n17046, ZN => n17039);
   U15809 : AOI222_X1 port map( A1 => n21026, A2 => n19521, B1 => n21020, B2 =>
                           n9153, C1 => n21014, C2 => n8769, ZN => n17046);
   U15810 : OAI221_X1 port map( B1 => n14122, B2 => n21038, C1 => n15653, C2 =>
                           n21032, A => n17027, ZN => n17020);
   U15811 : AOI222_X1 port map( A1 => n21026, A2 => n19501, B1 => n21020, B2 =>
                           n9149, C1 => n21014, C2 => n8765, ZN => n17027);
   U15812 : OAI221_X1 port map( B1 => n14121, B2 => n21038, C1 => n15652, C2 =>
                           n21032, A => n17008, ZN => n17001);
   U15813 : AOI222_X1 port map( A1 => n21026, A2 => n19481, B1 => n21020, B2 =>
                           n9145, C1 => n21014, C2 => n8761, ZN => n17008);
   U15814 : OAI221_X1 port map( B1 => n14120, B2 => n21038, C1 => n15651, C2 =>
                           n21032, A => n16989, ZN => n16982);
   U15815 : AOI222_X1 port map( A1 => n21026, A2 => n19461, B1 => n21020, B2 =>
                           n9141, C1 => n21014, C2 => n8757, ZN => n16989);
   U15816 : OAI221_X1 port map( B1 => n14119, B2 => n21038, C1 => n15650, C2 =>
                           n21032, A => n16970, ZN => n16963);
   U15817 : AOI222_X1 port map( A1 => n21026, A2 => n19441, B1 => n21020, B2 =>
                           n9137, C1 => n21014, C2 => n8753, ZN => n16970);
   U15818 : OAI221_X1 port map( B1 => n14118, B2 => n21038, C1 => n15649, C2 =>
                           n21032, A => n16951, ZN => n16944);
   U15819 : AOI222_X1 port map( A1 => n21026, A2 => n19421, B1 => n21020, B2 =>
                           n9133, C1 => n21014, C2 => n8749, ZN => n16951);
   U15820 : OAI221_X1 port map( B1 => n14117, B2 => n21038, C1 => n15648, C2 =>
                           n21032, A => n16932, ZN => n16925);
   U15821 : AOI222_X1 port map( A1 => n21026, A2 => n19401, B1 => n21020, B2 =>
                           n9129, C1 => n21014, C2 => n8745, ZN => n16932);
   U15822 : OAI221_X1 port map( B1 => n14116, B2 => n21038, C1 => n15647, C2 =>
                           n21032, A => n16913, ZN => n16906);
   U15823 : AOI222_X1 port map( A1 => n21026, A2 => n19381, B1 => n21020, B2 =>
                           n9125, C1 => n21014, C2 => n8741, ZN => n16913);
   U15824 : OAI221_X1 port map( B1 => n14115, B2 => n21038, C1 => n15646, C2 =>
                           n21032, A => n16894, ZN => n16887);
   U15825 : AOI222_X1 port map( A1 => n21026, A2 => n19361, B1 => n21020, B2 =>
                           n9121, C1 => n21014, C2 => n8737, ZN => n16894);
   U15826 : OAI221_X1 port map( B1 => n14114, B2 => n21038, C1 => n15645, C2 =>
                           n21032, A => n16875, ZN => n16868);
   U15827 : AOI222_X1 port map( A1 => n21026, A2 => n19341, B1 => n21020, B2 =>
                           n9117, C1 => n21014, C2 => n8733, ZN => n16875);
   U15828 : OAI221_X1 port map( B1 => n14113, B2 => n21039, C1 => n15644, C2 =>
                           n21033, A => n16856, ZN => n16849);
   U15829 : AOI222_X1 port map( A1 => n21027, A2 => n19321, B1 => n21021, B2 =>
                           n9113, C1 => n21015, C2 => n8729, ZN => n16856);
   U15830 : OAI221_X1 port map( B1 => n14112, B2 => n21039, C1 => n15643, C2 =>
                           n21033, A => n16837, ZN => n16830);
   U15831 : AOI222_X1 port map( A1 => n21027, A2 => n19301, B1 => n21021, B2 =>
                           n9109, C1 => n21015, C2 => n8725, ZN => n16837);
   U15832 : OAI221_X1 port map( B1 => n14111, B2 => n21039, C1 => n15642, C2 =>
                           n21033, A => n16818, ZN => n16811);
   U15833 : AOI222_X1 port map( A1 => n21027, A2 => n19281, B1 => n21021, B2 =>
                           n9105, C1 => n21015, C2 => n8721, ZN => n16818);
   U15834 : OAI221_X1 port map( B1 => n14110, B2 => n21039, C1 => n15641, C2 =>
                           n21033, A => n16799, ZN => n16792);
   U15835 : AOI222_X1 port map( A1 => n21027, A2 => n19261, B1 => n21021, B2 =>
                           n9101, C1 => n21015, C2 => n8717, ZN => n16799);
   U15836 : OAI221_X1 port map( B1 => n14109, B2 => n21039, C1 => n15640, C2 =>
                           n21033, A => n16780, ZN => n16773);
   U15837 : AOI222_X1 port map( A1 => n21027, A2 => n19241, B1 => n21021, B2 =>
                           n9097, C1 => n21015, C2 => n8713, ZN => n16780);
   U15838 : OAI221_X1 port map( B1 => n14108, B2 => n21039, C1 => n15639, C2 =>
                           n21033, A => n16761, ZN => n16754);
   U15839 : AOI222_X1 port map( A1 => n21027, A2 => n19221, B1 => n21021, B2 =>
                           n9093, C1 => n21015, C2 => n8709, ZN => n16761);
   U15840 : OAI221_X1 port map( B1 => n14107, B2 => n21039, C1 => n15638, C2 =>
                           n21033, A => n16742, ZN => n16735);
   U15841 : AOI222_X1 port map( A1 => n21027, A2 => n19201, B1 => n21021, B2 =>
                           n9089, C1 => n21015, C2 => n8705, ZN => n16742);
   U15842 : OAI221_X1 port map( B1 => n14106, B2 => n21039, C1 => n15637, C2 =>
                           n21033, A => n16723, ZN => n16716);
   U15843 : AOI222_X1 port map( A1 => n21027, A2 => n19181, B1 => n21021, B2 =>
                           n9085, C1 => n21015, C2 => n8701, ZN => n16723);
   U15844 : OAI221_X1 port map( B1 => n14105, B2 => n21039, C1 => n15636, C2 =>
                           n21033, A => n16704, ZN => n16697);
   U15845 : AOI222_X1 port map( A1 => n21027, A2 => n19161, B1 => n21021, B2 =>
                           n9081, C1 => n21015, C2 => n8697, ZN => n16704);
   U15846 : OAI221_X1 port map( B1 => n14104, B2 => n21039, C1 => n15635, C2 =>
                           n21033, A => n16685, ZN => n16678);
   U15847 : AOI222_X1 port map( A1 => n21027, A2 => n19141, B1 => n21021, B2 =>
                           n9077, C1 => n21015, C2 => n8693, ZN => n16685);
   U15848 : OAI221_X1 port map( B1 => n14103, B2 => n21039, C1 => n15634, C2 =>
                           n21033, A => n16666, ZN => n16659);
   U15849 : AOI222_X1 port map( A1 => n21027, A2 => n19121, B1 => n21021, B2 =>
                           n9073, C1 => n21015, C2 => n8689, ZN => n16666);
   U15850 : OAI221_X1 port map( B1 => n14102, B2 => n21039, C1 => n15633, C2 =>
                           n21033, A => n16647, ZN => n16640);
   U15851 : AOI222_X1 port map( A1 => n21027, A2 => n19101, B1 => n21021, B2 =>
                           n9069, C1 => n21015, C2 => n8685, ZN => n16647);
   U15852 : OAI221_X1 port map( B1 => n14101, B2 => n21040, C1 => n15632, C2 =>
                           n21034, A => n16628, ZN => n16621);
   U15853 : AOI222_X1 port map( A1 => n21028, A2 => n19081, B1 => n21022, B2 =>
                           n9065, C1 => n21016, C2 => n8681, ZN => n16628);
   U15854 : OAI221_X1 port map( B1 => n14100, B2 => n21040, C1 => n15631, C2 =>
                           n21034, A => n16609, ZN => n16602);
   U15855 : AOI222_X1 port map( A1 => n21028, A2 => n19061, B1 => n21022, B2 =>
                           n9061, C1 => n21016, C2 => n8677, ZN => n16609);
   U15856 : OAI221_X1 port map( B1 => n14099, B2 => n21040, C1 => n15630, C2 =>
                           n21034, A => n16590, ZN => n16583);
   U15857 : AOI222_X1 port map( A1 => n21028, A2 => n19041, B1 => n21022, B2 =>
                           n9057, C1 => n21016, C2 => n8673, ZN => n16590);
   U15858 : OAI221_X1 port map( B1 => n14098, B2 => n21040, C1 => n15629, C2 =>
                           n21034, A => n16571, ZN => n16564);
   U15859 : AOI222_X1 port map( A1 => n21028, A2 => n19021, B1 => n21022, B2 =>
                           n9053, C1 => n21016, C2 => n8669, ZN => n16571);
   U15860 : OAI221_X1 port map( B1 => n14097, B2 => n21040, C1 => n15628, C2 =>
                           n21034, A => n16552, ZN => n16545);
   U15861 : AOI222_X1 port map( A1 => n21028, A2 => n19001, B1 => n21022, B2 =>
                           n9049, C1 => n21016, C2 => n8665, ZN => n16552);
   U15862 : OAI221_X1 port map( B1 => n14096, B2 => n21040, C1 => n15627, C2 =>
                           n21034, A => n16533, ZN => n16526);
   U15863 : AOI222_X1 port map( A1 => n21028, A2 => n18981, B1 => n21022, B2 =>
                           n9045, C1 => n21016, C2 => n8661, ZN => n16533);
   U15864 : OAI221_X1 port map( B1 => n14095, B2 => n21040, C1 => n15626, C2 =>
                           n21034, A => n16514, ZN => n16507);
   U15865 : AOI222_X1 port map( A1 => n21028, A2 => n18961, B1 => n21022, B2 =>
                           n9041, C1 => n21016, C2 => n8657, ZN => n16514);
   U15866 : OAI221_X1 port map( B1 => n14094, B2 => n21040, C1 => n15625, C2 =>
                           n21034, A => n16495, ZN => n16488);
   U15867 : AOI222_X1 port map( A1 => n21028, A2 => n18941, B1 => n21022, B2 =>
                           n9037, C1 => n21016, C2 => n8653, ZN => n16495);
   U15868 : OAI221_X1 port map( B1 => n14093, B2 => n21040, C1 => n15624, C2 =>
                           n21034, A => n16476, ZN => n16469);
   U15869 : AOI222_X1 port map( A1 => n21028, A2 => n18921, B1 => n21022, B2 =>
                           n9033, C1 => n21016, C2 => n8649, ZN => n16476);
   U15870 : OAI221_X1 port map( B1 => n14092, B2 => n21040, C1 => n15623, C2 =>
                           n21034, A => n16457, ZN => n16450);
   U15871 : AOI222_X1 port map( A1 => n21028, A2 => n18901, B1 => n21022, B2 =>
                           n9029, C1 => n21016, C2 => n8645, ZN => n16457);
   U15872 : OAI221_X1 port map( B1 => n14091, B2 => n21040, C1 => n15622, C2 =>
                           n21034, A => n16438, ZN => n16431);
   U15873 : AOI222_X1 port map( A1 => n21028, A2 => n18881, B1 => n21022, B2 =>
                           n9025, C1 => n21016, C2 => n8641, ZN => n16438);
   U15874 : OAI221_X1 port map( B1 => n14090, B2 => n21040, C1 => n15621, C2 =>
                           n21034, A => n16419, ZN => n16412);
   U15875 : AOI222_X1 port map( A1 => n21028, A2 => n18861, B1 => n21022, B2 =>
                           n9021, C1 => n21016, C2 => n8637, ZN => n16419);
   U15876 : OAI221_X1 port map( B1 => n14089, B2 => n21041, C1 => n15620, C2 =>
                           n21035, A => n16400, ZN => n16393);
   U15877 : AOI222_X1 port map( A1 => n21029, A2 => n18841, B1 => n21023, B2 =>
                           n9017, C1 => n21017, C2 => n8633, ZN => n16400);
   U15878 : OAI221_X1 port map( B1 => n14088, B2 => n21041, C1 => n15619, C2 =>
                           n21035, A => n16381, ZN => n16374);
   U15879 : AOI222_X1 port map( A1 => n21029, A2 => n18821, B1 => n21023, B2 =>
                           n9013, C1 => n21017, C2 => n8629, ZN => n16381);
   U15880 : OAI221_X1 port map( B1 => n14087, B2 => n21041, C1 => n15618, C2 =>
                           n21035, A => n16362, ZN => n16355);
   U15881 : AOI222_X1 port map( A1 => n21029, A2 => n18801, B1 => n21023, B2 =>
                           n9009, C1 => n21017, C2 => n8625, ZN => n16362);
   U15882 : OAI221_X1 port map( B1 => n14086, B2 => n21041, C1 => n15617, C2 =>
                           n21035, A => n16343, ZN => n16336);
   U15883 : AOI222_X1 port map( A1 => n21029, A2 => n18781, B1 => n21023, B2 =>
                           n9005, C1 => n21017, C2 => n8621, ZN => n16343);
   U15884 : OAI221_X1 port map( B1 => n14085, B2 => n21041, C1 => n15616, C2 =>
                           n21035, A => n16324, ZN => n16317);
   U15885 : AOI222_X1 port map( A1 => n21029, A2 => n18761, B1 => n21023, B2 =>
                           n9001, C1 => n21017, C2 => n8617, ZN => n16324);
   U15886 : OAI221_X1 port map( B1 => n14084, B2 => n21041, C1 => n15615, C2 =>
                           n21035, A => n16305, ZN => n16298);
   U15887 : AOI222_X1 port map( A1 => n21029, A2 => n18741, B1 => n21023, B2 =>
                           n8997, C1 => n21017, C2 => n8613, ZN => n16305);
   U15888 : OAI221_X1 port map( B1 => n14083, B2 => n21041, C1 => n15614, C2 =>
                           n21035, A => n16286, ZN => n16279);
   U15889 : AOI222_X1 port map( A1 => n21029, A2 => n18721, B1 => n21023, B2 =>
                           n8993, C1 => n21017, C2 => n8609, ZN => n16286);
   U15890 : OAI221_X1 port map( B1 => n14082, B2 => n21041, C1 => n15613, C2 =>
                           n21035, A => n16267, ZN => n16260);
   U15891 : AOI222_X1 port map( A1 => n21029, A2 => n18701, B1 => n21023, B2 =>
                           n8989, C1 => n21017, C2 => n8605, ZN => n16267);
   U15892 : OAI221_X1 port map( B1 => n14081, B2 => n21041, C1 => n15612, C2 =>
                           n21035, A => n16248, ZN => n16241);
   U15893 : AOI222_X1 port map( A1 => n21029, A2 => n18681, B1 => n21023, B2 =>
                           n8985, C1 => n21017, C2 => n8601, ZN => n16248);
   U15894 : OAI221_X1 port map( B1 => n14080, B2 => n21041, C1 => n15611, C2 =>
                           n21035, A => n16229, ZN => n16222);
   U15895 : AOI222_X1 port map( A1 => n21029, A2 => n18661, B1 => n21023, B2 =>
                           n8981, C1 => n21017, C2 => n8597, ZN => n16229);
   U15896 : OAI221_X1 port map( B1 => n14079, B2 => n21041, C1 => n15610, C2 =>
                           n21035, A => n16210, ZN => n16203);
   U15897 : AOI222_X1 port map( A1 => n21029, A2 => n18641, B1 => n21023, B2 =>
                           n8977, C1 => n21017, C2 => n8593, ZN => n16210);
   U15898 : OAI221_X1 port map( B1 => n14078, B2 => n21041, C1 => n15609, C2 =>
                           n21035, A => n16191, ZN => n16184);
   U15899 : AOI222_X1 port map( A1 => n21029, A2 => n18621, B1 => n21023, B2 =>
                           n8973, C1 => n21017, C2 => n8589, ZN => n16191);
   U15900 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(3), A3 => n18532,
                           ZN => n18513);
   U15901 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(3), A3 => n17331,
                           ZN => n17312);
   U15902 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n17318);
   U15903 : NAND2_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(1), ZN => n14471);
   U15904 : NAND2_X1 port map( A1 => ADD_WR(2), A2 => n15738, ZN => n14338);
   U15905 : NAND2_X1 port map( A1 => ADD_WR(1), A2 => n15737, ZN => n14205);
   U15906 : OAI221_X1 port map( B1 => n14992, B2 => n20803, C1 => n15058, C2 =>
                           n20797, A => n18303, ZN => n18302);
   U15907 : AOI22_X1 port map( A1 => n20791, A2 => n8932, B1 => n20993, B2 => 
                           OUT2_12_port, ZN => n18303);
   U15908 : OAI221_X1 port map( B1 => n14991, B2 => n20803, C1 => n15057, C2 =>
                           n20797, A => n18285, ZN => n18284);
   U15909 : AOI22_X1 port map( A1 => n20791, A2 => n8930, B1 => n20993, B2 => 
                           OUT2_13_port, ZN => n18285);
   U15910 : OAI221_X1 port map( B1 => n14990, B2 => n20803, C1 => n15056, C2 =>
                           n20797, A => n18267, ZN => n18266);
   U15911 : AOI22_X1 port map( A1 => n20791, A2 => n8928, B1 => n20993, B2 => 
                           OUT2_14_port, ZN => n18267);
   U15912 : OAI221_X1 port map( B1 => n14989, B2 => n20803, C1 => n15055, C2 =>
                           n20797, A => n18249, ZN => n18248);
   U15913 : AOI22_X1 port map( A1 => n20791, A2 => n8926, B1 => n20993, B2 => 
                           OUT2_15_port, ZN => n18249);
   U15914 : OAI221_X1 port map( B1 => n14988, B2 => n20803, C1 => n15054, C2 =>
                           n20797, A => n18231, ZN => n18230);
   U15915 : AOI22_X1 port map( A1 => n20791, A2 => n8924, B1 => n20993, B2 => 
                           OUT2_16_port, ZN => n18231);
   U15916 : OAI221_X1 port map( B1 => n14987, B2 => n20803, C1 => n15053, C2 =>
                           n20797, A => n18213, ZN => n18212);
   U15917 : AOI22_X1 port map( A1 => n20791, A2 => n8922, B1 => n20993, B2 => 
                           OUT2_17_port, ZN => n18213);
   U15918 : OAI221_X1 port map( B1 => n14986, B2 => n20803, C1 => n15052, C2 =>
                           n20797, A => n18195, ZN => n18194);
   U15919 : AOI22_X1 port map( A1 => n20791, A2 => n8920, B1 => n20993, B2 => 
                           OUT2_18_port, ZN => n18195);
   U15920 : OAI221_X1 port map( B1 => n14985, B2 => n20803, C1 => n15051, C2 =>
                           n20797, A => n18177, ZN => n18176);
   U15921 : AOI22_X1 port map( A1 => n20791, A2 => n8918, B1 => n20993, B2 => 
                           OUT2_19_port, ZN => n18177);
   U15922 : OAI221_X1 port map( B1 => n14984, B2 => n20803, C1 => n15050, C2 =>
                           n20797, A => n18159, ZN => n18158);
   U15923 : AOI22_X1 port map( A1 => n20791, A2 => n8916, B1 => n20992, B2 => 
                           OUT2_20_port, ZN => n18159);
   U15924 : OAI221_X1 port map( B1 => n14983, B2 => n20803, C1 => n15049, C2 =>
                           n20797, A => n18141, ZN => n18140);
   U15925 : AOI22_X1 port map( A1 => n20791, A2 => n8914, B1 => n20992, B2 => 
                           OUT2_21_port, ZN => n18141);
   U15926 : OAI221_X1 port map( B1 => n14982, B2 => n20803, C1 => n15048, C2 =>
                           n20797, A => n18123, ZN => n18122);
   U15927 : AOI22_X1 port map( A1 => n20791, A2 => n8912, B1 => n20992, B2 => 
                           OUT2_22_port, ZN => n18123);
   U15928 : OAI221_X1 port map( B1 => n14981, B2 => n20803, C1 => n15047, C2 =>
                           n20797, A => n18105, ZN => n18104);
   U15929 : AOI22_X1 port map( A1 => n20791, A2 => n8910, B1 => n20992, B2 => 
                           OUT2_23_port, ZN => n18105);
   U15930 : OAI221_X1 port map( B1 => n14980, B2 => n20804, C1 => n15046, C2 =>
                           n20798, A => n18087, ZN => n18086);
   U15931 : AOI22_X1 port map( A1 => n20792, A2 => n8908, B1 => n20992, B2 => 
                           OUT2_24_port, ZN => n18087);
   U15932 : OAI221_X1 port map( B1 => n14979, B2 => n20804, C1 => n15045, C2 =>
                           n20798, A => n18069, ZN => n18068);
   U15933 : AOI22_X1 port map( A1 => n20792, A2 => n8906, B1 => n20992, B2 => 
                           OUT2_25_port, ZN => n18069);
   U15934 : OAI221_X1 port map( B1 => n14978, B2 => n20804, C1 => n15044, C2 =>
                           n20798, A => n18051, ZN => n18050);
   U15935 : AOI22_X1 port map( A1 => n20792, A2 => n8904, B1 => n20992, B2 => 
                           OUT2_26_port, ZN => n18051);
   U15936 : OAI221_X1 port map( B1 => n14977, B2 => n20804, C1 => n15043, C2 =>
                           n20798, A => n18033, ZN => n18032);
   U15937 : AOI22_X1 port map( A1 => n20792, A2 => n8902, B1 => n20992, B2 => 
                           OUT2_27_port, ZN => n18033);
   U15938 : OAI221_X1 port map( B1 => n14976, B2 => n20804, C1 => n15042, C2 =>
                           n20798, A => n18015, ZN => n18014);
   U15939 : AOI22_X1 port map( A1 => n20792, A2 => n8900, B1 => n20992, B2 => 
                           OUT2_28_port, ZN => n18015);
   U15940 : OAI221_X1 port map( B1 => n14975, B2 => n20804, C1 => n15041, C2 =>
                           n20798, A => n17997, ZN => n17996);
   U15941 : AOI22_X1 port map( A1 => n20792, A2 => n8898, B1 => n20992, B2 => 
                           OUT2_29_port, ZN => n17997);
   U15942 : OAI221_X1 port map( B1 => n14974, B2 => n20804, C1 => n15040, C2 =>
                           n20798, A => n17979, ZN => n17978);
   U15943 : AOI22_X1 port map( A1 => n20792, A2 => n8896, B1 => n20992, B2 => 
                           OUT2_30_port, ZN => n17979);
   U15944 : OAI221_X1 port map( B1 => n14973, B2 => n20804, C1 => n15039, C2 =>
                           n20798, A => n17961, ZN => n17960);
   U15945 : AOI22_X1 port map( A1 => n20792, A2 => n8894, B1 => n20992, B2 => 
                           OUT2_31_port, ZN => n17961);
   U15946 : OAI221_X1 port map( B1 => n14972, B2 => n20804, C1 => n15038, C2 =>
                           n20798, A => n17943, ZN => n17942);
   U15947 : AOI22_X1 port map( A1 => n20792, A2 => n8892, B1 => n20992, B2 => 
                           OUT2_32_port, ZN => n17943);
   U15948 : OAI221_X1 port map( B1 => n14971, B2 => n20804, C1 => n15037, C2 =>
                           n20798, A => n17925, ZN => n17924);
   U15949 : AOI22_X1 port map( A1 => n20792, A2 => n8890, B1 => n20991, B2 => 
                           OUT2_33_port, ZN => n17925);
   U15950 : OAI221_X1 port map( B1 => n14970, B2 => n20804, C1 => n15036, C2 =>
                           n20798, A => n17907, ZN => n17906);
   U15951 : AOI22_X1 port map( A1 => n20792, A2 => n8888, B1 => n20991, B2 => 
                           OUT2_34_port, ZN => n17907);
   U15952 : OAI221_X1 port map( B1 => n14969, B2 => n20804, C1 => n15035, C2 =>
                           n20798, A => n17889, ZN => n17888);
   U15953 : AOI22_X1 port map( A1 => n20792, A2 => n8886, B1 => n20991, B2 => 
                           OUT2_35_port, ZN => n17889);
   U15954 : OAI221_X1 port map( B1 => n14968, B2 => n20805, C1 => n15034, C2 =>
                           n20799, A => n17871, ZN => n17870);
   U15955 : AOI22_X1 port map( A1 => n20793, A2 => n8884, B1 => n20991, B2 => 
                           OUT2_36_port, ZN => n17871);
   U15956 : OAI221_X1 port map( B1 => n14967, B2 => n20805, C1 => n15033, C2 =>
                           n20799, A => n17853, ZN => n17852);
   U15957 : AOI22_X1 port map( A1 => n20793, A2 => n8882, B1 => n20991, B2 => 
                           OUT2_37_port, ZN => n17853);
   U15958 : OAI221_X1 port map( B1 => n14966, B2 => n20805, C1 => n15032, C2 =>
                           n20799, A => n17835, ZN => n17834);
   U15959 : AOI22_X1 port map( A1 => n20793, A2 => n8880, B1 => n20991, B2 => 
                           OUT2_38_port, ZN => n17835);
   U15960 : OAI221_X1 port map( B1 => n14965, B2 => n20805, C1 => n15031, C2 =>
                           n20799, A => n17817, ZN => n17816);
   U15961 : AOI22_X1 port map( A1 => n20793, A2 => n8878, B1 => n20991, B2 => 
                           OUT2_39_port, ZN => n17817);
   U15962 : OAI221_X1 port map( B1 => n14964, B2 => n20805, C1 => n15030, C2 =>
                           n20799, A => n17799, ZN => n17798);
   U15963 : AOI22_X1 port map( A1 => n20793, A2 => n8876, B1 => n20991, B2 => 
                           OUT2_40_port, ZN => n17799);
   U15964 : OAI221_X1 port map( B1 => n14963, B2 => n20805, C1 => n15029, C2 =>
                           n20799, A => n17781, ZN => n17780);
   U15965 : AOI22_X1 port map( A1 => n20793, A2 => n8874, B1 => n20991, B2 => 
                           OUT2_41_port, ZN => n17781);
   U15966 : OAI221_X1 port map( B1 => n14962, B2 => n20805, C1 => n15028, C2 =>
                           n20799, A => n17763, ZN => n17762);
   U15967 : AOI22_X1 port map( A1 => n20793, A2 => n8872, B1 => n20991, B2 => 
                           OUT2_42_port, ZN => n17763);
   U15968 : OAI221_X1 port map( B1 => n14961, B2 => n20805, C1 => n15027, C2 =>
                           n20799, A => n17745, ZN => n17744);
   U15969 : AOI22_X1 port map( A1 => n20793, A2 => n8870, B1 => n20991, B2 => 
                           OUT2_43_port, ZN => n17745);
   U15970 : OAI221_X1 port map( B1 => n14960, B2 => n20805, C1 => n15026, C2 =>
                           n20799, A => n17727, ZN => n17726);
   U15971 : AOI22_X1 port map( A1 => n20793, A2 => n8868, B1 => n20991, B2 => 
                           OUT2_44_port, ZN => n17727);
   U15972 : OAI221_X1 port map( B1 => n14959, B2 => n20805, C1 => n15025, C2 =>
                           n20799, A => n17709, ZN => n17708);
   U15973 : AOI22_X1 port map( A1 => n20793, A2 => n8866, B1 => n20991, B2 => 
                           OUT2_45_port, ZN => n17709);
   U15974 : OAI221_X1 port map( B1 => n14958, B2 => n20805, C1 => n15024, C2 =>
                           n20799, A => n17691, ZN => n17690);
   U15975 : AOI22_X1 port map( A1 => n20793, A2 => n8864, B1 => n20990, B2 => 
                           OUT2_46_port, ZN => n17691);
   U15976 : OAI221_X1 port map( B1 => n14957, B2 => n20805, C1 => n15023, C2 =>
                           n20799, A => n17673, ZN => n17672);
   U15977 : AOI22_X1 port map( A1 => n20793, A2 => n8862, B1 => n20990, B2 => 
                           OUT2_47_port, ZN => n17673);
   U15978 : OAI221_X1 port map( B1 => n14956, B2 => n20806, C1 => n15022, C2 =>
                           n20800, A => n17655, ZN => n17654);
   U15979 : AOI22_X1 port map( A1 => n20794, A2 => n8860, B1 => n20990, B2 => 
                           OUT2_48_port, ZN => n17655);
   U15980 : OAI221_X1 port map( B1 => n14955, B2 => n20806, C1 => n15021, C2 =>
                           n20800, A => n17637, ZN => n17636);
   U15981 : AOI22_X1 port map( A1 => n20794, A2 => n8858, B1 => n20990, B2 => 
                           OUT2_49_port, ZN => n17637);
   U15982 : OAI221_X1 port map( B1 => n14954, B2 => n20806, C1 => n15020, C2 =>
                           n20800, A => n17619, ZN => n17618);
   U15983 : AOI22_X1 port map( A1 => n20794, A2 => n8856, B1 => n20990, B2 => 
                           OUT2_50_port, ZN => n17619);
   U15984 : OAI221_X1 port map( B1 => n14953, B2 => n20806, C1 => n15019, C2 =>
                           n20800, A => n17601, ZN => n17600);
   U15985 : AOI22_X1 port map( A1 => n20794, A2 => n8854, B1 => n20990, B2 => 
                           OUT2_51_port, ZN => n17601);
   U15986 : OAI221_X1 port map( B1 => n14952, B2 => n20806, C1 => n15018, C2 =>
                           n20800, A => n17583, ZN => n17582);
   U15987 : AOI22_X1 port map( A1 => n20794, A2 => n8852, B1 => n20990, B2 => 
                           OUT2_52_port, ZN => n17583);
   U15988 : OAI221_X1 port map( B1 => n14951, B2 => n20806, C1 => n15017, C2 =>
                           n20800, A => n17565, ZN => n17564);
   U15989 : AOI22_X1 port map( A1 => n20794, A2 => n8850, B1 => n20990, B2 => 
                           OUT2_53_port, ZN => n17565);
   U15990 : OAI221_X1 port map( B1 => n14950, B2 => n20806, C1 => n15016, C2 =>
                           n20800, A => n17547, ZN => n17546);
   U15991 : AOI22_X1 port map( A1 => n20794, A2 => n8848, B1 => n20990, B2 => 
                           OUT2_54_port, ZN => n17547);
   U15992 : OAI221_X1 port map( B1 => n14949, B2 => n20806, C1 => n15015, C2 =>
                           n20800, A => n17529, ZN => n17528);
   U15993 : AOI22_X1 port map( A1 => n20794, A2 => n8846, B1 => n20990, B2 => 
                           OUT2_55_port, ZN => n17529);
   U15994 : OAI221_X1 port map( B1 => n14948, B2 => n20806, C1 => n15014, C2 =>
                           n20800, A => n17511, ZN => n17510);
   U15995 : AOI22_X1 port map( A1 => n20794, A2 => n8844, B1 => n20990, B2 => 
                           OUT2_56_port, ZN => n17511);
   U15996 : OAI221_X1 port map( B1 => n14947, B2 => n20806, C1 => n15013, C2 =>
                           n20800, A => n17493, ZN => n17492);
   U15997 : AOI22_X1 port map( A1 => n20794, A2 => n8842, B1 => n20990, B2 => 
                           OUT2_57_port, ZN => n17493);
   U15998 : OAI221_X1 port map( B1 => n14946, B2 => n20806, C1 => n15012, C2 =>
                           n20800, A => n17475, ZN => n17474);
   U15999 : AOI22_X1 port map( A1 => n20794, A2 => n8840, B1 => n20990, B2 => 
                           OUT2_58_port, ZN => n17475);
   U16000 : OAI221_X1 port map( B1 => n14945, B2 => n20806, C1 => n15011, C2 =>
                           n20800, A => n17457, ZN => n17456);
   U16001 : AOI22_X1 port map( A1 => n20794, A2 => n8838, B1 => n20989, B2 => 
                           OUT2_59_port, ZN => n17457);
   U16002 : OAI221_X1 port map( B1 => n14992, B2 => n21008, C1 => n15058, C2 =>
                           n21002, A => n17089, ZN => n17088);
   U16003 : AOI22_X1 port map( A1 => n20996, A2 => n8932, B1 => n20988, B2 => 
                           OUT1_12_port, ZN => n17089);
   U16004 : OAI221_X1 port map( B1 => n14991, B2 => n21008, C1 => n15057, C2 =>
                           n21002, A => n17070, ZN => n17069);
   U16005 : AOI22_X1 port map( A1 => n20996, A2 => n8930, B1 => n20988, B2 => 
                           OUT1_13_port, ZN => n17070);
   U16006 : OAI221_X1 port map( B1 => n14990, B2 => n21008, C1 => n15056, C2 =>
                           n21002, A => n17051, ZN => n17050);
   U16007 : AOI22_X1 port map( A1 => n20996, A2 => n8928, B1 => n20988, B2 => 
                           OUT1_14_port, ZN => n17051);
   U16008 : OAI221_X1 port map( B1 => n14989, B2 => n21008, C1 => n15055, C2 =>
                           n21002, A => n17032, ZN => n17031);
   U16009 : AOI22_X1 port map( A1 => n20996, A2 => n8926, B1 => n20988, B2 => 
                           OUT1_15_port, ZN => n17032);
   U16010 : OAI221_X1 port map( B1 => n14988, B2 => n21008, C1 => n15054, C2 =>
                           n21002, A => n17013, ZN => n17012);
   U16011 : AOI22_X1 port map( A1 => n20996, A2 => n8924, B1 => n20988, B2 => 
                           OUT1_16_port, ZN => n17013);
   U16012 : OAI221_X1 port map( B1 => n14987, B2 => n21008, C1 => n15053, C2 =>
                           n21002, A => n16994, ZN => n16993);
   U16013 : AOI22_X1 port map( A1 => n20996, A2 => n8922, B1 => n20988, B2 => 
                           OUT1_17_port, ZN => n16994);
   U16014 : OAI221_X1 port map( B1 => n14986, B2 => n21008, C1 => n15052, C2 =>
                           n21002, A => n16975, ZN => n16974);
   U16015 : AOI22_X1 port map( A1 => n20996, A2 => n8920, B1 => n20988, B2 => 
                           OUT1_18_port, ZN => n16975);
   U16016 : OAI221_X1 port map( B1 => n14985, B2 => n21008, C1 => n15051, C2 =>
                           n21002, A => n16956, ZN => n16955);
   U16017 : AOI22_X1 port map( A1 => n20996, A2 => n8918, B1 => n20987, B2 => 
                           OUT1_19_port, ZN => n16956);
   U16018 : OAI221_X1 port map( B1 => n14984, B2 => n21008, C1 => n15050, C2 =>
                           n21002, A => n16937, ZN => n16936);
   U16019 : AOI22_X1 port map( A1 => n20996, A2 => n8916, B1 => n20987, B2 => 
                           OUT1_20_port, ZN => n16937);
   U16020 : OAI221_X1 port map( B1 => n14983, B2 => n21008, C1 => n15049, C2 =>
                           n21002, A => n16918, ZN => n16917);
   U16021 : AOI22_X1 port map( A1 => n20996, A2 => n8914, B1 => n20987, B2 => 
                           OUT1_21_port, ZN => n16918);
   U16022 : OAI221_X1 port map( B1 => n14982, B2 => n21008, C1 => n15048, C2 =>
                           n21002, A => n16899, ZN => n16898);
   U16023 : AOI22_X1 port map( A1 => n20996, A2 => n8912, B1 => n20987, B2 => 
                           OUT1_22_port, ZN => n16899);
   U16024 : OAI221_X1 port map( B1 => n14981, B2 => n21008, C1 => n15047, C2 =>
                           n21002, A => n16880, ZN => n16879);
   U16025 : AOI22_X1 port map( A1 => n20996, A2 => n8910, B1 => n20987, B2 => 
                           OUT1_23_port, ZN => n16880);
   U16026 : OAI221_X1 port map( B1 => n14980, B2 => n21009, C1 => n15046, C2 =>
                           n21003, A => n16861, ZN => n16860);
   U16027 : AOI22_X1 port map( A1 => n20997, A2 => n8908, B1 => n20987, B2 => 
                           OUT1_24_port, ZN => n16861);
   U16028 : OAI221_X1 port map( B1 => n14979, B2 => n21009, C1 => n15045, C2 =>
                           n21003, A => n16842, ZN => n16841);
   U16029 : AOI22_X1 port map( A1 => n20997, A2 => n8906, B1 => n20987, B2 => 
                           OUT1_25_port, ZN => n16842);
   U16030 : OAI221_X1 port map( B1 => n14978, B2 => n21009, C1 => n15044, C2 =>
                           n21003, A => n16823, ZN => n16822);
   U16031 : AOI22_X1 port map( A1 => n20997, A2 => n8904, B1 => n20987, B2 => 
                           OUT1_26_port, ZN => n16823);
   U16032 : OAI221_X1 port map( B1 => n14977, B2 => n21009, C1 => n15043, C2 =>
                           n21003, A => n16804, ZN => n16803);
   U16033 : AOI22_X1 port map( A1 => n20997, A2 => n8902, B1 => n20987, B2 => 
                           OUT1_27_port, ZN => n16804);
   U16034 : OAI221_X1 port map( B1 => n14976, B2 => n21009, C1 => n15042, C2 =>
                           n21003, A => n16785, ZN => n16784);
   U16035 : AOI22_X1 port map( A1 => n20997, A2 => n8900, B1 => n20989, B2 => 
                           OUT1_28_port, ZN => n16785);
   U16036 : OAI221_X1 port map( B1 => n14975, B2 => n21009, C1 => n15041, C2 =>
                           n21003, A => n16766, ZN => n16765);
   U16037 : AOI22_X1 port map( A1 => n20997, A2 => n8898, B1 => n20987, B2 => 
                           OUT1_29_port, ZN => n16766);
   U16038 : OAI221_X1 port map( B1 => n14974, B2 => n21009, C1 => n15040, C2 =>
                           n21003, A => n16747, ZN => n16746);
   U16039 : AOI22_X1 port map( A1 => n20997, A2 => n8896, B1 => n20987, B2 => 
                           OUT1_30_port, ZN => n16747);
   U16040 : OAI221_X1 port map( B1 => n14973, B2 => n21009, C1 => n15039, C2 =>
                           n21003, A => n16728, ZN => n16727);
   U16041 : AOI22_X1 port map( A1 => n20997, A2 => n8894, B1 => n20986, B2 => 
                           OUT1_31_port, ZN => n16728);
   U16042 : OAI221_X1 port map( B1 => n14972, B2 => n21009, C1 => n15038, C2 =>
                           n21003, A => n16709, ZN => n16708);
   U16043 : AOI22_X1 port map( A1 => n20997, A2 => n8892, B1 => n20987, B2 => 
                           OUT1_32_port, ZN => n16709);
   U16044 : OAI221_X1 port map( B1 => n14971, B2 => n21009, C1 => n15037, C2 =>
                           n21003, A => n16690, ZN => n16689);
   U16045 : AOI22_X1 port map( A1 => n20997, A2 => n8890, B1 => n20986, B2 => 
                           OUT1_33_port, ZN => n16690);
   U16046 : OAI221_X1 port map( B1 => n14970, B2 => n21009, C1 => n15036, C2 =>
                           n21003, A => n16671, ZN => n16670);
   U16047 : AOI22_X1 port map( A1 => n20997, A2 => n8888, B1 => n20986, B2 => 
                           OUT1_34_port, ZN => n16671);
   U16048 : OAI221_X1 port map( B1 => n14969, B2 => n21009, C1 => n15035, C2 =>
                           n21003, A => n16652, ZN => n16651);
   U16049 : AOI22_X1 port map( A1 => n20997, A2 => n8886, B1 => n20986, B2 => 
                           OUT1_35_port, ZN => n16652);
   U16050 : OAI221_X1 port map( B1 => n14968, B2 => n21010, C1 => n15034, C2 =>
                           n21004, A => n16633, ZN => n16632);
   U16051 : AOI22_X1 port map( A1 => n20998, A2 => n8884, B1 => n20986, B2 => 
                           OUT1_36_port, ZN => n16633);
   U16052 : OAI221_X1 port map( B1 => n14967, B2 => n21010, C1 => n15033, C2 =>
                           n21004, A => n16614, ZN => n16613);
   U16053 : AOI22_X1 port map( A1 => n20998, A2 => n8882, B1 => n20986, B2 => 
                           OUT1_37_port, ZN => n16614);
   U16054 : OAI221_X1 port map( B1 => n14966, B2 => n21010, C1 => n15032, C2 =>
                           n21004, A => n16595, ZN => n16594);
   U16055 : AOI22_X1 port map( A1 => n20998, A2 => n8880, B1 => n20986, B2 => 
                           OUT1_38_port, ZN => n16595);
   U16056 : OAI221_X1 port map( B1 => n14965, B2 => n21010, C1 => n15031, C2 =>
                           n21004, A => n16576, ZN => n16575);
   U16057 : AOI22_X1 port map( A1 => n20998, A2 => n8878, B1 => n20986, B2 => 
                           OUT1_39_port, ZN => n16576);
   U16058 : OAI221_X1 port map( B1 => n14964, B2 => n21010, C1 => n15030, C2 =>
                           n21004, A => n16557, ZN => n16556);
   U16059 : AOI22_X1 port map( A1 => n20998, A2 => n8876, B1 => n20986, B2 => 
                           OUT1_40_port, ZN => n16557);
   U16060 : OAI221_X1 port map( B1 => n14963, B2 => n21010, C1 => n15029, C2 =>
                           n21004, A => n16538, ZN => n16537);
   U16061 : AOI22_X1 port map( A1 => n20998, A2 => n8874, B1 => n20986, B2 => 
                           OUT1_41_port, ZN => n16538);
   U16062 : OAI221_X1 port map( B1 => n14962, B2 => n21010, C1 => n15028, C2 =>
                           n21004, A => n16519, ZN => n16518);
   U16063 : AOI22_X1 port map( A1 => n20998, A2 => n8872, B1 => n20986, B2 => 
                           OUT1_42_port, ZN => n16519);
   U16064 : OAI221_X1 port map( B1 => n14961, B2 => n21010, C1 => n15027, C2 =>
                           n21004, A => n16500, ZN => n16499);
   U16065 : AOI22_X1 port map( A1 => n20998, A2 => n8870, B1 => n20986, B2 => 
                           OUT1_43_port, ZN => n16500);
   U16066 : OAI221_X1 port map( B1 => n14960, B2 => n21010, C1 => n15026, C2 =>
                           n21004, A => n16481, ZN => n16480);
   U16067 : AOI22_X1 port map( A1 => n20998, A2 => n8868, B1 => n20986, B2 => 
                           OUT1_44_port, ZN => n16481);
   U16068 : OAI221_X1 port map( B1 => n14959, B2 => n21010, C1 => n15025, C2 =>
                           n21004, A => n16462, ZN => n16461);
   U16069 : AOI22_X1 port map( A1 => n20998, A2 => n8866, B1 => n20985, B2 => 
                           OUT1_45_port, ZN => n16462);
   U16070 : OAI221_X1 port map( B1 => n14958, B2 => n21010, C1 => n15024, C2 =>
                           n21004, A => n16443, ZN => n16442);
   U16071 : AOI22_X1 port map( A1 => n20998, A2 => n8864, B1 => n20985, B2 => 
                           OUT1_46_port, ZN => n16443);
   U16072 : OAI221_X1 port map( B1 => n14957, B2 => n21010, C1 => n15023, C2 =>
                           n21004, A => n16424, ZN => n16423);
   U16073 : AOI22_X1 port map( A1 => n20998, A2 => n8862, B1 => n20985, B2 => 
                           OUT1_47_port, ZN => n16424);
   U16074 : OAI221_X1 port map( B1 => n14956, B2 => n21011, C1 => n15022, C2 =>
                           n21005, A => n16405, ZN => n16404);
   U16075 : AOI22_X1 port map( A1 => n20999, A2 => n8860, B1 => n20985, B2 => 
                           OUT1_48_port, ZN => n16405);
   U16076 : OAI221_X1 port map( B1 => n14955, B2 => n21011, C1 => n15021, C2 =>
                           n21005, A => n16386, ZN => n16385);
   U16077 : AOI22_X1 port map( A1 => n20999, A2 => n8858, B1 => n20985, B2 => 
                           OUT1_49_port, ZN => n16386);
   U16078 : OAI221_X1 port map( B1 => n14954, B2 => n21011, C1 => n15020, C2 =>
                           n21005, A => n16367, ZN => n16366);
   U16079 : AOI22_X1 port map( A1 => n20999, A2 => n8856, B1 => n20985, B2 => 
                           OUT1_50_port, ZN => n16367);
   U16080 : OAI221_X1 port map( B1 => n14953, B2 => n21011, C1 => n15019, C2 =>
                           n21005, A => n16348, ZN => n16347);
   U16081 : AOI22_X1 port map( A1 => n20999, A2 => n8854, B1 => n20985, B2 => 
                           OUT1_51_port, ZN => n16348);
   U16082 : OAI221_X1 port map( B1 => n14952, B2 => n21011, C1 => n15018, C2 =>
                           n21005, A => n16329, ZN => n16328);
   U16083 : AOI22_X1 port map( A1 => n20999, A2 => n8852, B1 => n20985, B2 => 
                           OUT1_52_port, ZN => n16329);
   U16084 : OAI221_X1 port map( B1 => n14951, B2 => n21011, C1 => n15017, C2 =>
                           n21005, A => n16310, ZN => n16309);
   U16085 : AOI22_X1 port map( A1 => n20999, A2 => n8850, B1 => n20985, B2 => 
                           OUT1_53_port, ZN => n16310);
   U16086 : OAI221_X1 port map( B1 => n14950, B2 => n21011, C1 => n15016, C2 =>
                           n21005, A => n16291, ZN => n16290);
   U16087 : AOI22_X1 port map( A1 => n20999, A2 => n8848, B1 => n20985, B2 => 
                           OUT1_54_port, ZN => n16291);
   U16088 : OAI221_X1 port map( B1 => n14949, B2 => n21011, C1 => n15015, C2 =>
                           n21005, A => n16272, ZN => n16271);
   U16089 : AOI22_X1 port map( A1 => n20999, A2 => n8846, B1 => n20985, B2 => 
                           OUT1_55_port, ZN => n16272);
   U16090 : OAI221_X1 port map( B1 => n14948, B2 => n21011, C1 => n15014, C2 =>
                           n21005, A => n16253, ZN => n16252);
   U16091 : AOI22_X1 port map( A1 => n20999, A2 => n8844, B1 => n20985, B2 => 
                           OUT1_56_port, ZN => n16253);
   U16092 : OAI221_X1 port map( B1 => n14947, B2 => n21011, C1 => n15013, C2 =>
                           n21005, A => n16234, ZN => n16233);
   U16093 : AOI22_X1 port map( A1 => n20999, A2 => n8842, B1 => n20984, B2 => 
                           OUT1_57_port, ZN => n16234);
   U16094 : OAI221_X1 port map( B1 => n14946, B2 => n21011, C1 => n15012, C2 =>
                           n21005, A => n16215, ZN => n16214);
   U16095 : AOI22_X1 port map( A1 => n20999, A2 => n8840, B1 => n20985, B2 => 
                           OUT1_58_port, ZN => n16215);
   U16096 : OAI221_X1 port map( B1 => n14945, B2 => n21011, C1 => n15011, C2 =>
                           n21005, A => n16196, ZN => n16195);
   U16097 : AOI22_X1 port map( A1 => n20999, A2 => n8838, B1 => n20984, B2 => 
                           OUT1_59_port, ZN => n16196);
   U16098 : OAI221_X1 port map( B1 => n14344, B2 => n20909, C1 => n14812, C2 =>
                           n20903, A => n17431, ZN => n17430);
   U16099 : AOI22_X1 port map( A1 => n20897, A2 => n18608, B1 => n20891, B2 => 
                           n18609, ZN => n17431);
   U16100 : OAI221_X1 port map( B1 => n14944, B2 => n20807, C1 => n15010, C2 =>
                           n20801, A => n17439, ZN => n17438);
   U16101 : AOI22_X1 port map( A1 => n20795, A2 => n8836, B1 => n20989, B2 => 
                           OUT2_60_port, ZN => n17439);
   U16102 : OAI221_X1 port map( B1 => n14343, B2 => n20909, C1 => n14811, C2 =>
                           n20903, A => n17413, ZN => n17412);
   U16103 : AOI22_X1 port map( A1 => n20897, A2 => n18588, B1 => n20891, B2 => 
                           n18589, ZN => n17413);
   U16104 : OAI221_X1 port map( B1 => n14943, B2 => n20807, C1 => n15009, C2 =>
                           n20801, A => n17421, ZN => n17420);
   U16105 : AOI22_X1 port map( A1 => n20795, A2 => n8834, B1 => n20989, B2 => 
                           OUT2_61_port, ZN => n17421);
   U16106 : OAI221_X1 port map( B1 => n14342, B2 => n20909, C1 => n14810, C2 =>
                           n20903, A => n17395, ZN => n17394);
   U16107 : AOI22_X1 port map( A1 => n20897, A2 => n18568, B1 => n20891, B2 => 
                           n18569, ZN => n17395);
   U16108 : OAI221_X1 port map( B1 => n14942, B2 => n20807, C1 => n15008, C2 =>
                           n20801, A => n17403, ZN => n17402);
   U16109 : AOI22_X1 port map( A1 => n20795, A2 => n8832, B1 => n20989, B2 => 
                           OUT2_62_port, ZN => n17403);
   U16110 : OAI221_X1 port map( B1 => n14340, B2 => n20909, C1 => n14808, C2 =>
                           n20903, A => n17347, ZN => n17344);
   U16111 : AOI22_X1 port map( A1 => n20897, A2 => n18548, B1 => n20891, B2 => 
                           n18549, ZN => n17347);
   U16112 : OAI221_X1 port map( B1 => n14940, B2 => n20807, C1 => n15006, C2 =>
                           n20801, A => n17372, ZN => n17369);
   U16113 : AOI22_X1 port map( A1 => n20795, A2 => n8830, B1 => n20989, B2 => 
                           OUT2_63_port, ZN => n17372);
   U16114 : OAI221_X1 port map( B1 => n14944, B2 => n21012, C1 => n15010, C2 =>
                           n21006, A => n16177, ZN => n16176);
   U16115 : AOI22_X1 port map( A1 => n21000, A2 => n8836, B1 => n20987, B2 => 
                           OUT1_60_port, ZN => n16177);
   U16116 : OAI221_X1 port map( B1 => n14943, B2 => n21012, C1 => n15009, C2 =>
                           n21006, A => n16158, ZN => n16157);
   U16117 : AOI22_X1 port map( A1 => n21000, A2 => n8834, B1 => n20984, B2 => 
                           OUT1_61_port, ZN => n16158);
   U16118 : OAI221_X1 port map( B1 => n14942, B2 => n21012, C1 => n15008, C2 =>
                           n21006, A => n16139, ZN => n16138);
   U16119 : AOI22_X1 port map( A1 => n21000, A2 => n8832, B1 => n20984, B2 => 
                           OUT1_62_port, ZN => n16139);
   U16120 : OAI221_X1 port map( B1 => n14340, B2 => n21115, C1 => n14808, C2 =>
                           n21109, A => n16080, ZN => n16077);
   U16121 : AOI22_X1 port map( A1 => n21103, A2 => n18548, B1 => n21097, B2 => 
                           n18549, ZN => n16080);
   U16122 : OAI221_X1 port map( B1 => n14940, B2 => n21012, C1 => n15006, C2 =>
                           n21006, A => n16106, ZN => n16103);
   U16123 : AOI22_X1 port map( A1 => n21000, A2 => n8830, B1 => n20989, B2 => 
                           OUT1_63_port, ZN => n16106);
   U16124 : OAI221_X1 port map( B1 => n15004, B2 => n20802, C1 => n15070, C2 =>
                           n20796, A => n18530, ZN => n18529);
   U16125 : AOI22_X1 port map( A1 => n20790, A2 => n8956, B1 => n20984, B2 => 
                           OUT2_0_port, ZN => n18530);
   U16126 : OAI221_X1 port map( B1 => n15003, B2 => n20802, C1 => n15069, C2 =>
                           n20796, A => n18501, ZN => n18500);
   U16127 : AOI22_X1 port map( A1 => n20790, A2 => n8954, B1 => n20994, B2 => 
                           OUT2_1_port, ZN => n18501);
   U16128 : OAI221_X1 port map( B1 => n15002, B2 => n20802, C1 => n15068, C2 =>
                           n20796, A => n18483, ZN => n18482);
   U16129 : AOI22_X1 port map( A1 => n20790, A2 => n8952, B1 => n20994, B2 => 
                           OUT2_2_port, ZN => n18483);
   U16130 : OAI221_X1 port map( B1 => n15001, B2 => n20802, C1 => n15067, C2 =>
                           n20796, A => n18465, ZN => n18464);
   U16131 : AOI22_X1 port map( A1 => n20790, A2 => n8950, B1 => n20994, B2 => 
                           OUT2_3_port, ZN => n18465);
   U16132 : OAI221_X1 port map( B1 => n15000, B2 => n20802, C1 => n15066, C2 =>
                           n20796, A => n18447, ZN => n18446);
   U16133 : AOI22_X1 port map( A1 => n20790, A2 => n8948, B1 => n20994, B2 => 
                           OUT2_4_port, ZN => n18447);
   U16134 : OAI221_X1 port map( B1 => n14999, B2 => n20802, C1 => n15065, C2 =>
                           n20796, A => n18429, ZN => n18428);
   U16135 : AOI22_X1 port map( A1 => n20790, A2 => n8946, B1 => n20994, B2 => 
                           OUT2_5_port, ZN => n18429);
   U16136 : OAI221_X1 port map( B1 => n14998, B2 => n20802, C1 => n15064, C2 =>
                           n20796, A => n18411, ZN => n18410);
   U16137 : AOI22_X1 port map( A1 => n20790, A2 => n8944, B1 => n20994, B2 => 
                           OUT2_6_port, ZN => n18411);
   U16138 : OAI221_X1 port map( B1 => n14997, B2 => n20802, C1 => n15063, C2 =>
                           n20796, A => n18393, ZN => n18392);
   U16139 : AOI22_X1 port map( A1 => n20790, A2 => n8942, B1 => n20993, B2 => 
                           OUT2_7_port, ZN => n18393);
   U16140 : OAI221_X1 port map( B1 => n14996, B2 => n20802, C1 => n15062, C2 =>
                           n20796, A => n18375, ZN => n18374);
   U16141 : AOI22_X1 port map( A1 => n20790, A2 => n8940, B1 => n20993, B2 => 
                           OUT2_8_port, ZN => n18375);
   U16142 : OAI221_X1 port map( B1 => n14995, B2 => n20802, C1 => n15061, C2 =>
                           n20796, A => n18357, ZN => n18356);
   U16143 : AOI22_X1 port map( A1 => n20790, A2 => n8938, B1 => n20993, B2 => 
                           OUT2_9_port, ZN => n18357);
   U16144 : OAI221_X1 port map( B1 => n14994, B2 => n20802, C1 => n15060, C2 =>
                           n20796, A => n18339, ZN => n18338);
   U16145 : AOI22_X1 port map( A1 => n20790, A2 => n8936, B1 => n20993, B2 => 
                           OUT2_10_port, ZN => n18339);
   U16146 : OAI221_X1 port map( B1 => n14993, B2 => n20802, C1 => n15059, C2 =>
                           n20796, A => n18321, ZN => n18320);
   U16147 : AOI22_X1 port map( A1 => n20790, A2 => n8934, B1 => n20993, B2 => 
                           OUT2_11_port, ZN => n18321);
   U16148 : OAI221_X1 port map( B1 => n15004, B2 => n21007, C1 => n15070, C2 =>
                           n21001, A => n17329, ZN => n17328);
   U16149 : AOI22_X1 port map( A1 => n20995, A2 => n8956, B1 => n20989, B2 => 
                           OUT1_0_port, ZN => n17329);
   U16150 : OAI221_X1 port map( B1 => n15003, B2 => n21007, C1 => n15069, C2 =>
                           n21001, A => n17298, ZN => n17297);
   U16151 : AOI22_X1 port map( A1 => n20995, A2 => n8954, B1 => n20989, B2 => 
                           OUT1_1_port, ZN => n17298);
   U16152 : OAI221_X1 port map( B1 => n15002, B2 => n21007, C1 => n15068, C2 =>
                           n21001, A => n17279, ZN => n17278);
   U16153 : AOI22_X1 port map( A1 => n20995, A2 => n8952, B1 => n20989, B2 => 
                           OUT1_2_port, ZN => n17279);
   U16154 : OAI221_X1 port map( B1 => n15001, B2 => n21007, C1 => n15067, C2 =>
                           n21001, A => n17260, ZN => n17259);
   U16155 : AOI22_X1 port map( A1 => n20995, A2 => n8950, B1 => n20989, B2 => 
                           OUT1_3_port, ZN => n17260);
   U16156 : OAI221_X1 port map( B1 => n15000, B2 => n21007, C1 => n15066, C2 =>
                           n21001, A => n17241, ZN => n17240);
   U16157 : AOI22_X1 port map( A1 => n20995, A2 => n8948, B1 => n20989, B2 => 
                           OUT1_4_port, ZN => n17241);
   U16158 : OAI221_X1 port map( B1 => n14999, B2 => n21007, C1 => n15065, C2 =>
                           n21001, A => n17222, ZN => n17221);
   U16159 : AOI22_X1 port map( A1 => n20995, A2 => n8946, B1 => n20988, B2 => 
                           OUT1_5_port, ZN => n17222);
   U16160 : OAI221_X1 port map( B1 => n14998, B2 => n21007, C1 => n15064, C2 =>
                           n21001, A => n17203, ZN => n17202);
   U16161 : AOI22_X1 port map( A1 => n20995, A2 => n8944, B1 => n20989, B2 => 
                           OUT1_6_port, ZN => n17203);
   U16162 : OAI221_X1 port map( B1 => n14997, B2 => n21007, C1 => n15063, C2 =>
                           n21001, A => n17184, ZN => n17183);
   U16163 : AOI22_X1 port map( A1 => n20995, A2 => n8942, B1 => n20988, B2 => 
                           OUT1_7_port, ZN => n17184);
   U16164 : OAI221_X1 port map( B1 => n14996, B2 => n21007, C1 => n15062, C2 =>
                           n21001, A => n17165, ZN => n17164);
   U16165 : AOI22_X1 port map( A1 => n20995, A2 => n8940, B1 => n20988, B2 => 
                           OUT1_8_port, ZN => n17165);
   U16166 : OAI221_X1 port map( B1 => n14995, B2 => n21007, C1 => n15061, C2 =>
                           n21001, A => n17146, ZN => n17145);
   U16167 : AOI22_X1 port map( A1 => n20995, A2 => n8938, B1 => n20988, B2 => 
                           OUT1_9_port, ZN => n17146);
   U16168 : OAI221_X1 port map( B1 => n14994, B2 => n21007, C1 => n15060, C2 =>
                           n21001, A => n17127, ZN => n17126);
   U16169 : AOI22_X1 port map( A1 => n20995, A2 => n8936, B1 => n20988, B2 => 
                           OUT1_10_port, ZN => n17127);
   U16170 : OAI221_X1 port map( B1 => n14993, B2 => n21007, C1 => n15059, C2 =>
                           n21001, A => n17108, ZN => n17107);
   U16171 : AOI22_X1 port map( A1 => n20995, A2 => n8934, B1 => n20988, B2 => 
                           OUT1_11_port, ZN => n17108);
   U16172 : OAI221_X1 port map( B1 => n17074, B2 => n20881, C1 => n14325, C2 =>
                           n20875, A => n18296, ZN => n18293);
   U16173 : AOI22_X1 port map( A1 => n20869, A2 => n9164, B1 => n20863, B2 => 
                           n8780, ZN => n18296);
   U16174 : OAI221_X1 port map( B1 => n17055, B2 => n20881, C1 => n14324, C2 =>
                           n20875, A => n18278, ZN => n18275);
   U16175 : AOI22_X1 port map( A1 => n20869, A2 => n9160, B1 => n20863, B2 => 
                           n8776, ZN => n18278);
   U16176 : OAI221_X1 port map( B1 => n17036, B2 => n20881, C1 => n14323, C2 =>
                           n20875, A => n18260, ZN => n18257);
   U16177 : AOI22_X1 port map( A1 => n20869, A2 => n9156, B1 => n20863, B2 => 
                           n8772, ZN => n18260);
   U16178 : OAI221_X1 port map( B1 => n17017, B2 => n20881, C1 => n14322, C2 =>
                           n20875, A => n18242, ZN => n18239);
   U16179 : AOI22_X1 port map( A1 => n20869, A2 => n9152, B1 => n20863, B2 => 
                           n8768, ZN => n18242);
   U16180 : OAI221_X1 port map( B1 => n16998, B2 => n20881, C1 => n14321, C2 =>
                           n20875, A => n18224, ZN => n18221);
   U16181 : AOI22_X1 port map( A1 => n20869, A2 => n9148, B1 => n20863, B2 => 
                           n8764, ZN => n18224);
   U16182 : OAI221_X1 port map( B1 => n16979, B2 => n20881, C1 => n14320, C2 =>
                           n20875, A => n18206, ZN => n18203);
   U16183 : AOI22_X1 port map( A1 => n20869, A2 => n9144, B1 => n20863, B2 => 
                           n8760, ZN => n18206);
   U16184 : OAI221_X1 port map( B1 => n16960, B2 => n20881, C1 => n14319, C2 =>
                           n20875, A => n18188, ZN => n18185);
   U16185 : AOI22_X1 port map( A1 => n20869, A2 => n9140, B1 => n20863, B2 => 
                           n8756, ZN => n18188);
   U16186 : OAI221_X1 port map( B1 => n16941, B2 => n20881, C1 => n14318, C2 =>
                           n20875, A => n18170, ZN => n18167);
   U16187 : AOI22_X1 port map( A1 => n20869, A2 => n9136, B1 => n20863, B2 => 
                           n8752, ZN => n18170);
   U16188 : OAI221_X1 port map( B1 => n16922, B2 => n20881, C1 => n14317, C2 =>
                           n20875, A => n18152, ZN => n18149);
   U16189 : AOI22_X1 port map( A1 => n20869, A2 => n9132, B1 => n20863, B2 => 
                           n8748, ZN => n18152);
   U16190 : OAI221_X1 port map( B1 => n16903, B2 => n20881, C1 => n14316, C2 =>
                           n20875, A => n18134, ZN => n18131);
   U16191 : AOI22_X1 port map( A1 => n20869, A2 => n9128, B1 => n20863, B2 => 
                           n8744, ZN => n18134);
   U16192 : OAI221_X1 port map( B1 => n16884, B2 => n20881, C1 => n14315, C2 =>
                           n20875, A => n18116, ZN => n18113);
   U16193 : AOI22_X1 port map( A1 => n20869, A2 => n9124, B1 => n20863, B2 => 
                           n8740, ZN => n18116);
   U16194 : OAI221_X1 port map( B1 => n16865, B2 => n20881, C1 => n14314, C2 =>
                           n20875, A => n18098, ZN => n18095);
   U16195 : AOI22_X1 port map( A1 => n20869, A2 => n9120, B1 => n20863, B2 => 
                           n8736, ZN => n18098);
   U16196 : OAI221_X1 port map( B1 => n16846, B2 => n20882, C1 => n14313, C2 =>
                           n20876, A => n18080, ZN => n18077);
   U16197 : AOI22_X1 port map( A1 => n20870, A2 => n9116, B1 => n20864, B2 => 
                           n8732, ZN => n18080);
   U16198 : OAI221_X1 port map( B1 => n16827, B2 => n20882, C1 => n14312, C2 =>
                           n20876, A => n18062, ZN => n18059);
   U16199 : AOI22_X1 port map( A1 => n20870, A2 => n9112, B1 => n20864, B2 => 
                           n8728, ZN => n18062);
   U16200 : OAI221_X1 port map( B1 => n16808, B2 => n20882, C1 => n14311, C2 =>
                           n20876, A => n18044, ZN => n18041);
   U16201 : AOI22_X1 port map( A1 => n20870, A2 => n9108, B1 => n20864, B2 => 
                           n8724, ZN => n18044);
   U16202 : OAI221_X1 port map( B1 => n16789, B2 => n20882, C1 => n14310, C2 =>
                           n20876, A => n18026, ZN => n18023);
   U16203 : AOI22_X1 port map( A1 => n20870, A2 => n9104, B1 => n20864, B2 => 
                           n8720, ZN => n18026);
   U16204 : OAI221_X1 port map( B1 => n16770, B2 => n20882, C1 => n14309, C2 =>
                           n20876, A => n18008, ZN => n18005);
   U16205 : AOI22_X1 port map( A1 => n20870, A2 => n9100, B1 => n20864, B2 => 
                           n8716, ZN => n18008);
   U16206 : OAI221_X1 port map( B1 => n16751, B2 => n20882, C1 => n14308, C2 =>
                           n20876, A => n17990, ZN => n17987);
   U16207 : AOI22_X1 port map( A1 => n20870, A2 => n9096, B1 => n20864, B2 => 
                           n8712, ZN => n17990);
   U16208 : OAI221_X1 port map( B1 => n16732, B2 => n20882, C1 => n14307, C2 =>
                           n20876, A => n17972, ZN => n17969);
   U16209 : AOI22_X1 port map( A1 => n20870, A2 => n9092, B1 => n20864, B2 => 
                           n8708, ZN => n17972);
   U16210 : OAI221_X1 port map( B1 => n16713, B2 => n20882, C1 => n14306, C2 =>
                           n20876, A => n17954, ZN => n17951);
   U16211 : AOI22_X1 port map( A1 => n20870, A2 => n9088, B1 => n20864, B2 => 
                           n8704, ZN => n17954);
   U16212 : OAI221_X1 port map( B1 => n16694, B2 => n20882, C1 => n14305, C2 =>
                           n20876, A => n17936, ZN => n17933);
   U16213 : AOI22_X1 port map( A1 => n20870, A2 => n9084, B1 => n20864, B2 => 
                           n8700, ZN => n17936);
   U16214 : OAI221_X1 port map( B1 => n16675, B2 => n20882, C1 => n14304, C2 =>
                           n20876, A => n17918, ZN => n17915);
   U16215 : AOI22_X1 port map( A1 => n20870, A2 => n9080, B1 => n20864, B2 => 
                           n8696, ZN => n17918);
   U16216 : OAI221_X1 port map( B1 => n16656, B2 => n20882, C1 => n14303, C2 =>
                           n20876, A => n17900, ZN => n17897);
   U16217 : AOI22_X1 port map( A1 => n20870, A2 => n9076, B1 => n20864, B2 => 
                           n8692, ZN => n17900);
   U16218 : OAI221_X1 port map( B1 => n16637, B2 => n20882, C1 => n14302, C2 =>
                           n20876, A => n17882, ZN => n17879);
   U16219 : AOI22_X1 port map( A1 => n20870, A2 => n9072, B1 => n20864, B2 => 
                           n8688, ZN => n17882);
   U16220 : OAI221_X1 port map( B1 => n16618, B2 => n20883, C1 => n14301, C2 =>
                           n20877, A => n17864, ZN => n17861);
   U16221 : AOI22_X1 port map( A1 => n20871, A2 => n9068, B1 => n20865, B2 => 
                           n8684, ZN => n17864);
   U16222 : OAI221_X1 port map( B1 => n16599, B2 => n20883, C1 => n14300, C2 =>
                           n20877, A => n17846, ZN => n17843);
   U16223 : AOI22_X1 port map( A1 => n20871, A2 => n9064, B1 => n20865, B2 => 
                           n8680, ZN => n17846);
   U16224 : OAI221_X1 port map( B1 => n16580, B2 => n20883, C1 => n14299, C2 =>
                           n20877, A => n17828, ZN => n17825);
   U16225 : AOI22_X1 port map( A1 => n20871, A2 => n9060, B1 => n20865, B2 => 
                           n8676, ZN => n17828);
   U16226 : OAI221_X1 port map( B1 => n16561, B2 => n20883, C1 => n14298, C2 =>
                           n20877, A => n17810, ZN => n17807);
   U16227 : AOI22_X1 port map( A1 => n20871, A2 => n9056, B1 => n20865, B2 => 
                           n8672, ZN => n17810);
   U16228 : OAI221_X1 port map( B1 => n16542, B2 => n20883, C1 => n14297, C2 =>
                           n20877, A => n17792, ZN => n17789);
   U16229 : AOI22_X1 port map( A1 => n20871, A2 => n9052, B1 => n20865, B2 => 
                           n8668, ZN => n17792);
   U16230 : OAI221_X1 port map( B1 => n16523, B2 => n20883, C1 => n14296, C2 =>
                           n20877, A => n17774, ZN => n17771);
   U16231 : AOI22_X1 port map( A1 => n20871, A2 => n9048, B1 => n20865, B2 => 
                           n8664, ZN => n17774);
   U16232 : OAI221_X1 port map( B1 => n16504, B2 => n20883, C1 => n14295, C2 =>
                           n20877, A => n17756, ZN => n17753);
   U16233 : AOI22_X1 port map( A1 => n20871, A2 => n9044, B1 => n20865, B2 => 
                           n8660, ZN => n17756);
   U16234 : OAI221_X1 port map( B1 => n16485, B2 => n20883, C1 => n14294, C2 =>
                           n20877, A => n17738, ZN => n17735);
   U16235 : AOI22_X1 port map( A1 => n20871, A2 => n9040, B1 => n20865, B2 => 
                           n8656, ZN => n17738);
   U16236 : OAI221_X1 port map( B1 => n16466, B2 => n20883, C1 => n14293, C2 =>
                           n20877, A => n17720, ZN => n17717);
   U16237 : AOI22_X1 port map( A1 => n20871, A2 => n9036, B1 => n20865, B2 => 
                           n8652, ZN => n17720);
   U16238 : OAI221_X1 port map( B1 => n16447, B2 => n20883, C1 => n14292, C2 =>
                           n20877, A => n17702, ZN => n17699);
   U16239 : AOI22_X1 port map( A1 => n20871, A2 => n9032, B1 => n20865, B2 => 
                           n8648, ZN => n17702);
   U16240 : OAI221_X1 port map( B1 => n16428, B2 => n20883, C1 => n14291, C2 =>
                           n20877, A => n17684, ZN => n17681);
   U16241 : AOI22_X1 port map( A1 => n20871, A2 => n9028, B1 => n20865, B2 => 
                           n8644, ZN => n17684);
   U16242 : OAI221_X1 port map( B1 => n16409, B2 => n20883, C1 => n14290, C2 =>
                           n20877, A => n17666, ZN => n17663);
   U16243 : AOI22_X1 port map( A1 => n20871, A2 => n9024, B1 => n20865, B2 => 
                           n8640, ZN => n17666);
   U16244 : OAI221_X1 port map( B1 => n16390, B2 => n20884, C1 => n14289, C2 =>
                           n20878, A => n17648, ZN => n17645);
   U16245 : AOI22_X1 port map( A1 => n20872, A2 => n9020, B1 => n20866, B2 => 
                           n8636, ZN => n17648);
   U16246 : OAI221_X1 port map( B1 => n16371, B2 => n20884, C1 => n14288, C2 =>
                           n20878, A => n17630, ZN => n17627);
   U16247 : AOI22_X1 port map( A1 => n20872, A2 => n9016, B1 => n20866, B2 => 
                           n8632, ZN => n17630);
   U16248 : OAI221_X1 port map( B1 => n16352, B2 => n20884, C1 => n14287, C2 =>
                           n20878, A => n17612, ZN => n17609);
   U16249 : AOI22_X1 port map( A1 => n20872, A2 => n9012, B1 => n20866, B2 => 
                           n8628, ZN => n17612);
   U16250 : OAI221_X1 port map( B1 => n16333, B2 => n20884, C1 => n14286, C2 =>
                           n20878, A => n17594, ZN => n17591);
   U16251 : AOI22_X1 port map( A1 => n20872, A2 => n9008, B1 => n20866, B2 => 
                           n8624, ZN => n17594);
   U16252 : OAI221_X1 port map( B1 => n16314, B2 => n20884, C1 => n14285, C2 =>
                           n20878, A => n17576, ZN => n17573);
   U16253 : AOI22_X1 port map( A1 => n20872, A2 => n9004, B1 => n20866, B2 => 
                           n8620, ZN => n17576);
   U16254 : OAI221_X1 port map( B1 => n16295, B2 => n20884, C1 => n14284, C2 =>
                           n20878, A => n17558, ZN => n17555);
   U16255 : AOI22_X1 port map( A1 => n20872, A2 => n9000, B1 => n20866, B2 => 
                           n8616, ZN => n17558);
   U16256 : OAI221_X1 port map( B1 => n16276, B2 => n20884, C1 => n14283, C2 =>
                           n20878, A => n17540, ZN => n17537);
   U16257 : AOI22_X1 port map( A1 => n20872, A2 => n8996, B1 => n20866, B2 => 
                           n8612, ZN => n17540);
   U16258 : OAI221_X1 port map( B1 => n16257, B2 => n20884, C1 => n14282, C2 =>
                           n20878, A => n17522, ZN => n17519);
   U16259 : AOI22_X1 port map( A1 => n20872, A2 => n8992, B1 => n20866, B2 => 
                           n8608, ZN => n17522);
   U16260 : OAI221_X1 port map( B1 => n16238, B2 => n20884, C1 => n14281, C2 =>
                           n20878, A => n17504, ZN => n17501);
   U16261 : AOI22_X1 port map( A1 => n20872, A2 => n8988, B1 => n20866, B2 => 
                           n8604, ZN => n17504);
   U16262 : OAI221_X1 port map( B1 => n16219, B2 => n20884, C1 => n14280, C2 =>
                           n20878, A => n17486, ZN => n17483);
   U16263 : AOI22_X1 port map( A1 => n20872, A2 => n8984, B1 => n20866, B2 => 
                           n8600, ZN => n17486);
   U16264 : OAI221_X1 port map( B1 => n16200, B2 => n20884, C1 => n14279, C2 =>
                           n20878, A => n17468, ZN => n17465);
   U16265 : AOI22_X1 port map( A1 => n20872, A2 => n8980, B1 => n20866, B2 => 
                           n8596, ZN => n17468);
   U16266 : OAI221_X1 port map( B1 => n16181, B2 => n20884, C1 => n14278, C2 =>
                           n20878, A => n17450, ZN => n17447);
   U16267 : AOI22_X1 port map( A1 => n20872, A2 => n8976, B1 => n20866, B2 => 
                           n8592, ZN => n17450);
   U16268 : OAI221_X1 port map( B1 => n14597, B2 => n21077, C1 => n14929, C2 =>
                           n21067, A => n17139, ZN => n17136);
   U16269 : AOI22_X1 port map( A1 => n19624, A2 => n21086, B1 => n21084, B2 => 
                           n19625, ZN => n17139);
   U16270 : OAI221_X1 port map( B1 => n14596, B2 => n21077, C1 => n14928, C2 =>
                           n21067, A => n17120, ZN => n17117);
   U16271 : AOI22_X1 port map( A1 => n19604, A2 => n21086, B1 => n21084, B2 => 
                           n19605, ZN => n17120);
   U16272 : OAI221_X1 port map( B1 => n14595, B2 => n21077, C1 => n14927, C2 =>
                           n21067, A => n17101, ZN => n17098);
   U16273 : AOI22_X1 port map( A1 => n19584, A2 => n21086, B1 => n21084, B2 => 
                           n19585, ZN => n17101);
   U16274 : OAI221_X1 port map( B1 => n14594, B2 => n21077, C1 => n14926, C2 =>
                           n21068, A => n17082, ZN => n17079);
   U16275 : AOI22_X1 port map( A1 => n19564, A2 => n21087, B1 => n21084, B2 => 
                           n19565, ZN => n17082);
   U16276 : OAI221_X1 port map( B1 => n14593, B2 => n21077, C1 => n14925, C2 =>
                           n21068, A => n17063, ZN => n17060);
   U16277 : AOI22_X1 port map( A1 => n19544, A2 => n21087, B1 => n21084, B2 => 
                           n19545, ZN => n17063);
   U16278 : OAI221_X1 port map( B1 => n14592, B2 => n21077, C1 => n14924, C2 =>
                           n21068, A => n17044, ZN => n17041);
   U16279 : AOI22_X1 port map( A1 => n19524, A2 => n21087, B1 => n21084, B2 => 
                           n19525, ZN => n17044);
   U16280 : OAI221_X1 port map( B1 => n14591, B2 => n21077, C1 => n14923, C2 =>
                           n21068, A => n17025, ZN => n17022);
   U16281 : AOI22_X1 port map( A1 => n19504, A2 => n21087, B1 => n21084, B2 => 
                           n19505, ZN => n17025);
   U16282 : OAI221_X1 port map( B1 => n14590, B2 => n21076, C1 => n14922, C2 =>
                           n21068, A => n17006, ZN => n17003);
   U16283 : AOI22_X1 port map( A1 => n19484, A2 => n21087, B1 => n21084, B2 => 
                           n19485, ZN => n17006);
   U16284 : OAI221_X1 port map( B1 => n14589, B2 => n21076, C1 => n14921, C2 =>
                           n21068, A => n16987, ZN => n16984);
   U16285 : AOI22_X1 port map( A1 => n19464, A2 => n21087, B1 => n21084, B2 => 
                           n19465, ZN => n16987);
   U16286 : OAI221_X1 port map( B1 => n14588, B2 => n21076, C1 => n14920, C2 =>
                           n21068, A => n16968, ZN => n16965);
   U16287 : AOI22_X1 port map( A1 => n19444, A2 => n21087, B1 => n21084, B2 => 
                           n19445, ZN => n16968);
   U16288 : OAI221_X1 port map( B1 => n14587, B2 => n21076, C1 => n14919, C2 =>
                           n21068, A => n16949, ZN => n16946);
   U16289 : AOI22_X1 port map( A1 => n19424, A2 => n21087, B1 => n21084, B2 => 
                           n19425, ZN => n16949);
   U16290 : OAI221_X1 port map( B1 => n14586, B2 => n21076, C1 => n14918, C2 =>
                           n21068, A => n16930, ZN => n16927);
   U16291 : AOI22_X1 port map( A1 => n19404, A2 => n21087, B1 => n21084, B2 => 
                           n19405, ZN => n16930);
   U16292 : OAI221_X1 port map( B1 => n14585, B2 => n21076, C1 => n14917, C2 =>
                           n21068, A => n16911, ZN => n16908);
   U16293 : AOI22_X1 port map( A1 => n19384, A2 => n21087, B1 => n21084, B2 => 
                           n19385, ZN => n16911);
   U16294 : OAI221_X1 port map( B1 => n14584, B2 => n21076, C1 => n14916, C2 =>
                           n21068, A => n16892, ZN => n16889);
   U16295 : AOI22_X1 port map( A1 => n19364, A2 => n21087, B1 => n21084, B2 => 
                           n19365, ZN => n16892);
   U16296 : OAI221_X1 port map( B1 => n14583, B2 => n21076, C1 => n14915, C2 =>
                           n21068, A => n16873, ZN => n16870);
   U16297 : AOI22_X1 port map( A1 => n19344, A2 => n21087, B1 => n21083, B2 => 
                           n19345, ZN => n16873);
   U16298 : OAI221_X1 port map( B1 => n14582, B2 => n21076, C1 => n14914, C2 =>
                           n21069, A => n16854, ZN => n16851);
   U16299 : AOI22_X1 port map( A1 => n19324, A2 => n21088, B1 => n21083, B2 => 
                           n19325, ZN => n16854);
   U16300 : OAI221_X1 port map( B1 => n14581, B2 => n21076, C1 => n14913, C2 =>
                           n21069, A => n16835, ZN => n16832);
   U16301 : AOI22_X1 port map( A1 => n19304, A2 => n21088, B1 => n21083, B2 => 
                           n19305, ZN => n16835);
   U16302 : OAI221_X1 port map( B1 => n14580, B2 => n21076, C1 => n14912, C2 =>
                           n21069, A => n16816, ZN => n16813);
   U16303 : AOI22_X1 port map( A1 => n19284, A2 => n21088, B1 => n21083, B2 => 
                           n19285, ZN => n16816);
   U16304 : OAI221_X1 port map( B1 => n14579, B2 => n21076, C1 => n14911, C2 =>
                           n21069, A => n16797, ZN => n16794);
   U16305 : AOI22_X1 port map( A1 => n19264, A2 => n21088, B1 => n21083, B2 => 
                           n19265, ZN => n16797);
   U16306 : OAI221_X1 port map( B1 => n14578, B2 => n21075, C1 => n14910, C2 =>
                           n21069, A => n16778, ZN => n16775);
   U16307 : AOI22_X1 port map( A1 => n19244, A2 => n21088, B1 => n21083, B2 => 
                           n19245, ZN => n16778);
   U16308 : OAI221_X1 port map( B1 => n14577, B2 => n21075, C1 => n14909, C2 =>
                           n21069, A => n16759, ZN => n16756);
   U16309 : AOI22_X1 port map( A1 => n19224, A2 => n21088, B1 => n21083, B2 => 
                           n19225, ZN => n16759);
   U16310 : OAI221_X1 port map( B1 => n14576, B2 => n21075, C1 => n14908, C2 =>
                           n21069, A => n16740, ZN => n16737);
   U16311 : AOI22_X1 port map( A1 => n19204, A2 => n21088, B1 => n21083, B2 => 
                           n19205, ZN => n16740);
   U16312 : OAI221_X1 port map( B1 => n14575, B2 => n21075, C1 => n14907, C2 =>
                           n21069, A => n16721, ZN => n16718);
   U16313 : AOI22_X1 port map( A1 => n19184, A2 => n21088, B1 => n21083, B2 => 
                           n19185, ZN => n16721);
   U16314 : OAI221_X1 port map( B1 => n14574, B2 => n21075, C1 => n14906, C2 =>
                           n21069, A => n16702, ZN => n16699);
   U16315 : AOI22_X1 port map( A1 => n19164, A2 => n21088, B1 => n21083, B2 => 
                           n19165, ZN => n16702);
   U16316 : OAI221_X1 port map( B1 => n14573, B2 => n21075, C1 => n14905, C2 =>
                           n21069, A => n16683, ZN => n16680);
   U16317 : AOI22_X1 port map( A1 => n19144, A2 => n21088, B1 => n21083, B2 => 
                           n19145, ZN => n16683);
   U16318 : OAI221_X1 port map( B1 => n14572, B2 => n21075, C1 => n14904, C2 =>
                           n21069, A => n16664, ZN => n16661);
   U16319 : AOI22_X1 port map( A1 => n19124, A2 => n21088, B1 => n21083, B2 => 
                           n19125, ZN => n16664);
   U16320 : OAI221_X1 port map( B1 => n14571, B2 => n21075, C1 => n14903, C2 =>
                           n21069, A => n16645, ZN => n16642);
   U16321 : AOI22_X1 port map( A1 => n19104, A2 => n21088, B1 => n21083, B2 => 
                           n19105, ZN => n16645);
   U16322 : OAI221_X1 port map( B1 => n14570, B2 => n21075, C1 => n14902, C2 =>
                           n21070, A => n16626, ZN => n16623);
   U16323 : AOI22_X1 port map( A1 => n19084, A2 => n21089, B1 => n21083, B2 => 
                           n19085, ZN => n16626);
   U16324 : OAI221_X1 port map( B1 => n14569, B2 => n21075, C1 => n14901, C2 =>
                           n21070, A => n16607, ZN => n16604);
   U16325 : AOI22_X1 port map( A1 => n19064, A2 => n21089, B1 => n21082, B2 => 
                           n19065, ZN => n16607);
   U16326 : OAI221_X1 port map( B1 => n14568, B2 => n21075, C1 => n14900, C2 =>
                           n21070, A => n16588, ZN => n16585);
   U16327 : AOI22_X1 port map( A1 => n19044, A2 => n21089, B1 => n21082, B2 => 
                           n19045, ZN => n16588);
   U16328 : OAI221_X1 port map( B1 => n14567, B2 => n21075, C1 => n14899, C2 =>
                           n21070, A => n16569, ZN => n16566);
   U16329 : AOI22_X1 port map( A1 => n19024, A2 => n21089, B1 => n21082, B2 => 
                           n19025, ZN => n16569);
   U16330 : OAI221_X1 port map( B1 => n14566, B2 => n21074, C1 => n14898, C2 =>
                           n21070, A => n16550, ZN => n16547);
   U16331 : AOI22_X1 port map( A1 => n19004, A2 => n21089, B1 => n21082, B2 => 
                           n19005, ZN => n16550);
   U16332 : OAI221_X1 port map( B1 => n14565, B2 => n21074, C1 => n14897, C2 =>
                           n21070, A => n16531, ZN => n16528);
   U16333 : AOI22_X1 port map( A1 => n18984, A2 => n21089, B1 => n21082, B2 => 
                           n18985, ZN => n16531);
   U16334 : OAI221_X1 port map( B1 => n14564, B2 => n21074, C1 => n14896, C2 =>
                           n21070, A => n16512, ZN => n16509);
   U16335 : AOI22_X1 port map( A1 => n18964, A2 => n21089, B1 => n21082, B2 => 
                           n18965, ZN => n16512);
   U16336 : OAI221_X1 port map( B1 => n14563, B2 => n21074, C1 => n14895, C2 =>
                           n21070, A => n16493, ZN => n16490);
   U16337 : AOI22_X1 port map( A1 => n18944, A2 => n21089, B1 => n21082, B2 => 
                           n18945, ZN => n16493);
   U16338 : OAI221_X1 port map( B1 => n14562, B2 => n21074, C1 => n14894, C2 =>
                           n21070, A => n16474, ZN => n16471);
   U16339 : AOI22_X1 port map( A1 => n18924, A2 => n21089, B1 => n21082, B2 => 
                           n18925, ZN => n16474);
   U16340 : OAI221_X1 port map( B1 => n14561, B2 => n21074, C1 => n14893, C2 =>
                           n21070, A => n16455, ZN => n16452);
   U16341 : AOI22_X1 port map( A1 => n18904, A2 => n21089, B1 => n21082, B2 => 
                           n18905, ZN => n16455);
   U16342 : OAI221_X1 port map( B1 => n14560, B2 => n21074, C1 => n14892, C2 =>
                           n21070, A => n16436, ZN => n16433);
   U16343 : AOI22_X1 port map( A1 => n18884, A2 => n21089, B1 => n21082, B2 => 
                           n18885, ZN => n16436);
   U16344 : OAI221_X1 port map( B1 => n14559, B2 => n21074, C1 => n14891, C2 =>
                           n21070, A => n16417, ZN => n16414);
   U16345 : AOI22_X1 port map( A1 => n18864, A2 => n21089, B1 => n21082, B2 => 
                           n18865, ZN => n16417);
   U16346 : OAI221_X1 port map( B1 => n14558, B2 => n21074, C1 => n14890, C2 =>
                           n21071, A => n16398, ZN => n16395);
   U16347 : AOI22_X1 port map( A1 => n18844, A2 => n21090, B1 => n21082, B2 => 
                           n18845, ZN => n16398);
   U16348 : OAI221_X1 port map( B1 => n14557, B2 => n21074, C1 => n14889, C2 =>
                           n21071, A => n16379, ZN => n16376);
   U16349 : AOI22_X1 port map( A1 => n18824, A2 => n21090, B1 => n21082, B2 => 
                           n18825, ZN => n16379);
   U16350 : OAI221_X1 port map( B1 => n14556, B2 => n21074, C1 => n14888, C2 =>
                           n21071, A => n16360, ZN => n16357);
   U16351 : AOI22_X1 port map( A1 => n18804, A2 => n21090, B1 => n21082, B2 => 
                           n18805, ZN => n16360);
   U16352 : OAI221_X1 port map( B1 => n14555, B2 => n21074, C1 => n14887, C2 =>
                           n21071, A => n16341, ZN => n16338);
   U16353 : AOI22_X1 port map( A1 => n18784, A2 => n21090, B1 => n21081, B2 => 
                           n18785, ZN => n16341);
   U16354 : OAI221_X1 port map( B1 => n16162, B2 => n20885, C1 => n14277, C2 =>
                           n20879, A => n17432, ZN => n17429);
   U16355 : AOI22_X1 port map( A1 => n20873, A2 => n8972, B1 => n20867, B2 => 
                           n8588, ZN => n17432);
   U16356 : OAI221_X1 port map( B1 => n15744, B2 => n20789, C1 => n14746, C2 =>
                           n20783, A => n17440, ZN => n17437);
   U16357 : AOI22_X1 port map( A1 => n20777, A2 => n8835, B1 => n20771, B2 => 
                           n18619, ZN => n17440);
   U16358 : OAI221_X1 port map( B1 => n16143, B2 => n20885, C1 => n14276, C2 =>
                           n20879, A => n17414, ZN => n17411);
   U16359 : AOI22_X1 port map( A1 => n20873, A2 => n8968, B1 => n20867, B2 => 
                           n8584, ZN => n17414);
   U16360 : OAI221_X1 port map( B1 => n15743, B2 => n20789, C1 => n14745, C2 =>
                           n20783, A => n17422, ZN => n17419);
   U16361 : AOI22_X1 port map( A1 => n20777, A2 => n8833, B1 => n20771, B2 => 
                           n18599, ZN => n17422);
   U16362 : OAI221_X1 port map( B1 => n16124, B2 => n20885, C1 => n14275, C2 =>
                           n20879, A => n17396, ZN => n17393);
   U16363 : AOI22_X1 port map( A1 => n20873, A2 => n8964, B1 => n20867, B2 => 
                           n8580, ZN => n17396);
   U16364 : OAI221_X1 port map( B1 => n15742, B2 => n20789, C1 => n14744, C2 =>
                           n20783, A => n17404, ZN => n17401);
   U16365 : AOI22_X1 port map( A1 => n20777, A2 => n8831, B1 => n20771, B2 => 
                           n18579, ZN => n17404);
   U16366 : OAI221_X1 port map( B1 => n16070, B2 => n20885, C1 => n14273, C2 =>
                           n20879, A => n17352, ZN => n17343);
   U16367 : AOI22_X1 port map( A1 => n20873, A2 => n8960, B1 => n20867, B2 => 
                           n8576, ZN => n17352);
   U16368 : OAI221_X1 port map( B1 => n15740, B2 => n20789, C1 => n14742, C2 =>
                           n20783, A => n17376, ZN => n17368);
   U16369 : AOI22_X1 port map( A1 => n20777, A2 => n8829, B1 => n20771, B2 => 
                           n18559, ZN => n17376);
   U16370 : OAI221_X1 port map( B1 => n14606, B2 => n21078, C1 => n14938, C2 =>
                           n21067, A => n17317, ZN => n17308);
   U16371 : AOI22_X1 port map( A1 => n19804, A2 => n21086, B1 => n21085, B2 => 
                           n19805, ZN => n17317);
   U16372 : OAI221_X1 port map( B1 => n14605, B2 => n21078, C1 => n14937, C2 =>
                           n21067, A => n17291, ZN => n17288);
   U16373 : AOI22_X1 port map( A1 => n19784, A2 => n21086, B1 => n21085, B2 => 
                           n19785, ZN => n17291);
   U16374 : OAI221_X1 port map( B1 => n14604, B2 => n21078, C1 => n14936, C2 =>
                           n21067, A => n17272, ZN => n17269);
   U16375 : AOI22_X1 port map( A1 => n19764, A2 => n21086, B1 => n21085, B2 => 
                           n19765, ZN => n17272);
   U16376 : OAI221_X1 port map( B1 => n14603, B2 => n21078, C1 => n14935, C2 =>
                           n21067, A => n17253, ZN => n17250);
   U16377 : AOI22_X1 port map( A1 => n19744, A2 => n21086, B1 => n21085, B2 => 
                           n19745, ZN => n17253);
   U16378 : OAI221_X1 port map( B1 => n15744, B2 => n20981, C1 => n14746, C2 =>
                           n20975, A => n16178, ZN => n16175);
   U16379 : AOI22_X1 port map( A1 => n20969, A2 => n8835, B1 => n20963, B2 => 
                           n18619, ZN => n16178);
   U16380 : OAI221_X1 port map( B1 => n15743, B2 => n20981, C1 => n14745, C2 =>
                           n20975, A => n16159, ZN => n16156);
   U16381 : AOI22_X1 port map( A1 => n20969, A2 => n8833, B1 => n20963, B2 => 
                           n18599, ZN => n16159);
   U16382 : OAI221_X1 port map( B1 => n15742, B2 => n20981, C1 => n14744, C2 =>
                           n20975, A => n16140, ZN => n16137);
   U16383 : AOI22_X1 port map( A1 => n20969, A2 => n8831, B1 => n20963, B2 => 
                           n18579, ZN => n16140);
   U16384 : OAI221_X1 port map( B1 => n15740, B2 => n20981, C1 => n14742, C2 =>
                           n20975, A => n16111, ZN => n16102);
   U16385 : AOI22_X1 port map( A1 => n20969, A2 => n8829, B1 => n20963, B2 => 
                           n18559, ZN => n16111);
   U16386 : OAI221_X1 port map( B1 => n15457, B2 => n20857, C1 => n16056, C2 =>
                           n20851, A => n18297, ZN => n18292);
   U16387 : AOI22_X1 port map( A1 => n20845, A2 => n9163, B1 => n20839, B2 => 
                           n8779, ZN => n18297);
   U16388 : OAI221_X1 port map( B1 => n14259, B2 => n20761, C1 => n15325, C2 =>
                           n20755, A => n18305, ZN => n18300);
   U16389 : AOI22_X1 port map( A1 => n20749, A2 => n19574, B1 => n20743, B2 => 
                           n19575, ZN => n18305);
   U16390 : OAI221_X1 port map( B1 => n15456, B2 => n20857, C1 => n16055, C2 =>
                           n20851, A => n18279, ZN => n18274);
   U16391 : AOI22_X1 port map( A1 => n20845, A2 => n9159, B1 => n20839, B2 => 
                           n8775, ZN => n18279);
   U16392 : OAI221_X1 port map( B1 => n14258, B2 => n20761, C1 => n15324, C2 =>
                           n20755, A => n18287, ZN => n18282);
   U16393 : AOI22_X1 port map( A1 => n20749, A2 => n19554, B1 => n20743, B2 => 
                           n19555, ZN => n18287);
   U16394 : OAI221_X1 port map( B1 => n15455, B2 => n20857, C1 => n16054, C2 =>
                           n20851, A => n18261, ZN => n18256);
   U16395 : AOI22_X1 port map( A1 => n20845, A2 => n9155, B1 => n20839, B2 => 
                           n8771, ZN => n18261);
   U16396 : OAI221_X1 port map( B1 => n14257, B2 => n20761, C1 => n15323, C2 =>
                           n20755, A => n18269, ZN => n18264);
   U16397 : AOI22_X1 port map( A1 => n20749, A2 => n19534, B1 => n20743, B2 => 
                           n19535, ZN => n18269);
   U16398 : OAI221_X1 port map( B1 => n15454, B2 => n20857, C1 => n16053, C2 =>
                           n20851, A => n18243, ZN => n18238);
   U16399 : AOI22_X1 port map( A1 => n20845, A2 => n9151, B1 => n20839, B2 => 
                           n8767, ZN => n18243);
   U16400 : OAI221_X1 port map( B1 => n14256, B2 => n20761, C1 => n15322, C2 =>
                           n20755, A => n18251, ZN => n18246);
   U16401 : AOI22_X1 port map( A1 => n20749, A2 => n19514, B1 => n20743, B2 => 
                           n19515, ZN => n18251);
   U16402 : OAI221_X1 port map( B1 => n15453, B2 => n20857, C1 => n16052, C2 =>
                           n20851, A => n18225, ZN => n18220);
   U16403 : AOI22_X1 port map( A1 => n20845, A2 => n9147, B1 => n20839, B2 => 
                           n8763, ZN => n18225);
   U16404 : OAI221_X1 port map( B1 => n14255, B2 => n20761, C1 => n15321, C2 =>
                           n20755, A => n18233, ZN => n18228);
   U16405 : AOI22_X1 port map( A1 => n20749, A2 => n19494, B1 => n20743, B2 => 
                           n19495, ZN => n18233);
   U16406 : OAI221_X1 port map( B1 => n15452, B2 => n20857, C1 => n16051, C2 =>
                           n20851, A => n18207, ZN => n18202);
   U16407 : AOI22_X1 port map( A1 => n20845, A2 => n9143, B1 => n20839, B2 => 
                           n8759, ZN => n18207);
   U16408 : OAI221_X1 port map( B1 => n14254, B2 => n20761, C1 => n15320, C2 =>
                           n20755, A => n18215, ZN => n18210);
   U16409 : AOI22_X1 port map( A1 => n20749, A2 => n19474, B1 => n20743, B2 => 
                           n19475, ZN => n18215);
   U16410 : OAI221_X1 port map( B1 => n15451, B2 => n20857, C1 => n16050, C2 =>
                           n20851, A => n18189, ZN => n18184);
   U16411 : AOI22_X1 port map( A1 => n20845, A2 => n9139, B1 => n20839, B2 => 
                           n8755, ZN => n18189);
   U16412 : OAI221_X1 port map( B1 => n14253, B2 => n20761, C1 => n15319, C2 =>
                           n20755, A => n18197, ZN => n18192);
   U16413 : AOI22_X1 port map( A1 => n20749, A2 => n19454, B1 => n20743, B2 => 
                           n19455, ZN => n18197);
   U16414 : OAI221_X1 port map( B1 => n15450, B2 => n20857, C1 => n16049, C2 =>
                           n20851, A => n18171, ZN => n18166);
   U16415 : AOI22_X1 port map( A1 => n20845, A2 => n9135, B1 => n20839, B2 => 
                           n8751, ZN => n18171);
   U16416 : OAI221_X1 port map( B1 => n14252, B2 => n20761, C1 => n15318, C2 =>
                           n20755, A => n18179, ZN => n18174);
   U16417 : AOI22_X1 port map( A1 => n20749, A2 => n19434, B1 => n20743, B2 => 
                           n19435, ZN => n18179);
   U16418 : OAI221_X1 port map( B1 => n15449, B2 => n20857, C1 => n16048, C2 =>
                           n20851, A => n18153, ZN => n18148);
   U16419 : AOI22_X1 port map( A1 => n20845, A2 => n9131, B1 => n20839, B2 => 
                           n8747, ZN => n18153);
   U16420 : OAI221_X1 port map( B1 => n14251, B2 => n20761, C1 => n15317, C2 =>
                           n20755, A => n18161, ZN => n18156);
   U16421 : AOI22_X1 port map( A1 => n20749, A2 => n19414, B1 => n20743, B2 => 
                           n19415, ZN => n18161);
   U16422 : OAI221_X1 port map( B1 => n15448, B2 => n20857, C1 => n16047, C2 =>
                           n20851, A => n18135, ZN => n18130);
   U16423 : AOI22_X1 port map( A1 => n20845, A2 => n9127, B1 => n20839, B2 => 
                           n8743, ZN => n18135);
   U16424 : OAI221_X1 port map( B1 => n14250, B2 => n20761, C1 => n15316, C2 =>
                           n20755, A => n18143, ZN => n18138);
   U16425 : AOI22_X1 port map( A1 => n20749, A2 => n19394, B1 => n20743, B2 => 
                           n19395, ZN => n18143);
   U16426 : OAI221_X1 port map( B1 => n15447, B2 => n20857, C1 => n16046, C2 =>
                           n20851, A => n18117, ZN => n18112);
   U16427 : AOI22_X1 port map( A1 => n20845, A2 => n9123, B1 => n20839, B2 => 
                           n8739, ZN => n18117);
   U16428 : OAI221_X1 port map( B1 => n14249, B2 => n20761, C1 => n15315, C2 =>
                           n20755, A => n18125, ZN => n18120);
   U16429 : AOI22_X1 port map( A1 => n20749, A2 => n19374, B1 => n20743, B2 => 
                           n19375, ZN => n18125);
   U16430 : OAI221_X1 port map( B1 => n15446, B2 => n20857, C1 => n16045, C2 =>
                           n20851, A => n18099, ZN => n18094);
   U16431 : AOI22_X1 port map( A1 => n20845, A2 => n9119, B1 => n20839, B2 => 
                           n8735, ZN => n18099);
   U16432 : OAI221_X1 port map( B1 => n14248, B2 => n20761, C1 => n15314, C2 =>
                           n20755, A => n18107, ZN => n18102);
   U16433 : AOI22_X1 port map( A1 => n20749, A2 => n19354, B1 => n20743, B2 => 
                           n19355, ZN => n18107);
   U16434 : OAI221_X1 port map( B1 => n15445, B2 => n20858, C1 => n16044, C2 =>
                           n20852, A => n18081, ZN => n18076);
   U16435 : AOI22_X1 port map( A1 => n20846, A2 => n9115, B1 => n20840, B2 => 
                           n8731, ZN => n18081);
   U16436 : OAI221_X1 port map( B1 => n14247, B2 => n20762, C1 => n15313, C2 =>
                           n20756, A => n18089, ZN => n18084);
   U16437 : AOI22_X1 port map( A1 => n20750, A2 => n19334, B1 => n20744, B2 => 
                           n19335, ZN => n18089);
   U16438 : OAI221_X1 port map( B1 => n15444, B2 => n20858, C1 => n16043, C2 =>
                           n20852, A => n18063, ZN => n18058);
   U16439 : AOI22_X1 port map( A1 => n20846, A2 => n9111, B1 => n20840, B2 => 
                           n8727, ZN => n18063);
   U16440 : OAI221_X1 port map( B1 => n14246, B2 => n20762, C1 => n15312, C2 =>
                           n20756, A => n18071, ZN => n18066);
   U16441 : AOI22_X1 port map( A1 => n20750, A2 => n19314, B1 => n20744, B2 => 
                           n19315, ZN => n18071);
   U16442 : OAI221_X1 port map( B1 => n15443, B2 => n20858, C1 => n16042, C2 =>
                           n20852, A => n18045, ZN => n18040);
   U16443 : AOI22_X1 port map( A1 => n20846, A2 => n9107, B1 => n20840, B2 => 
                           n8723, ZN => n18045);
   U16444 : OAI221_X1 port map( B1 => n14245, B2 => n20762, C1 => n15311, C2 =>
                           n20756, A => n18053, ZN => n18048);
   U16445 : AOI22_X1 port map( A1 => n20750, A2 => n19294, B1 => n20744, B2 => 
                           n19295, ZN => n18053);
   U16446 : OAI221_X1 port map( B1 => n15442, B2 => n20858, C1 => n16041, C2 =>
                           n20852, A => n18027, ZN => n18022);
   U16447 : AOI22_X1 port map( A1 => n20846, A2 => n9103, B1 => n20840, B2 => 
                           n8719, ZN => n18027);
   U16448 : OAI221_X1 port map( B1 => n14244, B2 => n20762, C1 => n15310, C2 =>
                           n20756, A => n18035, ZN => n18030);
   U16449 : AOI22_X1 port map( A1 => n20750, A2 => n19274, B1 => n20744, B2 => 
                           n19275, ZN => n18035);
   U16450 : OAI221_X1 port map( B1 => n15441, B2 => n20858, C1 => n16040, C2 =>
                           n20852, A => n18009, ZN => n18004);
   U16451 : AOI22_X1 port map( A1 => n20846, A2 => n9099, B1 => n20840, B2 => 
                           n8715, ZN => n18009);
   U16452 : OAI221_X1 port map( B1 => n14243, B2 => n20762, C1 => n15309, C2 =>
                           n20756, A => n18017, ZN => n18012);
   U16453 : AOI22_X1 port map( A1 => n20750, A2 => n19254, B1 => n20744, B2 => 
                           n19255, ZN => n18017);
   U16454 : OAI221_X1 port map( B1 => n15440, B2 => n20858, C1 => n16039, C2 =>
                           n20852, A => n17991, ZN => n17986);
   U16455 : AOI22_X1 port map( A1 => n20846, A2 => n9095, B1 => n20840, B2 => 
                           n8711, ZN => n17991);
   U16456 : OAI221_X1 port map( B1 => n14242, B2 => n20762, C1 => n15308, C2 =>
                           n20756, A => n17999, ZN => n17994);
   U16457 : AOI22_X1 port map( A1 => n20750, A2 => n19234, B1 => n20744, B2 => 
                           n19235, ZN => n17999);
   U16458 : OAI221_X1 port map( B1 => n15439, B2 => n20858, C1 => n16038, C2 =>
                           n20852, A => n17973, ZN => n17968);
   U16459 : AOI22_X1 port map( A1 => n20846, A2 => n9091, B1 => n20840, B2 => 
                           n8707, ZN => n17973);
   U16460 : OAI221_X1 port map( B1 => n14241, B2 => n20762, C1 => n15307, C2 =>
                           n20756, A => n17981, ZN => n17976);
   U16461 : AOI22_X1 port map( A1 => n20750, A2 => n19214, B1 => n20744, B2 => 
                           n19215, ZN => n17981);
   U16462 : OAI221_X1 port map( B1 => n15438, B2 => n20858, C1 => n16037, C2 =>
                           n20852, A => n17955, ZN => n17950);
   U16463 : AOI22_X1 port map( A1 => n20846, A2 => n9087, B1 => n20840, B2 => 
                           n8703, ZN => n17955);
   U16464 : OAI221_X1 port map( B1 => n14240, B2 => n20762, C1 => n15306, C2 =>
                           n20756, A => n17963, ZN => n17958);
   U16465 : AOI22_X1 port map( A1 => n20750, A2 => n19194, B1 => n20744, B2 => 
                           n19195, ZN => n17963);
   U16466 : OAI221_X1 port map( B1 => n15437, B2 => n20858, C1 => n16036, C2 =>
                           n20852, A => n17937, ZN => n17932);
   U16467 : AOI22_X1 port map( A1 => n20846, A2 => n9083, B1 => n20840, B2 => 
                           n8699, ZN => n17937);
   U16468 : OAI221_X1 port map( B1 => n14239, B2 => n20762, C1 => n15305, C2 =>
                           n20756, A => n17945, ZN => n17940);
   U16469 : AOI22_X1 port map( A1 => n20750, A2 => n19174, B1 => n20744, B2 => 
                           n19175, ZN => n17945);
   U16470 : OAI221_X1 port map( B1 => n15436, B2 => n20858, C1 => n16035, C2 =>
                           n20852, A => n17919, ZN => n17914);
   U16471 : AOI22_X1 port map( A1 => n20846, A2 => n9079, B1 => n20840, B2 => 
                           n8695, ZN => n17919);
   U16472 : OAI221_X1 port map( B1 => n14238, B2 => n20762, C1 => n15304, C2 =>
                           n20756, A => n17927, ZN => n17922);
   U16473 : AOI22_X1 port map( A1 => n20750, A2 => n19154, B1 => n20744, B2 => 
                           n19155, ZN => n17927);
   U16474 : OAI221_X1 port map( B1 => n15435, B2 => n20858, C1 => n16034, C2 =>
                           n20852, A => n17901, ZN => n17896);
   U16475 : AOI22_X1 port map( A1 => n20846, A2 => n9075, B1 => n20840, B2 => 
                           n8691, ZN => n17901);
   U16476 : OAI221_X1 port map( B1 => n14237, B2 => n20762, C1 => n15303, C2 =>
                           n20756, A => n17909, ZN => n17904);
   U16477 : AOI22_X1 port map( A1 => n20750, A2 => n19134, B1 => n20744, B2 => 
                           n19135, ZN => n17909);
   U16478 : OAI221_X1 port map( B1 => n15434, B2 => n20858, C1 => n16033, C2 =>
                           n20852, A => n17883, ZN => n17878);
   U16479 : AOI22_X1 port map( A1 => n20846, A2 => n9071, B1 => n20840, B2 => 
                           n8687, ZN => n17883);
   U16480 : OAI221_X1 port map( B1 => n14236, B2 => n20762, C1 => n15302, C2 =>
                           n20756, A => n17891, ZN => n17886);
   U16481 : AOI22_X1 port map( A1 => n20750, A2 => n19114, B1 => n20744, B2 => 
                           n19115, ZN => n17891);
   U16482 : OAI221_X1 port map( B1 => n15433, B2 => n20859, C1 => n16032, C2 =>
                           n20853, A => n17865, ZN => n17860);
   U16483 : AOI22_X1 port map( A1 => n20847, A2 => n9067, B1 => n20841, B2 => 
                           n8683, ZN => n17865);
   U16484 : OAI221_X1 port map( B1 => n14235, B2 => n20763, C1 => n15301, C2 =>
                           n20757, A => n17873, ZN => n17868);
   U16485 : AOI22_X1 port map( A1 => n20751, A2 => n19094, B1 => n20745, B2 => 
                           n19095, ZN => n17873);
   U16486 : OAI221_X1 port map( B1 => n15432, B2 => n20859, C1 => n16031, C2 =>
                           n20853, A => n17847, ZN => n17842);
   U16487 : AOI22_X1 port map( A1 => n20847, A2 => n9063, B1 => n20841, B2 => 
                           n8679, ZN => n17847);
   U16488 : OAI221_X1 port map( B1 => n14234, B2 => n20763, C1 => n15300, C2 =>
                           n20757, A => n17855, ZN => n17850);
   U16489 : AOI22_X1 port map( A1 => n20751, A2 => n19074, B1 => n20745, B2 => 
                           n19075, ZN => n17855);
   U16490 : OAI221_X1 port map( B1 => n15431, B2 => n20859, C1 => n16030, C2 =>
                           n20853, A => n17829, ZN => n17824);
   U16491 : AOI22_X1 port map( A1 => n20847, A2 => n9059, B1 => n20841, B2 => 
                           n8675, ZN => n17829);
   U16492 : OAI221_X1 port map( B1 => n14233, B2 => n20763, C1 => n15299, C2 =>
                           n20757, A => n17837, ZN => n17832);
   U16493 : AOI22_X1 port map( A1 => n20751, A2 => n19054, B1 => n20745, B2 => 
                           n19055, ZN => n17837);
   U16494 : OAI221_X1 port map( B1 => n15430, B2 => n20859, C1 => n16029, C2 =>
                           n20853, A => n17811, ZN => n17806);
   U16495 : AOI22_X1 port map( A1 => n20847, A2 => n9055, B1 => n20841, B2 => 
                           n8671, ZN => n17811);
   U16496 : OAI221_X1 port map( B1 => n14232, B2 => n20763, C1 => n15298, C2 =>
                           n20757, A => n17819, ZN => n17814);
   U16497 : AOI22_X1 port map( A1 => n20751, A2 => n19034, B1 => n20745, B2 => 
                           n19035, ZN => n17819);
   U16498 : OAI221_X1 port map( B1 => n15429, B2 => n20859, C1 => n16028, C2 =>
                           n20853, A => n17793, ZN => n17788);
   U16499 : AOI22_X1 port map( A1 => n20847, A2 => n9051, B1 => n20841, B2 => 
                           n8667, ZN => n17793);
   U16500 : OAI221_X1 port map( B1 => n14231, B2 => n20763, C1 => n15297, C2 =>
                           n20757, A => n17801, ZN => n17796);
   U16501 : AOI22_X1 port map( A1 => n20751, A2 => n19014, B1 => n20745, B2 => 
                           n19015, ZN => n17801);
   U16502 : OAI221_X1 port map( B1 => n15428, B2 => n20859, C1 => n16027, C2 =>
                           n20853, A => n17775, ZN => n17770);
   U16503 : AOI22_X1 port map( A1 => n20847, A2 => n9047, B1 => n20841, B2 => 
                           n8663, ZN => n17775);
   U16504 : OAI221_X1 port map( B1 => n14230, B2 => n20763, C1 => n15296, C2 =>
                           n20757, A => n17783, ZN => n17778);
   U16505 : AOI22_X1 port map( A1 => n20751, A2 => n18994, B1 => n20745, B2 => 
                           n18995, ZN => n17783);
   U16506 : OAI221_X1 port map( B1 => n15427, B2 => n20859, C1 => n16026, C2 =>
                           n20853, A => n17757, ZN => n17752);
   U16507 : AOI22_X1 port map( A1 => n20847, A2 => n9043, B1 => n20841, B2 => 
                           n8659, ZN => n17757);
   U16508 : OAI221_X1 port map( B1 => n14229, B2 => n20763, C1 => n15295, C2 =>
                           n20757, A => n17765, ZN => n17760);
   U16509 : AOI22_X1 port map( A1 => n20751, A2 => n18974, B1 => n20745, B2 => 
                           n18975, ZN => n17765);
   U16510 : OAI221_X1 port map( B1 => n15426, B2 => n20859, C1 => n16025, C2 =>
                           n20853, A => n17739, ZN => n17734);
   U16511 : AOI22_X1 port map( A1 => n20847, A2 => n9039, B1 => n20841, B2 => 
                           n8655, ZN => n17739);
   U16512 : OAI221_X1 port map( B1 => n14228, B2 => n20763, C1 => n15294, C2 =>
                           n20757, A => n17747, ZN => n17742);
   U16513 : AOI22_X1 port map( A1 => n20751, A2 => n18954, B1 => n20745, B2 => 
                           n18955, ZN => n17747);
   U16514 : OAI221_X1 port map( B1 => n15425, B2 => n20859, C1 => n16024, C2 =>
                           n20853, A => n17721, ZN => n17716);
   U16515 : AOI22_X1 port map( A1 => n20847, A2 => n9035, B1 => n20841, B2 => 
                           n8651, ZN => n17721);
   U16516 : OAI221_X1 port map( B1 => n14227, B2 => n20763, C1 => n15293, C2 =>
                           n20757, A => n17729, ZN => n17724);
   U16517 : AOI22_X1 port map( A1 => n20751, A2 => n18934, B1 => n20745, B2 => 
                           n18935, ZN => n17729);
   U16518 : OAI221_X1 port map( B1 => n15424, B2 => n20859, C1 => n16023, C2 =>
                           n20853, A => n17703, ZN => n17698);
   U16519 : AOI22_X1 port map( A1 => n20847, A2 => n9031, B1 => n20841, B2 => 
                           n8647, ZN => n17703);
   U16520 : OAI221_X1 port map( B1 => n14226, B2 => n20763, C1 => n15292, C2 =>
                           n20757, A => n17711, ZN => n17706);
   U16521 : AOI22_X1 port map( A1 => n20751, A2 => n18914, B1 => n20745, B2 => 
                           n18915, ZN => n17711);
   U16522 : OAI221_X1 port map( B1 => n15423, B2 => n20859, C1 => n16022, C2 =>
                           n20853, A => n17685, ZN => n17680);
   U16523 : AOI22_X1 port map( A1 => n20847, A2 => n9027, B1 => n20841, B2 => 
                           n8643, ZN => n17685);
   U16524 : OAI221_X1 port map( B1 => n14225, B2 => n20763, C1 => n15291, C2 =>
                           n20757, A => n17693, ZN => n17688);
   U16525 : AOI22_X1 port map( A1 => n20751, A2 => n18894, B1 => n20745, B2 => 
                           n18895, ZN => n17693);
   U16526 : OAI221_X1 port map( B1 => n15422, B2 => n20859, C1 => n16021, C2 =>
                           n20853, A => n17667, ZN => n17662);
   U16527 : AOI22_X1 port map( A1 => n20847, A2 => n9023, B1 => n20841, B2 => 
                           n8639, ZN => n17667);
   U16528 : OAI221_X1 port map( B1 => n14224, B2 => n20763, C1 => n15290, C2 =>
                           n20757, A => n17675, ZN => n17670);
   U16529 : AOI22_X1 port map( A1 => n20751, A2 => n18874, B1 => n20745, B2 => 
                           n18875, ZN => n17675);
   U16530 : OAI221_X1 port map( B1 => n15421, B2 => n20860, C1 => n16020, C2 =>
                           n20854, A => n17649, ZN => n17644);
   U16531 : AOI22_X1 port map( A1 => n20848, A2 => n9019, B1 => n20842, B2 => 
                           n8635, ZN => n17649);
   U16532 : OAI221_X1 port map( B1 => n14223, B2 => n20764, C1 => n15289, C2 =>
                           n20758, A => n17657, ZN => n17652);
   U16533 : AOI22_X1 port map( A1 => n20752, A2 => n18854, B1 => n20746, B2 => 
                           n18855, ZN => n17657);
   U16534 : OAI221_X1 port map( B1 => n15420, B2 => n20860, C1 => n16019, C2 =>
                           n20854, A => n17631, ZN => n17626);
   U16535 : AOI22_X1 port map( A1 => n20848, A2 => n9015, B1 => n20842, B2 => 
                           n8631, ZN => n17631);
   U16536 : OAI221_X1 port map( B1 => n14222, B2 => n20764, C1 => n15288, C2 =>
                           n20758, A => n17639, ZN => n17634);
   U16537 : AOI22_X1 port map( A1 => n20752, A2 => n18834, B1 => n20746, B2 => 
                           n18835, ZN => n17639);
   U16538 : OAI221_X1 port map( B1 => n15419, B2 => n20860, C1 => n16018, C2 =>
                           n20854, A => n17613, ZN => n17608);
   U16539 : AOI22_X1 port map( A1 => n20848, A2 => n9011, B1 => n20842, B2 => 
                           n8627, ZN => n17613);
   U16540 : OAI221_X1 port map( B1 => n14221, B2 => n20764, C1 => n15287, C2 =>
                           n20758, A => n17621, ZN => n17616);
   U16541 : AOI22_X1 port map( A1 => n20752, A2 => n18814, B1 => n20746, B2 => 
                           n18815, ZN => n17621);
   U16542 : OAI221_X1 port map( B1 => n15418, B2 => n20860, C1 => n16017, C2 =>
                           n20854, A => n17595, ZN => n17590);
   U16543 : AOI22_X1 port map( A1 => n20848, A2 => n9007, B1 => n20842, B2 => 
                           n8623, ZN => n17595);
   U16544 : OAI221_X1 port map( B1 => n14220, B2 => n20764, C1 => n15286, C2 =>
                           n20758, A => n17603, ZN => n17598);
   U16545 : AOI22_X1 port map( A1 => n20752, A2 => n18794, B1 => n20746, B2 => 
                           n18795, ZN => n17603);
   U16546 : OAI221_X1 port map( B1 => n15417, B2 => n20860, C1 => n16016, C2 =>
                           n20854, A => n17577, ZN => n17572);
   U16547 : AOI22_X1 port map( A1 => n20848, A2 => n9003, B1 => n20842, B2 => 
                           n8619, ZN => n17577);
   U16548 : OAI221_X1 port map( B1 => n14219, B2 => n20764, C1 => n15285, C2 =>
                           n20758, A => n17585, ZN => n17580);
   U16549 : AOI22_X1 port map( A1 => n20752, A2 => n18774, B1 => n20746, B2 => 
                           n18775, ZN => n17585);
   U16550 : OAI221_X1 port map( B1 => n15416, B2 => n20860, C1 => n16015, C2 =>
                           n20854, A => n17559, ZN => n17554);
   U16551 : AOI22_X1 port map( A1 => n20848, A2 => n8999, B1 => n20842, B2 => 
                           n8615, ZN => n17559);
   U16552 : OAI221_X1 port map( B1 => n14218, B2 => n20764, C1 => n15284, C2 =>
                           n20758, A => n17567, ZN => n17562);
   U16553 : AOI22_X1 port map( A1 => n20752, A2 => n18754, B1 => n20746, B2 => 
                           n18755, ZN => n17567);
   U16554 : OAI221_X1 port map( B1 => n15415, B2 => n20860, C1 => n16014, C2 =>
                           n20854, A => n17541, ZN => n17536);
   U16555 : AOI22_X1 port map( A1 => n20848, A2 => n8995, B1 => n20842, B2 => 
                           n8611, ZN => n17541);
   U16556 : OAI221_X1 port map( B1 => n14217, B2 => n20764, C1 => n15283, C2 =>
                           n20758, A => n17549, ZN => n17544);
   U16557 : AOI22_X1 port map( A1 => n20752, A2 => n18734, B1 => n20746, B2 => 
                           n18735, ZN => n17549);
   U16558 : OAI221_X1 port map( B1 => n15414, B2 => n20860, C1 => n16013, C2 =>
                           n20854, A => n17523, ZN => n17518);
   U16559 : AOI22_X1 port map( A1 => n20848, A2 => n8991, B1 => n20842, B2 => 
                           n8607, ZN => n17523);
   U16560 : OAI221_X1 port map( B1 => n14216, B2 => n20764, C1 => n15282, C2 =>
                           n20758, A => n17531, ZN => n17526);
   U16561 : AOI22_X1 port map( A1 => n20752, A2 => n18714, B1 => n20746, B2 => 
                           n18715, ZN => n17531);
   U16562 : OAI221_X1 port map( B1 => n15413, B2 => n20860, C1 => n16012, C2 =>
                           n20854, A => n17505, ZN => n17500);
   U16563 : AOI22_X1 port map( A1 => n20848, A2 => n8987, B1 => n20842, B2 => 
                           n8603, ZN => n17505);
   U16564 : OAI221_X1 port map( B1 => n14215, B2 => n20764, C1 => n15281, C2 =>
                           n20758, A => n17513, ZN => n17508);
   U16565 : AOI22_X1 port map( A1 => n20752, A2 => n18694, B1 => n20746, B2 => 
                           n18695, ZN => n17513);
   U16566 : OAI221_X1 port map( B1 => n15412, B2 => n20860, C1 => n16011, C2 =>
                           n20854, A => n17487, ZN => n17482);
   U16567 : AOI22_X1 port map( A1 => n20848, A2 => n8983, B1 => n20842, B2 => 
                           n8599, ZN => n17487);
   U16568 : OAI221_X1 port map( B1 => n14214, B2 => n20764, C1 => n15280, C2 =>
                           n20758, A => n17495, ZN => n17490);
   U16569 : AOI22_X1 port map( A1 => n20752, A2 => n18674, B1 => n20746, B2 => 
                           n18675, ZN => n17495);
   U16570 : OAI221_X1 port map( B1 => n15411, B2 => n20860, C1 => n16010, C2 =>
                           n20854, A => n17469, ZN => n17464);
   U16571 : AOI22_X1 port map( A1 => n20848, A2 => n8979, B1 => n20842, B2 => 
                           n8595, ZN => n17469);
   U16572 : OAI221_X1 port map( B1 => n14213, B2 => n20764, C1 => n15279, C2 =>
                           n20758, A => n17477, ZN => n17472);
   U16573 : AOI22_X1 port map( A1 => n20752, A2 => n18654, B1 => n20746, B2 => 
                           n18655, ZN => n17477);
   U16574 : OAI221_X1 port map( B1 => n15410, B2 => n20860, C1 => n16009, C2 =>
                           n20854, A => n17451, ZN => n17446);
   U16575 : AOI22_X1 port map( A1 => n20848, A2 => n8975, B1 => n20842, B2 => 
                           n8591, ZN => n17451);
   U16576 : OAI221_X1 port map( B1 => n14212, B2 => n20764, C1 => n15278, C2 =>
                           n20758, A => n17459, ZN => n17454);
   U16577 : AOI22_X1 port map( A1 => n20752, A2 => n18634, B1 => n20746, B2 => 
                           n18635, ZN => n17459);
   U16578 : OAI221_X1 port map( B1 => n14259, B2 => n20953, C1 => n15325, C2 =>
                           n20947, A => n17091, ZN => n17086);
   U16579 : AOI22_X1 port map( A1 => n20941, A2 => n19574, B1 => n20935, B2 => 
                           n19575, ZN => n17091);
   U16580 : OAI221_X1 port map( B1 => n14258, B2 => n20953, C1 => n15324, C2 =>
                           n20947, A => n17072, ZN => n17067);
   U16581 : AOI22_X1 port map( A1 => n20941, A2 => n19554, B1 => n20935, B2 => 
                           n19555, ZN => n17072);
   U16582 : OAI221_X1 port map( B1 => n14257, B2 => n20953, C1 => n15323, C2 =>
                           n20947, A => n17053, ZN => n17048);
   U16583 : AOI22_X1 port map( A1 => n20941, A2 => n19534, B1 => n20935, B2 => 
                           n19535, ZN => n17053);
   U16584 : OAI221_X1 port map( B1 => n14256, B2 => n20953, C1 => n15322, C2 =>
                           n20947, A => n17034, ZN => n17029);
   U16585 : AOI22_X1 port map( A1 => n20941, A2 => n19514, B1 => n20935, B2 => 
                           n19515, ZN => n17034);
   U16586 : OAI221_X1 port map( B1 => n14255, B2 => n20953, C1 => n15321, C2 =>
                           n20947, A => n17015, ZN => n17010);
   U16587 : AOI22_X1 port map( A1 => n20941, A2 => n19494, B1 => n20935, B2 => 
                           n19495, ZN => n17015);
   U16588 : OAI221_X1 port map( B1 => n14254, B2 => n20953, C1 => n15320, C2 =>
                           n20947, A => n16996, ZN => n16991);
   U16589 : AOI22_X1 port map( A1 => n20941, A2 => n19474, B1 => n20935, B2 => 
                           n19475, ZN => n16996);
   U16590 : OAI221_X1 port map( B1 => n14253, B2 => n20953, C1 => n15319, C2 =>
                           n20947, A => n16977, ZN => n16972);
   U16591 : AOI22_X1 port map( A1 => n20941, A2 => n19454, B1 => n20935, B2 => 
                           n19455, ZN => n16977);
   U16592 : OAI221_X1 port map( B1 => n14252, B2 => n20953, C1 => n15318, C2 =>
                           n20947, A => n16958, ZN => n16953);
   U16593 : AOI22_X1 port map( A1 => n20941, A2 => n19434, B1 => n20935, B2 => 
                           n19435, ZN => n16958);
   U16594 : OAI221_X1 port map( B1 => n14251, B2 => n20953, C1 => n15317, C2 =>
                           n20947, A => n16939, ZN => n16934);
   U16595 : AOI22_X1 port map( A1 => n20941, A2 => n19414, B1 => n20935, B2 => 
                           n19415, ZN => n16939);
   U16596 : OAI221_X1 port map( B1 => n14250, B2 => n20953, C1 => n15316, C2 =>
                           n20947, A => n16920, ZN => n16915);
   U16597 : AOI22_X1 port map( A1 => n20941, A2 => n19394, B1 => n20935, B2 => 
                           n19395, ZN => n16920);
   U16598 : OAI221_X1 port map( B1 => n14249, B2 => n20953, C1 => n15315, C2 =>
                           n20947, A => n16901, ZN => n16896);
   U16599 : AOI22_X1 port map( A1 => n20941, A2 => n19374, B1 => n20935, B2 => 
                           n19375, ZN => n16901);
   U16600 : OAI221_X1 port map( B1 => n14248, B2 => n20953, C1 => n15314, C2 =>
                           n20947, A => n16882, ZN => n16877);
   U16601 : AOI22_X1 port map( A1 => n20941, A2 => n19354, B1 => n20935, B2 => 
                           n19355, ZN => n16882);
   U16602 : OAI221_X1 port map( B1 => n14247, B2 => n20954, C1 => n15313, C2 =>
                           n20948, A => n16863, ZN => n16858);
   U16603 : AOI22_X1 port map( A1 => n20942, A2 => n19334, B1 => n20936, B2 => 
                           n19335, ZN => n16863);
   U16604 : OAI221_X1 port map( B1 => n14246, B2 => n20954, C1 => n15312, C2 =>
                           n20948, A => n16844, ZN => n16839);
   U16605 : AOI22_X1 port map( A1 => n20942, A2 => n19314, B1 => n20936, B2 => 
                           n19315, ZN => n16844);
   U16606 : OAI221_X1 port map( B1 => n14245, B2 => n20954, C1 => n15311, C2 =>
                           n20948, A => n16825, ZN => n16820);
   U16607 : AOI22_X1 port map( A1 => n20942, A2 => n19294, B1 => n20936, B2 => 
                           n19295, ZN => n16825);
   U16608 : OAI221_X1 port map( B1 => n14244, B2 => n20954, C1 => n15310, C2 =>
                           n20948, A => n16806, ZN => n16801);
   U16609 : AOI22_X1 port map( A1 => n20942, A2 => n19274, B1 => n20936, B2 => 
                           n19275, ZN => n16806);
   U16610 : OAI221_X1 port map( B1 => n14243, B2 => n20954, C1 => n15309, C2 =>
                           n20948, A => n16787, ZN => n16782);
   U16611 : AOI22_X1 port map( A1 => n20942, A2 => n19254, B1 => n20936, B2 => 
                           n19255, ZN => n16787);
   U16612 : OAI221_X1 port map( B1 => n14242, B2 => n20954, C1 => n15308, C2 =>
                           n20948, A => n16768, ZN => n16763);
   U16613 : AOI22_X1 port map( A1 => n20942, A2 => n19234, B1 => n20936, B2 => 
                           n19235, ZN => n16768);
   U16614 : OAI221_X1 port map( B1 => n14241, B2 => n20954, C1 => n15307, C2 =>
                           n20948, A => n16749, ZN => n16744);
   U16615 : AOI22_X1 port map( A1 => n20942, A2 => n19214, B1 => n20936, B2 => 
                           n19215, ZN => n16749);
   U16616 : OAI221_X1 port map( B1 => n14240, B2 => n20954, C1 => n15306, C2 =>
                           n20948, A => n16730, ZN => n16725);
   U16617 : AOI22_X1 port map( A1 => n20942, A2 => n19194, B1 => n20936, B2 => 
                           n19195, ZN => n16730);
   U16618 : OAI221_X1 port map( B1 => n14239, B2 => n20954, C1 => n15305, C2 =>
                           n20948, A => n16711, ZN => n16706);
   U16619 : AOI22_X1 port map( A1 => n20942, A2 => n19174, B1 => n20936, B2 => 
                           n19175, ZN => n16711);
   U16620 : OAI221_X1 port map( B1 => n14238, B2 => n20954, C1 => n15304, C2 =>
                           n20948, A => n16692, ZN => n16687);
   U16621 : AOI22_X1 port map( A1 => n20942, A2 => n19154, B1 => n20936, B2 => 
                           n19155, ZN => n16692);
   U16622 : OAI221_X1 port map( B1 => n14237, B2 => n20954, C1 => n15303, C2 =>
                           n20948, A => n16673, ZN => n16668);
   U16623 : AOI22_X1 port map( A1 => n20942, A2 => n19134, B1 => n20936, B2 => 
                           n19135, ZN => n16673);
   U16624 : OAI221_X1 port map( B1 => n14236, B2 => n20954, C1 => n15302, C2 =>
                           n20948, A => n16654, ZN => n16649);
   U16625 : AOI22_X1 port map( A1 => n20942, A2 => n19114, B1 => n20936, B2 => 
                           n19115, ZN => n16654);
   U16626 : OAI221_X1 port map( B1 => n14235, B2 => n20955, C1 => n15301, C2 =>
                           n20949, A => n16635, ZN => n16630);
   U16627 : AOI22_X1 port map( A1 => n20943, A2 => n19094, B1 => n20937, B2 => 
                           n19095, ZN => n16635);
   U16628 : OAI221_X1 port map( B1 => n14234, B2 => n20955, C1 => n15300, C2 =>
                           n20949, A => n16616, ZN => n16611);
   U16629 : AOI22_X1 port map( A1 => n20943, A2 => n19074, B1 => n20937, B2 => 
                           n19075, ZN => n16616);
   U16630 : OAI221_X1 port map( B1 => n14233, B2 => n20955, C1 => n15299, C2 =>
                           n20949, A => n16597, ZN => n16592);
   U16631 : AOI22_X1 port map( A1 => n20943, A2 => n19054, B1 => n20937, B2 => 
                           n19055, ZN => n16597);
   U16632 : OAI221_X1 port map( B1 => n14232, B2 => n20955, C1 => n15298, C2 =>
                           n20949, A => n16578, ZN => n16573);
   U16633 : AOI22_X1 port map( A1 => n20943, A2 => n19034, B1 => n20937, B2 => 
                           n19035, ZN => n16578);
   U16634 : OAI221_X1 port map( B1 => n14231, B2 => n20955, C1 => n15297, C2 =>
                           n20949, A => n16559, ZN => n16554);
   U16635 : AOI22_X1 port map( A1 => n20943, A2 => n19014, B1 => n20937, B2 => 
                           n19015, ZN => n16559);
   U16636 : OAI221_X1 port map( B1 => n14230, B2 => n20955, C1 => n15296, C2 =>
                           n20949, A => n16540, ZN => n16535);
   U16637 : AOI22_X1 port map( A1 => n20943, A2 => n18994, B1 => n20937, B2 => 
                           n18995, ZN => n16540);
   U16638 : OAI221_X1 port map( B1 => n14229, B2 => n20955, C1 => n15295, C2 =>
                           n20949, A => n16521, ZN => n16516);
   U16639 : AOI22_X1 port map( A1 => n20943, A2 => n18974, B1 => n20937, B2 => 
                           n18975, ZN => n16521);
   U16640 : OAI221_X1 port map( B1 => n14228, B2 => n20955, C1 => n15294, C2 =>
                           n20949, A => n16502, ZN => n16497);
   U16641 : AOI22_X1 port map( A1 => n20943, A2 => n18954, B1 => n20937, B2 => 
                           n18955, ZN => n16502);
   U16642 : OAI221_X1 port map( B1 => n14227, B2 => n20955, C1 => n15293, C2 =>
                           n20949, A => n16483, ZN => n16478);
   U16643 : AOI22_X1 port map( A1 => n20943, A2 => n18934, B1 => n20937, B2 => 
                           n18935, ZN => n16483);
   U16644 : OAI221_X1 port map( B1 => n14226, B2 => n20955, C1 => n15292, C2 =>
                           n20949, A => n16464, ZN => n16459);
   U16645 : AOI22_X1 port map( A1 => n20943, A2 => n18914, B1 => n20937, B2 => 
                           n18915, ZN => n16464);
   U16646 : OAI221_X1 port map( B1 => n14225, B2 => n20955, C1 => n15291, C2 =>
                           n20949, A => n16445, ZN => n16440);
   U16647 : AOI22_X1 port map( A1 => n20943, A2 => n18894, B1 => n20937, B2 => 
                           n18895, ZN => n16445);
   U16648 : OAI221_X1 port map( B1 => n14224, B2 => n20955, C1 => n15290, C2 =>
                           n20949, A => n16426, ZN => n16421);
   U16649 : AOI22_X1 port map( A1 => n20943, A2 => n18874, B1 => n20937, B2 => 
                           n18875, ZN => n16426);
   U16650 : OAI221_X1 port map( B1 => n14223, B2 => n20956, C1 => n15289, C2 =>
                           n20950, A => n16407, ZN => n16402);
   U16651 : AOI22_X1 port map( A1 => n20944, A2 => n18854, B1 => n20938, B2 => 
                           n18855, ZN => n16407);
   U16652 : OAI221_X1 port map( B1 => n14222, B2 => n20956, C1 => n15288, C2 =>
                           n20950, A => n16388, ZN => n16383);
   U16653 : AOI22_X1 port map( A1 => n20944, A2 => n18834, B1 => n20938, B2 => 
                           n18835, ZN => n16388);
   U16654 : OAI221_X1 port map( B1 => n14221, B2 => n20956, C1 => n15287, C2 =>
                           n20950, A => n16369, ZN => n16364);
   U16655 : AOI22_X1 port map( A1 => n20944, A2 => n18814, B1 => n20938, B2 => 
                           n18815, ZN => n16369);
   U16656 : OAI221_X1 port map( B1 => n14220, B2 => n20956, C1 => n15286, C2 =>
                           n20950, A => n16350, ZN => n16345);
   U16657 : AOI22_X1 port map( A1 => n20944, A2 => n18794, B1 => n20938, B2 => 
                           n18795, ZN => n16350);
   U16658 : OAI221_X1 port map( B1 => n14219, B2 => n20956, C1 => n15285, C2 =>
                           n20950, A => n16331, ZN => n16326);
   U16659 : AOI22_X1 port map( A1 => n20944, A2 => n18774, B1 => n20938, B2 => 
                           n18775, ZN => n16331);
   U16660 : OAI221_X1 port map( B1 => n14218, B2 => n20956, C1 => n15284, C2 =>
                           n20950, A => n16312, ZN => n16307);
   U16661 : AOI22_X1 port map( A1 => n20944, A2 => n18754, B1 => n20938, B2 => 
                           n18755, ZN => n16312);
   U16662 : OAI221_X1 port map( B1 => n14217, B2 => n20956, C1 => n15283, C2 =>
                           n20950, A => n16293, ZN => n16288);
   U16663 : AOI22_X1 port map( A1 => n20944, A2 => n18734, B1 => n20938, B2 => 
                           n18735, ZN => n16293);
   U16664 : OAI221_X1 port map( B1 => n14216, B2 => n20956, C1 => n15282, C2 =>
                           n20950, A => n16274, ZN => n16269);
   U16665 : AOI22_X1 port map( A1 => n20944, A2 => n18714, B1 => n20938, B2 => 
                           n18715, ZN => n16274);
   U16666 : OAI221_X1 port map( B1 => n14215, B2 => n20956, C1 => n15281, C2 =>
                           n20950, A => n16255, ZN => n16250);
   U16667 : AOI22_X1 port map( A1 => n20944, A2 => n18694, B1 => n20938, B2 => 
                           n18695, ZN => n16255);
   U16668 : OAI221_X1 port map( B1 => n14214, B2 => n20956, C1 => n15280, C2 =>
                           n20950, A => n16236, ZN => n16231);
   U16669 : AOI22_X1 port map( A1 => n20944, A2 => n18674, B1 => n20938, B2 => 
                           n18675, ZN => n16236);
   U16670 : OAI221_X1 port map( B1 => n14213, B2 => n20956, C1 => n15279, C2 =>
                           n20950, A => n16217, ZN => n16212);
   U16671 : AOI22_X1 port map( A1 => n20944, A2 => n18654, B1 => n20938, B2 => 
                           n18655, ZN => n16217);
   U16672 : OAI221_X1 port map( B1 => n14212, B2 => n20956, C1 => n15278, C2 =>
                           n20950, A => n16198, ZN => n16193);
   U16673 : AOI22_X1 port map( A1 => n20944, A2 => n18634, B1 => n20938, B2 => 
                           n18635, ZN => n16198);
   U16674 : OAI221_X1 port map( B1 => n15409, B2 => n20861, C1 => n16008, C2 =>
                           n20855, A => n17433, ZN => n17428);
   U16675 : AOI22_X1 port map( A1 => n20849, A2 => n8971, B1 => n20843, B2 => 
                           n8587, ZN => n17433);
   U16676 : OAI221_X1 port map( B1 => n14211, B2 => n20765, C1 => n15277, C2 =>
                           n20759, A => n17441, ZN => n17436);
   U16677 : AOI22_X1 port map( A1 => n20753, A2 => n18614, B1 => n20747, B2 => 
                           n18615, ZN => n17441);
   U16678 : OAI221_X1 port map( B1 => n15408, B2 => n20861, C1 => n16007, C2 =>
                           n20855, A => n17415, ZN => n17410);
   U16679 : AOI22_X1 port map( A1 => n20849, A2 => n8967, B1 => n20843, B2 => 
                           n8583, ZN => n17415);
   U16680 : OAI221_X1 port map( B1 => n14210, B2 => n20765, C1 => n15276, C2 =>
                           n20759, A => n17423, ZN => n17418);
   U16681 : AOI22_X1 port map( A1 => n20753, A2 => n18594, B1 => n20747, B2 => 
                           n18595, ZN => n17423);
   U16682 : OAI221_X1 port map( B1 => n15407, B2 => n20861, C1 => n16006, C2 =>
                           n20855, A => n17397, ZN => n17392);
   U16683 : AOI22_X1 port map( A1 => n20849, A2 => n8963, B1 => n20843, B2 => 
                           n8579, ZN => n17397);
   U16684 : OAI221_X1 port map( B1 => n14209, B2 => n20765, C1 => n15275, C2 =>
                           n20759, A => n17405, ZN => n17400);
   U16685 : AOI22_X1 port map( A1 => n20753, A2 => n18574, B1 => n20747, B2 => 
                           n18575, ZN => n17405);
   U16686 : OAI221_X1 port map( B1 => n15405, B2 => n20861, C1 => n16004, C2 =>
                           n20855, A => n17357, ZN => n17342);
   U16687 : AOI22_X1 port map( A1 => n20849, A2 => n8959, B1 => n20843, B2 => 
                           n8575, ZN => n17357);
   U16688 : OAI221_X1 port map( B1 => n14207, B2 => n20765, C1 => n15273, C2 =>
                           n20759, A => n17381, ZN => n17367);
   U16689 : AOI22_X1 port map( A1 => n20753, A2 => n18554, B1 => n20747, B2 => 
                           n18555, ZN => n17381);
   U16690 : OAI221_X1 port map( B1 => n15409, B2 => n21066, C1 => n16008, C2 =>
                           n21060, A => n16171, ZN => n16166);
   U16691 : AOI22_X1 port map( A1 => n21054, A2 => n8971, B1 => n21048, B2 => 
                           n8587, ZN => n16171);
   U16692 : OAI221_X1 port map( B1 => n14211, B2 => n20957, C1 => n15277, C2 =>
                           n20951, A => n16179, ZN => n16174);
   U16693 : AOI22_X1 port map( A1 => n20945, A2 => n18614, B1 => n20939, B2 => 
                           n18615, ZN => n16179);
   U16694 : OAI221_X1 port map( B1 => n15408, B2 => n21066, C1 => n16007, C2 =>
                           n21060, A => n16152, ZN => n16147);
   U16695 : AOI22_X1 port map( A1 => n21054, A2 => n8967, B1 => n21048, B2 => 
                           n8583, ZN => n16152);
   U16696 : OAI221_X1 port map( B1 => n14210, B2 => n20957, C1 => n15276, C2 =>
                           n20951, A => n16160, ZN => n16155);
   U16697 : AOI22_X1 port map( A1 => n20945, A2 => n18594, B1 => n20939, B2 => 
                           n18595, ZN => n16160);
   U16698 : OAI221_X1 port map( B1 => n15407, B2 => n21066, C1 => n16006, C2 =>
                           n21060, A => n16133, ZN => n16128);
   U16699 : AOI22_X1 port map( A1 => n21054, A2 => n8963, B1 => n21048, B2 => 
                           n8579, ZN => n16133);
   U16700 : OAI221_X1 port map( B1 => n14209, B2 => n20957, C1 => n15275, C2 =>
                           n20951, A => n16141, ZN => n16136);
   U16701 : AOI22_X1 port map( A1 => n20945, A2 => n18574, B1 => n20939, B2 => 
                           n18575, ZN => n16141);
   U16702 : OAI221_X1 port map( B1 => n15405, B2 => n21066, C1 => n16004, C2 =>
                           n21060, A => n16091, ZN => n16075);
   U16703 : AOI22_X1 port map( A1 => n21054, A2 => n8959, B1 => n21048, B2 => 
                           n8575, ZN => n16091);
   U16704 : OAI221_X1 port map( B1 => n14207, B2 => n20957, C1 => n15273, C2 =>
                           n20951, A => n16116, ZN => n16101);
   U16705 : AOI22_X1 port map( A1 => n20945, A2 => n18554, B1 => n20939, B2 => 
                           n18555, ZN => n16116);
   U16706 : OAI221_X1 port map( B1 => n14125, B2 => n20833, C1 => n15656, C2 =>
                           n20827, A => n18298, ZN => n18291);
   U16707 : AOI222_X1 port map( A1 => n20821, A2 => n19561, B1 => n20815, B2 =>
                           n9161, C1 => n20809, C2 => n8777, ZN => n18298);
   U16708 : OAI221_X1 port map( B1 => n14124, B2 => n20833, C1 => n15655, C2 =>
                           n20827, A => n18280, ZN => n18273);
   U16709 : AOI222_X1 port map( A1 => n20821, A2 => n19541, B1 => n20815, B2 =>
                           n9157, C1 => n20809, C2 => n8773, ZN => n18280);
   U16710 : OAI221_X1 port map( B1 => n14123, B2 => n20833, C1 => n15654, C2 =>
                           n20827, A => n18262, ZN => n18255);
   U16711 : AOI222_X1 port map( A1 => n20821, A2 => n19521, B1 => n20815, B2 =>
                           n9153, C1 => n20809, C2 => n8769, ZN => n18262);
   U16712 : OAI221_X1 port map( B1 => n14122, B2 => n20833, C1 => n15653, C2 =>
                           n20827, A => n18244, ZN => n18237);
   U16713 : AOI222_X1 port map( A1 => n20821, A2 => n19501, B1 => n20815, B2 =>
                           n9149, C1 => n20809, C2 => n8765, ZN => n18244);
   U16714 : OAI221_X1 port map( B1 => n14121, B2 => n20833, C1 => n15652, C2 =>
                           n20827, A => n18226, ZN => n18219);
   U16715 : AOI222_X1 port map( A1 => n20821, A2 => n19481, B1 => n20815, B2 =>
                           n9145, C1 => n20809, C2 => n8761, ZN => n18226);
   U16716 : OAI221_X1 port map( B1 => n14120, B2 => n20833, C1 => n15651, C2 =>
                           n20827, A => n18208, ZN => n18201);
   U16717 : AOI222_X1 port map( A1 => n20821, A2 => n19461, B1 => n20815, B2 =>
                           n9141, C1 => n20809, C2 => n8757, ZN => n18208);
   U16718 : OAI221_X1 port map( B1 => n14119, B2 => n20833, C1 => n15650, C2 =>
                           n20827, A => n18190, ZN => n18183);
   U16719 : AOI222_X1 port map( A1 => n20821, A2 => n19441, B1 => n20815, B2 =>
                           n9137, C1 => n20809, C2 => n8753, ZN => n18190);
   U16720 : OAI221_X1 port map( B1 => n14118, B2 => n20833, C1 => n15649, C2 =>
                           n20827, A => n18172, ZN => n18165);
   U16721 : AOI222_X1 port map( A1 => n20821, A2 => n19421, B1 => n20815, B2 =>
                           n9133, C1 => n20809, C2 => n8749, ZN => n18172);
   U16722 : OAI221_X1 port map( B1 => n14117, B2 => n20833, C1 => n15648, C2 =>
                           n20827, A => n18154, ZN => n18147);
   U16723 : AOI222_X1 port map( A1 => n20821, A2 => n19401, B1 => n20815, B2 =>
                           n9129, C1 => n20809, C2 => n8745, ZN => n18154);
   U16724 : OAI221_X1 port map( B1 => n14116, B2 => n20833, C1 => n15647, C2 =>
                           n20827, A => n18136, ZN => n18129);
   U16725 : AOI222_X1 port map( A1 => n20821, A2 => n19381, B1 => n20815, B2 =>
                           n9125, C1 => n20809, C2 => n8741, ZN => n18136);
   U16726 : OAI221_X1 port map( B1 => n14115, B2 => n20833, C1 => n15646, C2 =>
                           n20827, A => n18118, ZN => n18111);
   U16727 : AOI222_X1 port map( A1 => n20821, A2 => n19361, B1 => n20815, B2 =>
                           n9121, C1 => n20809, C2 => n8737, ZN => n18118);
   U16728 : OAI221_X1 port map( B1 => n14114, B2 => n20833, C1 => n15645, C2 =>
                           n20827, A => n18100, ZN => n18093);
   U16729 : AOI222_X1 port map( A1 => n20821, A2 => n19341, B1 => n20815, B2 =>
                           n9117, C1 => n20809, C2 => n8733, ZN => n18100);
   U16730 : OAI221_X1 port map( B1 => n14113, B2 => n20834, C1 => n15644, C2 =>
                           n20828, A => n18082, ZN => n18075);
   U16731 : AOI222_X1 port map( A1 => n20822, A2 => n19321, B1 => n20816, B2 =>
                           n9113, C1 => n20810, C2 => n8729, ZN => n18082);
   U16732 : OAI221_X1 port map( B1 => n14112, B2 => n20834, C1 => n15643, C2 =>
                           n20828, A => n18064, ZN => n18057);
   U16733 : AOI222_X1 port map( A1 => n20822, A2 => n19301, B1 => n20816, B2 =>
                           n9109, C1 => n20810, C2 => n8725, ZN => n18064);
   U16734 : OAI221_X1 port map( B1 => n14111, B2 => n20834, C1 => n15642, C2 =>
                           n20828, A => n18046, ZN => n18039);
   U16735 : AOI222_X1 port map( A1 => n20822, A2 => n19281, B1 => n20816, B2 =>
                           n9105, C1 => n20810, C2 => n8721, ZN => n18046);
   U16736 : OAI221_X1 port map( B1 => n14110, B2 => n20834, C1 => n15641, C2 =>
                           n20828, A => n18028, ZN => n18021);
   U16737 : AOI222_X1 port map( A1 => n20822, A2 => n19261, B1 => n20816, B2 =>
                           n9101, C1 => n20810, C2 => n8717, ZN => n18028);
   U16738 : OAI221_X1 port map( B1 => n14109, B2 => n20834, C1 => n15640, C2 =>
                           n20828, A => n18010, ZN => n18003);
   U16739 : AOI222_X1 port map( A1 => n20822, A2 => n19241, B1 => n20816, B2 =>
                           n9097, C1 => n20810, C2 => n8713, ZN => n18010);
   U16740 : OAI221_X1 port map( B1 => n14108, B2 => n20834, C1 => n15639, C2 =>
                           n20828, A => n17992, ZN => n17985);
   U16741 : AOI222_X1 port map( A1 => n20822, A2 => n19221, B1 => n20816, B2 =>
                           n9093, C1 => n20810, C2 => n8709, ZN => n17992);
   U16742 : OAI221_X1 port map( B1 => n14107, B2 => n20834, C1 => n15638, C2 =>
                           n20828, A => n17974, ZN => n17967);
   U16743 : AOI222_X1 port map( A1 => n20822, A2 => n19201, B1 => n20816, B2 =>
                           n9089, C1 => n20810, C2 => n8705, ZN => n17974);
   U16744 : OAI221_X1 port map( B1 => n14106, B2 => n20834, C1 => n15637, C2 =>
                           n20828, A => n17956, ZN => n17949);
   U16745 : AOI222_X1 port map( A1 => n20822, A2 => n19181, B1 => n20816, B2 =>
                           n9085, C1 => n20810, C2 => n8701, ZN => n17956);
   U16746 : OAI221_X1 port map( B1 => n14105, B2 => n20834, C1 => n15636, C2 =>
                           n20828, A => n17938, ZN => n17931);
   U16747 : AOI222_X1 port map( A1 => n20822, A2 => n19161, B1 => n20816, B2 =>
                           n9081, C1 => n20810, C2 => n8697, ZN => n17938);
   U16748 : OAI221_X1 port map( B1 => n14104, B2 => n20834, C1 => n15635, C2 =>
                           n20828, A => n17920, ZN => n17913);
   U16749 : AOI222_X1 port map( A1 => n20822, A2 => n19141, B1 => n20816, B2 =>
                           n9077, C1 => n20810, C2 => n8693, ZN => n17920);
   U16750 : OAI221_X1 port map( B1 => n14103, B2 => n20834, C1 => n15634, C2 =>
                           n20828, A => n17902, ZN => n17895);
   U16751 : AOI222_X1 port map( A1 => n20822, A2 => n19121, B1 => n20816, B2 =>
                           n9073, C1 => n20810, C2 => n8689, ZN => n17902);
   U16752 : OAI221_X1 port map( B1 => n14102, B2 => n20834, C1 => n15633, C2 =>
                           n20828, A => n17884, ZN => n17877);
   U16753 : AOI222_X1 port map( A1 => n20822, A2 => n19101, B1 => n20816, B2 =>
                           n9069, C1 => n20810, C2 => n8685, ZN => n17884);
   U16754 : OAI221_X1 port map( B1 => n14101, B2 => n20835, C1 => n15632, C2 =>
                           n20829, A => n17866, ZN => n17859);
   U16755 : AOI222_X1 port map( A1 => n20823, A2 => n19081, B1 => n20817, B2 =>
                           n9065, C1 => n20811, C2 => n8681, ZN => n17866);
   U16756 : OAI221_X1 port map( B1 => n14100, B2 => n20835, C1 => n15631, C2 =>
                           n20829, A => n17848, ZN => n17841);
   U16757 : AOI222_X1 port map( A1 => n20823, A2 => n19061, B1 => n20817, B2 =>
                           n9061, C1 => n20811, C2 => n8677, ZN => n17848);
   U16758 : OAI221_X1 port map( B1 => n14099, B2 => n20835, C1 => n15630, C2 =>
                           n20829, A => n17830, ZN => n17823);
   U16759 : AOI222_X1 port map( A1 => n20823, A2 => n19041, B1 => n20817, B2 =>
                           n9057, C1 => n20811, C2 => n8673, ZN => n17830);
   U16760 : OAI221_X1 port map( B1 => n14098, B2 => n20835, C1 => n15629, C2 =>
                           n20829, A => n17812, ZN => n17805);
   U16761 : AOI222_X1 port map( A1 => n20823, A2 => n19021, B1 => n20817, B2 =>
                           n9053, C1 => n20811, C2 => n8669, ZN => n17812);
   U16762 : OAI221_X1 port map( B1 => n14097, B2 => n20835, C1 => n15628, C2 =>
                           n20829, A => n17794, ZN => n17787);
   U16763 : AOI222_X1 port map( A1 => n20823, A2 => n19001, B1 => n20817, B2 =>
                           n9049, C1 => n20811, C2 => n8665, ZN => n17794);
   U16764 : OAI221_X1 port map( B1 => n14096, B2 => n20835, C1 => n15627, C2 =>
                           n20829, A => n17776, ZN => n17769);
   U16765 : AOI222_X1 port map( A1 => n20823, A2 => n18981, B1 => n20817, B2 =>
                           n9045, C1 => n20811, C2 => n8661, ZN => n17776);
   U16766 : OAI221_X1 port map( B1 => n14095, B2 => n20835, C1 => n15626, C2 =>
                           n20829, A => n17758, ZN => n17751);
   U16767 : AOI222_X1 port map( A1 => n20823, A2 => n18961, B1 => n20817, B2 =>
                           n9041, C1 => n20811, C2 => n8657, ZN => n17758);
   U16768 : OAI221_X1 port map( B1 => n14094, B2 => n20835, C1 => n15625, C2 =>
                           n20829, A => n17740, ZN => n17733);
   U16769 : AOI222_X1 port map( A1 => n20823, A2 => n18941, B1 => n20817, B2 =>
                           n9037, C1 => n20811, C2 => n8653, ZN => n17740);
   U16770 : OAI221_X1 port map( B1 => n14093, B2 => n20835, C1 => n15624, C2 =>
                           n20829, A => n17722, ZN => n17715);
   U16771 : AOI222_X1 port map( A1 => n20823, A2 => n18921, B1 => n20817, B2 =>
                           n9033, C1 => n20811, C2 => n8649, ZN => n17722);
   U16772 : OAI221_X1 port map( B1 => n14092, B2 => n20835, C1 => n15623, C2 =>
                           n20829, A => n17704, ZN => n17697);
   U16773 : AOI222_X1 port map( A1 => n20823, A2 => n18901, B1 => n20817, B2 =>
                           n9029, C1 => n20811, C2 => n8645, ZN => n17704);
   U16774 : OAI221_X1 port map( B1 => n14091, B2 => n20835, C1 => n15622, C2 =>
                           n20829, A => n17686, ZN => n17679);
   U16775 : AOI222_X1 port map( A1 => n20823, A2 => n18881, B1 => n20817, B2 =>
                           n9025, C1 => n20811, C2 => n8641, ZN => n17686);
   U16776 : OAI221_X1 port map( B1 => n14090, B2 => n20835, C1 => n15621, C2 =>
                           n20829, A => n17668, ZN => n17661);
   U16777 : AOI222_X1 port map( A1 => n20823, A2 => n18861, B1 => n20817, B2 =>
                           n9021, C1 => n20811, C2 => n8637, ZN => n17668);
   U16778 : OAI221_X1 port map( B1 => n14089, B2 => n20836, C1 => n15620, C2 =>
                           n20830, A => n17650, ZN => n17643);
   U16779 : AOI222_X1 port map( A1 => n20824, A2 => n18841, B1 => n20818, B2 =>
                           n9017, C1 => n20812, C2 => n8633, ZN => n17650);
   U16780 : OAI221_X1 port map( B1 => n14088, B2 => n20836, C1 => n15619, C2 =>
                           n20830, A => n17632, ZN => n17625);
   U16781 : AOI222_X1 port map( A1 => n20824, A2 => n18821, B1 => n20818, B2 =>
                           n9013, C1 => n20812, C2 => n8629, ZN => n17632);
   U16782 : OAI221_X1 port map( B1 => n14087, B2 => n20836, C1 => n15618, C2 =>
                           n20830, A => n17614, ZN => n17607);
   U16783 : AOI222_X1 port map( A1 => n20824, A2 => n18801, B1 => n20818, B2 =>
                           n9009, C1 => n20812, C2 => n8625, ZN => n17614);
   U16784 : OAI221_X1 port map( B1 => n14086, B2 => n20836, C1 => n15617, C2 =>
                           n20830, A => n17596, ZN => n17589);
   U16785 : AOI222_X1 port map( A1 => n20824, A2 => n18781, B1 => n20818, B2 =>
                           n9005, C1 => n20812, C2 => n8621, ZN => n17596);
   U16786 : OAI221_X1 port map( B1 => n14085, B2 => n20836, C1 => n15616, C2 =>
                           n20830, A => n17578, ZN => n17571);
   U16787 : AOI222_X1 port map( A1 => n20824, A2 => n18761, B1 => n20818, B2 =>
                           n9001, C1 => n20812, C2 => n8617, ZN => n17578);
   U16788 : OAI221_X1 port map( B1 => n14084, B2 => n20836, C1 => n15615, C2 =>
                           n20830, A => n17560, ZN => n17553);
   U16789 : AOI222_X1 port map( A1 => n20824, A2 => n18741, B1 => n20818, B2 =>
                           n8997, C1 => n20812, C2 => n8613, ZN => n17560);
   U16790 : OAI221_X1 port map( B1 => n14083, B2 => n20836, C1 => n15614, C2 =>
                           n20830, A => n17542, ZN => n17535);
   U16791 : AOI222_X1 port map( A1 => n20824, A2 => n18721, B1 => n20818, B2 =>
                           n8993, C1 => n20812, C2 => n8609, ZN => n17542);
   U16792 : OAI221_X1 port map( B1 => n14082, B2 => n20836, C1 => n15613, C2 =>
                           n20830, A => n17524, ZN => n17517);
   U16793 : AOI222_X1 port map( A1 => n20824, A2 => n18701, B1 => n20818, B2 =>
                           n8989, C1 => n20812, C2 => n8605, ZN => n17524);
   U16794 : OAI221_X1 port map( B1 => n14081, B2 => n20836, C1 => n15612, C2 =>
                           n20830, A => n17506, ZN => n17499);
   U16795 : AOI222_X1 port map( A1 => n20824, A2 => n18681, B1 => n20818, B2 =>
                           n8985, C1 => n20812, C2 => n8601, ZN => n17506);
   U16796 : OAI221_X1 port map( B1 => n14080, B2 => n20836, C1 => n15611, C2 =>
                           n20830, A => n17488, ZN => n17481);
   U16797 : AOI222_X1 port map( A1 => n20824, A2 => n18661, B1 => n20818, B2 =>
                           n8981, C1 => n20812, C2 => n8597, ZN => n17488);
   U16798 : OAI221_X1 port map( B1 => n14079, B2 => n20836, C1 => n15610, C2 =>
                           n20830, A => n17470, ZN => n17463);
   U16799 : AOI222_X1 port map( A1 => n20824, A2 => n18641, B1 => n20818, B2 =>
                           n8977, C1 => n20812, C2 => n8593, ZN => n17470);
   U16800 : OAI221_X1 port map( B1 => n14078, B2 => n20836, C1 => n15609, C2 =>
                           n20830, A => n17452, ZN => n17445);
   U16801 : AOI222_X1 port map( A1 => n20824, A2 => n18621, B1 => n20818, B2 =>
                           n8973, C1 => n20812, C2 => n8589, ZN => n17452);
   U16802 : OAI221_X1 port map( B1 => n14077, B2 => n20837, C1 => n15608, C2 =>
                           n20831, A => n17434, ZN => n17427);
   U16803 : AOI222_X1 port map( A1 => n20825, A2 => n18601, B1 => n20819, B2 =>
                           n8969, C1 => n20813, C2 => n8585, ZN => n17434);
   U16804 : OAI221_X1 port map( B1 => n14076, B2 => n20837, C1 => n15607, C2 =>
                           n20831, A => n17416, ZN => n17409);
   U16805 : AOI222_X1 port map( A1 => n20825, A2 => n18581, B1 => n20819, B2 =>
                           n8965, C1 => n20813, C2 => n8581, ZN => n17416);
   U16806 : OAI221_X1 port map( B1 => n14075, B2 => n20837, C1 => n15606, C2 =>
                           n20831, A => n17398, ZN => n17391);
   U16807 : AOI222_X1 port map( A1 => n20825, A2 => n18561, B1 => n20819, B2 =>
                           n8961, C1 => n20813, C2 => n8577, ZN => n17398);
   U16808 : OAI221_X1 port map( B1 => n14073, B2 => n20837, C1 => n15604, C2 =>
                           n20831, A => n17362, ZN => n17341);
   U16809 : AOI222_X1 port map( A1 => n20825, A2 => n18541, B1 => n20819, B2 =>
                           n8957, C1 => n20813, C2 => n8573, ZN => n17362);
   U16810 : OAI221_X1 port map( B1 => n14077, B2 => n21042, C1 => n15608, C2 =>
                           n21036, A => n16172, ZN => n16165);
   U16811 : AOI222_X1 port map( A1 => n21030, A2 => n18601, B1 => n21024, B2 =>
                           n8969, C1 => n21018, C2 => n8585, ZN => n16172);
   U16812 : OAI221_X1 port map( B1 => n14076, B2 => n21042, C1 => n15607, C2 =>
                           n21036, A => n16153, ZN => n16146);
   U16813 : AOI222_X1 port map( A1 => n21030, A2 => n18581, B1 => n21024, B2 =>
                           n8965, C1 => n21018, C2 => n8581, ZN => n16153);
   U16814 : OAI221_X1 port map( B1 => n14075, B2 => n21042, C1 => n15606, C2 =>
                           n21036, A => n16134, ZN => n16127);
   U16815 : AOI222_X1 port map( A1 => n21030, A2 => n18561, B1 => n21024, B2 =>
                           n8961, C1 => n21018, C2 => n8577, ZN => n16134);
   U16816 : OAI221_X1 port map( B1 => n14073, B2 => n21042, C1 => n15604, C2 =>
                           n21036, A => n16096, ZN => n16074);
   U16817 : AOI222_X1 port map( A1 => n21030, A2 => n18541, B1 => n21024, B2 =>
                           n8957, C1 => n21018, C2 => n8573, ZN => n16096);
   U16818 : OAI221_X1 port map( B1 => n15469, B2 => n20856, C1 => n16068, C2 =>
                           n20850, A => n18522, ZN => n18508);
   U16819 : AOI22_X1 port map( A1 => n20844, A2 => n9211, B1 => n20838, B2 => 
                           n8827, ZN => n18522);
   U16820 : OAI221_X1 port map( B1 => n15468, B2 => n20856, C1 => n16067, C2 =>
                           n20850, A => n18495, ZN => n18490);
   U16821 : AOI22_X1 port map( A1 => n20844, A2 => n9207, B1 => n20838, B2 => 
                           n8823, ZN => n18495);
   U16822 : OAI221_X1 port map( B1 => n15467, B2 => n20856, C1 => n16066, C2 =>
                           n20850, A => n18477, ZN => n18472);
   U16823 : AOI22_X1 port map( A1 => n20844, A2 => n9203, B1 => n20838, B2 => 
                           n8819, ZN => n18477);
   U16824 : OAI221_X1 port map( B1 => n15466, B2 => n20856, C1 => n16065, C2 =>
                           n20850, A => n18459, ZN => n18454);
   U16825 : AOI22_X1 port map( A1 => n20844, A2 => n9199, B1 => n20838, B2 => 
                           n8815, ZN => n18459);
   U16826 : OAI221_X1 port map( B1 => n15465, B2 => n20856, C1 => n16064, C2 =>
                           n20850, A => n18441, ZN => n18436);
   U16827 : AOI22_X1 port map( A1 => n20844, A2 => n9195, B1 => n20838, B2 => 
                           n8811, ZN => n18441);
   U16828 : OAI221_X1 port map( B1 => n15464, B2 => n20856, C1 => n16063, C2 =>
                           n20850, A => n18423, ZN => n18418);
   U16829 : AOI22_X1 port map( A1 => n20844, A2 => n9191, B1 => n20838, B2 => 
                           n8807, ZN => n18423);
   U16830 : OAI221_X1 port map( B1 => n15463, B2 => n20856, C1 => n16062, C2 =>
                           n20850, A => n18405, ZN => n18400);
   U16831 : AOI22_X1 port map( A1 => n20844, A2 => n9187, B1 => n20838, B2 => 
                           n8803, ZN => n18405);
   U16832 : OAI221_X1 port map( B1 => n15462, B2 => n20856, C1 => n16061, C2 =>
                           n20850, A => n18387, ZN => n18382);
   U16833 : AOI22_X1 port map( A1 => n20844, A2 => n9183, B1 => n20838, B2 => 
                           n8799, ZN => n18387);
   U16834 : OAI221_X1 port map( B1 => n15461, B2 => n20856, C1 => n16060, C2 =>
                           n20850, A => n18369, ZN => n18364);
   U16835 : AOI22_X1 port map( A1 => n20844, A2 => n9179, B1 => n20838, B2 => 
                           n8795, ZN => n18369);
   U16836 : OAI221_X1 port map( B1 => n15460, B2 => n20856, C1 => n16059, C2 =>
                           n20850, A => n18351, ZN => n18346);
   U16837 : AOI22_X1 port map( A1 => n20844, A2 => n9175, B1 => n20838, B2 => 
                           n8791, ZN => n18351);
   U16838 : OAI221_X1 port map( B1 => n15459, B2 => n20856, C1 => n16058, C2 =>
                           n20850, A => n18333, ZN => n18328);
   U16839 : AOI22_X1 port map( A1 => n20844, A2 => n9171, B1 => n20838, B2 => 
                           n8787, ZN => n18333);
   U16840 : OAI221_X1 port map( B1 => n15458, B2 => n20856, C1 => n16057, C2 =>
                           n20850, A => n18315, ZN => n18310);
   U16841 : AOI22_X1 port map( A1 => n20844, A2 => n9167, B1 => n20838, B2 => 
                           n8783, ZN => n18315);
   U16842 : OAI221_X1 port map( B1 => n14137, B2 => n20832, C1 => n15668, C2 =>
                           n20826, A => n18525, ZN => n18507);
   U16843 : AOI222_X1 port map( A1 => n20820, A2 => n19801, B1 => n20814, B2 =>
                           n9209, C1 => n20808, C2 => n8825, ZN => n18525);
   U16844 : OAI221_X1 port map( B1 => n14136, B2 => n20832, C1 => n15667, C2 =>
                           n20826, A => n18496, ZN => n18489);
   U16845 : AOI222_X1 port map( A1 => n20820, A2 => n19781, B1 => n20814, B2 =>
                           n9205, C1 => n20808, C2 => n8821, ZN => n18496);
   U16846 : OAI221_X1 port map( B1 => n14135, B2 => n20832, C1 => n15666, C2 =>
                           n20826, A => n18478, ZN => n18471);
   U16847 : AOI222_X1 port map( A1 => n20820, A2 => n19761, B1 => n20814, B2 =>
                           n9201, C1 => n20808, C2 => n8817, ZN => n18478);
   U16848 : OAI221_X1 port map( B1 => n14134, B2 => n20832, C1 => n15665, C2 =>
                           n20826, A => n18460, ZN => n18453);
   U16849 : AOI222_X1 port map( A1 => n20820, A2 => n19741, B1 => n20814, B2 =>
                           n9197, C1 => n20808, C2 => n8813, ZN => n18460);
   U16850 : OAI221_X1 port map( B1 => n14133, B2 => n20832, C1 => n15664, C2 =>
                           n20826, A => n18442, ZN => n18435);
   U16851 : AOI222_X1 port map( A1 => n20820, A2 => n19721, B1 => n20814, B2 =>
                           n9193, C1 => n20808, C2 => n8809, ZN => n18442);
   U16852 : OAI221_X1 port map( B1 => n14132, B2 => n20832, C1 => n15663, C2 =>
                           n20826, A => n18424, ZN => n18417);
   U16853 : AOI222_X1 port map( A1 => n20820, A2 => n19701, B1 => n20814, B2 =>
                           n9189, C1 => n20808, C2 => n8805, ZN => n18424);
   U16854 : OAI221_X1 port map( B1 => n14131, B2 => n20832, C1 => n15662, C2 =>
                           n20826, A => n18406, ZN => n18399);
   U16855 : AOI222_X1 port map( A1 => n20820, A2 => n19681, B1 => n20814, B2 =>
                           n9185, C1 => n20808, C2 => n8801, ZN => n18406);
   U16856 : OAI221_X1 port map( B1 => n14130, B2 => n20832, C1 => n15661, C2 =>
                           n20826, A => n18388, ZN => n18381);
   U16857 : AOI222_X1 port map( A1 => n20820, A2 => n19661, B1 => n20814, B2 =>
                           n9181, C1 => n20808, C2 => n8797, ZN => n18388);
   U16858 : OAI221_X1 port map( B1 => n14129, B2 => n20832, C1 => n15660, C2 =>
                           n20826, A => n18370, ZN => n18363);
   U16859 : AOI222_X1 port map( A1 => n20820, A2 => n19641, B1 => n20814, B2 =>
                           n9177, C1 => n20808, C2 => n8793, ZN => n18370);
   U16860 : OAI221_X1 port map( B1 => n14128, B2 => n20832, C1 => n15659, C2 =>
                           n20826, A => n18352, ZN => n18345);
   U16861 : AOI222_X1 port map( A1 => n20820, A2 => n19621, B1 => n20814, B2 =>
                           n9173, C1 => n20808, C2 => n8789, ZN => n18352);
   U16862 : OAI221_X1 port map( B1 => n14127, B2 => n20832, C1 => n15658, C2 =>
                           n20826, A => n18334, ZN => n18327);
   U16863 : AOI222_X1 port map( A1 => n20820, A2 => n19601, B1 => n20814, B2 =>
                           n9169, C1 => n20808, C2 => n8785, ZN => n18334);
   U16864 : OAI221_X1 port map( B1 => n14126, B2 => n20832, C1 => n15657, C2 =>
                           n20826, A => n18316, ZN => n18309);
   U16865 : AOI222_X1 port map( A1 => n20820, A2 => n19581, B1 => n20814, B2 =>
                           n9165, C1 => n20808, C2 => n8781, ZN => n18316);
   U16866 : NOR2_X1 port map( A1 => RD2, A2 => RD1, ZN => n18540);
   U16867 : INV_X1 port map( A => n16083, ZN => n16076);
   U16868 : AOI221_X1 port map( B1 => n18544, B2 => n21091, C1 => n18545, C2 =>
                           n21081, A => n16086, ZN => n16083);
   U16869 : OAI22_X1 port map( A1 => n21073, A2 => n14542, B1 => n21072, B2 => 
                           n14874, ZN => n16086);
   U16870 : NOR2_X1 port map( A1 => n15071, A2 => ADD_WR(4), ZN => n14474);
   U16871 : NOR2_X1 port map( A1 => n17303, A2 => n15071, ZN => n15536);
   U16872 : INV_X1 port map( A => ADD_WR(4), ZN => n17303);
   U16873 : OAI22_X1 port map( A1 => n21727, A2 => n14043, B1 => n21719, B2 => 
                           n21562, ZN => n7369);
   U16874 : OAI22_X1 port map( A1 => n21727, A2 => n14041, B1 => n21719, B2 => 
                           n21565, ZN => n7370);
   U16875 : OAI22_X1 port map( A1 => n21727, A2 => n14039, B1 => n21719, B2 => 
                           n21568, ZN => n7371);
   U16876 : OAI22_X1 port map( A1 => n21727, A2 => n14037, B1 => n21719, B2 => 
                           n21571, ZN => n7372);
   U16877 : OAI22_X1 port map( A1 => n21727, A2 => n14035, B1 => n21719, B2 => 
                           n21574, ZN => n7373);
   U16878 : OAI22_X1 port map( A1 => n21727, A2 => n14033, B1 => n21719, B2 => 
                           n21577, ZN => n7374);
   U16879 : OAI22_X1 port map( A1 => n21727, A2 => n14031, B1 => n21719, B2 => 
                           n21580, ZN => n7375);
   U16880 : OAI22_X1 port map( A1 => n21727, A2 => n14029, B1 => n21719, B2 => 
                           n21583, ZN => n7376);
   U16881 : OAI22_X1 port map( A1 => n21727, A2 => n14027, B1 => n21719, B2 => 
                           n21586, ZN => n7377);
   U16882 : OAI22_X1 port map( A1 => n21727, A2 => n14025, B1 => n21719, B2 => 
                           n21589, ZN => n7378);
   U16883 : OAI22_X1 port map( A1 => n21727, A2 => n14023, B1 => n21719, B2 => 
                           n21592, ZN => n7379);
   U16884 : OAI22_X1 port map( A1 => n21727, A2 => n14021, B1 => n21719, B2 => 
                           n21595, ZN => n7380);
   U16885 : OAI22_X1 port map( A1 => n21727, A2 => n14019, B1 => n21720, B2 => 
                           n21598, ZN => n7381);
   U16886 : OAI22_X1 port map( A1 => n21728, A2 => n14017, B1 => n21720, B2 => 
                           n21601, ZN => n7382);
   U16887 : OAI22_X1 port map( A1 => n21728, A2 => n14015, B1 => n21720, B2 => 
                           n21604, ZN => n7383);
   U16888 : OAI22_X1 port map( A1 => n21728, A2 => n14013, B1 => n21720, B2 => 
                           n21607, ZN => n7384);
   U16889 : OAI22_X1 port map( A1 => n21728, A2 => n14011, B1 => n21720, B2 => 
                           n21610, ZN => n7385);
   U16890 : OAI22_X1 port map( A1 => n21728, A2 => n14009, B1 => n21720, B2 => 
                           n21613, ZN => n7386);
   U16891 : OAI22_X1 port map( A1 => n21728, A2 => n14007, B1 => n21720, B2 => 
                           n21616, ZN => n7387);
   U16892 : OAI22_X1 port map( A1 => n21728, A2 => n14005, B1 => n21720, B2 => 
                           n21619, ZN => n7388);
   U16893 : OAI22_X1 port map( A1 => n21728, A2 => n14003, B1 => n21720, B2 => 
                           n21622, ZN => n7389);
   U16894 : OAI22_X1 port map( A1 => n21728, A2 => n14001, B1 => n21720, B2 => 
                           n21625, ZN => n7390);
   U16895 : OAI22_X1 port map( A1 => n21728, A2 => n13999, B1 => n21720, B2 => 
                           n21628, ZN => n7391);
   U16896 : OAI22_X1 port map( A1 => n21728, A2 => n13997, B1 => n21720, B2 => 
                           n21631, ZN => n7392);
   U16897 : OAI22_X1 port map( A1 => n21728, A2 => n13995, B1 => n21721, B2 => 
                           n21634, ZN => n7393);
   U16898 : OAI22_X1 port map( A1 => n21728, A2 => n13993, B1 => n21721, B2 => 
                           n21637, ZN => n7394);
   U16899 : OAI22_X1 port map( A1 => n21729, A2 => n13991, B1 => n21721, B2 => 
                           n21640, ZN => n7395);
   U16900 : OAI22_X1 port map( A1 => n21729, A2 => n13989, B1 => n21721, B2 => 
                           n21643, ZN => n7396);
   U16901 : OAI22_X1 port map( A1 => n21729, A2 => n13987, B1 => n21721, B2 => 
                           n21646, ZN => n7397);
   U16902 : OAI22_X1 port map( A1 => n21729, A2 => n13985, B1 => n21721, B2 => 
                           n21649, ZN => n7398);
   U16903 : OAI22_X1 port map( A1 => n21729, A2 => n13983, B1 => n21721, B2 => 
                           n21652, ZN => n7399);
   U16904 : OAI22_X1 port map( A1 => n21729, A2 => n13981, B1 => n21721, B2 => 
                           n21655, ZN => n7400);
   U16905 : OAI22_X1 port map( A1 => n21729, A2 => n13979, B1 => n21721, B2 => 
                           n21658, ZN => n7401);
   U16906 : OAI22_X1 port map( A1 => n21729, A2 => n13977, B1 => n21721, B2 => 
                           n21661, ZN => n7402);
   U16907 : OAI22_X1 port map( A1 => n21729, A2 => n13975, B1 => n21721, B2 => 
                           n21664, ZN => n7403);
   U16908 : OAI22_X1 port map( A1 => n21729, A2 => n13973, B1 => n21721, B2 => 
                           n21667, ZN => n7404);
   U16909 : OAI22_X1 port map( A1 => n21729, A2 => n13971, B1 => n21722, B2 => 
                           n21670, ZN => n7405);
   U16910 : OAI22_X1 port map( A1 => n21729, A2 => n13969, B1 => n21722, B2 => 
                           n21673, ZN => n7406);
   U16911 : OAI22_X1 port map( A1 => n21729, A2 => n13967, B1 => n21722, B2 => 
                           n21676, ZN => n7407);
   U16912 : OAI22_X1 port map( A1 => n21730, A2 => n13965, B1 => n21722, B2 => 
                           n21679, ZN => n7408);
   U16913 : OAI22_X1 port map( A1 => n21730, A2 => n13963, B1 => n21722, B2 => 
                           n21682, ZN => n7409);
   U16914 : OAI22_X1 port map( A1 => n21730, A2 => n13961, B1 => n21722, B2 => 
                           n21685, ZN => n7410);
   U16915 : OAI22_X1 port map( A1 => n21730, A2 => n13959, B1 => n21722, B2 => 
                           n21688, ZN => n7411);
   U16916 : OAI22_X1 port map( A1 => n21730, A2 => n13957, B1 => n21722, B2 => 
                           n21691, ZN => n7412);
   U16917 : OAI22_X1 port map( A1 => n21730, A2 => n13955, B1 => n21722, B2 => 
                           n21694, ZN => n7413);
   U16918 : OAI22_X1 port map( A1 => n21730, A2 => n13953, B1 => n21722, B2 => 
                           n21697, ZN => n7414);
   U16919 : OAI22_X1 port map( A1 => n21730, A2 => n13951, B1 => n21722, B2 => 
                           n21700, ZN => n7415);
   U16920 : OAI22_X1 port map( A1 => n21730, A2 => n13949, B1 => n21722, B2 => 
                           n21703, ZN => n7416);
   U16921 : OAI22_X1 port map( A1 => n21730, A2 => n13947, B1 => n21723, B2 => 
                           n21706, ZN => n7417);
   U16922 : OAI22_X1 port map( A1 => n21730, A2 => n13945, B1 => n21723, B2 => 
                           n21709, ZN => n7418);
   U16923 : OAI22_X1 port map( A1 => n21730, A2 => n13943, B1 => n21723, B2 => 
                           n21712, ZN => n7419);
   U16924 : OAI22_X1 port map( A1 => n21730, A2 => n13940, B1 => n21723, B2 => 
                           n21715, ZN => n7420);
   U16925 : OAI221_X1 port map( B1 => n14546, B2 => n21073, C1 => n14878, C2 =>
                           n21072, A => n16170, ZN => n16167);
   U16926 : AOI22_X1 port map( A1 => n18604, A2 => n21091, B1 => n21081, B2 => 
                           n18605, ZN => n16170);
   U16927 : OAI221_X1 port map( B1 => n14545, B2 => n21073, C1 => n14877, C2 =>
                           n21072, A => n16151, ZN => n16148);
   U16928 : AOI22_X1 port map( A1 => n18584, A2 => n21091, B1 => n21081, B2 => 
                           n18585, ZN => n16151);
   U16929 : OAI221_X1 port map( B1 => n14544, B2 => n21073, C1 => n14876, C2 =>
                           n21072, A => n16132, ZN => n16129);
   U16930 : AOI22_X1 port map( A1 => n18564, A2 => n21091, B1 => n21081, B2 => 
                           n18565, ZN => n16132);
   U16931 : OAI22_X1 port map( A1 => n21154, A2 => n15942, B1 => n21708, B2 => 
                           n21147, ZN => n5561);
   U16932 : OAI22_X1 port map( A1 => n21154, A2 => n15941, B1 => n21711, B2 => 
                           n21147, ZN => n5562);
   U16933 : OAI22_X1 port map( A1 => n21154, A2 => n15940, B1 => n21714, B2 => 
                           n21147, ZN => n5563);
   U16934 : OAI22_X1 port map( A1 => n21154, A2 => n15938, B1 => n21717, B2 => 
                           n21147, ZN => n5564);
   U16935 : OAI22_X1 port map( A1 => n21180, A2 => n15810, B1 => n21708, B2 => 
                           n21173, ZN => n5689);
   U16936 : OAI22_X1 port map( A1 => n21180, A2 => n15809, B1 => n21711, B2 => 
                           n21173, ZN => n5690);
   U16937 : OAI22_X1 port map( A1 => n21180, A2 => n15808, B1 => n21714, B2 => 
                           n21173, ZN => n5691);
   U16938 : OAI22_X1 port map( A1 => n21180, A2 => n15806, B1 => n21717, B2 => 
                           n21173, ZN => n5692);
   U16939 : OAI22_X1 port map( A1 => n21206, A2 => n15675, B1 => n21708, B2 => 
                           n21199, ZN => n5817);
   U16940 : OAI22_X1 port map( A1 => n21206, A2 => n15674, B1 => n21711, B2 => 
                           n21199, ZN => n5818);
   U16941 : OAI22_X1 port map( A1 => n21206, A2 => n15673, B1 => n21714, B2 => 
                           n21199, ZN => n5819);
   U16942 : OAI22_X1 port map( A1 => n21206, A2 => n15671, B1 => n21717, B2 => 
                           n21199, ZN => n5820);
   U16943 : OAI22_X1 port map( A1 => n21232, A2 => n15542, B1 => n21707, B2 => 
                           n21225, ZN => n5945);
   U16944 : OAI22_X1 port map( A1 => n21232, A2 => n15541, B1 => n21710, B2 => 
                           n21225, ZN => n5946);
   U16945 : OAI22_X1 port map( A1 => n21232, A2 => n15540, B1 => n21713, B2 => 
                           n21225, ZN => n5947);
   U16946 : OAI22_X1 port map( A1 => n21232, A2 => n15538, B1 => n21716, B2 => 
                           n21225, ZN => n5948);
   U16947 : OAI22_X1 port map( A1 => n21245, A2 => n15475, B1 => n21707, B2 => 
                           n21238, ZN => n6009);
   U16948 : OAI22_X1 port map( A1 => n21245, A2 => n15474, B1 => n21710, B2 => 
                           n21238, ZN => n6010);
   U16949 : OAI22_X1 port map( A1 => n21245, A2 => n15473, B1 => n21713, B2 => 
                           n21238, ZN => n6011);
   U16950 : OAI22_X1 port map( A1 => n21245, A2 => n15471, B1 => n21716, B2 => 
                           n21238, ZN => n6012);
   U16951 : OAI22_X1 port map( A1 => n21271, A2 => n15343, B1 => n21707, B2 => 
                           n21264, ZN => n6137);
   U16952 : OAI22_X1 port map( A1 => n21271, A2 => n15342, B1 => n21710, B2 => 
                           n21264, ZN => n6138);
   U16953 : OAI22_X1 port map( A1 => n21271, A2 => n15341, B1 => n21713, B2 => 
                           n21264, ZN => n6139);
   U16954 : OAI22_X1 port map( A1 => n21271, A2 => n15339, B1 => n21716, B2 => 
                           n21264, ZN => n6140);
   U16955 : OAI22_X1 port map( A1 => n21297, A2 => n15211, B1 => n21707, B2 => 
                           n21290, ZN => n6265);
   U16956 : OAI22_X1 port map( A1 => n21297, A2 => n15210, B1 => n21710, B2 => 
                           n21290, ZN => n6266);
   U16957 : OAI22_X1 port map( A1 => n21297, A2 => n15209, B1 => n21713, B2 => 
                           n21290, ZN => n6267);
   U16958 : OAI22_X1 port map( A1 => n21297, A2 => n15207, B1 => n21716, B2 => 
                           n21290, ZN => n6268);
   U16959 : OAI22_X1 port map( A1 => n21310, A2 => n15144, B1 => n21707, B2 => 
                           n21303, ZN => n6329);
   U16960 : OAI22_X1 port map( A1 => n21310, A2 => n15143, B1 => n21710, B2 => 
                           n21303, ZN => n6330);
   U16961 : OAI22_X1 port map( A1 => n21310, A2 => n15142, B1 => n21713, B2 => 
                           n21303, ZN => n6331);
   U16962 : OAI22_X1 port map( A1 => n21310, A2 => n15140, B1 => n21716, B2 => 
                           n21303, ZN => n6332);
   U16963 : OAI22_X1 port map( A1 => n21323, A2 => n15077, B1 => n21707, B2 => 
                           n21316, ZN => n6393);
   U16964 : OAI22_X1 port map( A1 => n21323, A2 => n15076, B1 => n21710, B2 => 
                           n21316, ZN => n6394);
   U16965 : OAI22_X1 port map( A1 => n21323, A2 => n15075, B1 => n21713, B2 => 
                           n21316, ZN => n6395);
   U16966 : OAI22_X1 port map( A1 => n21323, A2 => n15073, B1 => n21716, B2 => 
                           n21316, ZN => n6396);
   U16967 : OAI22_X1 port map( A1 => n21401, A2 => n14680, B1 => n21706, B2 => 
                           n21394, ZN => n6777);
   U16968 : OAI22_X1 port map( A1 => n21401, A2 => n14679, B1 => n21709, B2 => 
                           n21394, ZN => n6778);
   U16969 : OAI22_X1 port map( A1 => n21401, A2 => n14678, B1 => n21712, B2 => 
                           n21394, ZN => n6779);
   U16970 : OAI22_X1 port map( A1 => n21401, A2 => n14676, B1 => n21715, B2 => 
                           n21394, ZN => n6780);
   U16971 : OAI22_X1 port map( A1 => n21414, A2 => n14613, B1 => n21706, B2 => 
                           n21407, ZN => n6841);
   U16972 : OAI22_X1 port map( A1 => n21414, A2 => n14612, B1 => n21709, B2 => 
                           n21407, ZN => n6842);
   U16973 : OAI22_X1 port map( A1 => n21414, A2 => n14611, B1 => n21712, B2 => 
                           n21407, ZN => n6843);
   U16974 : OAI22_X1 port map( A1 => n21414, A2 => n14609, B1 => n21715, B2 => 
                           n21407, ZN => n6844);
   U16975 : OAI22_X1 port map( A1 => n21453, A2 => n14410, B1 => n21706, B2 => 
                           n21446, ZN => n7033);
   U16976 : OAI22_X1 port map( A1 => n21453, A2 => n14409, B1 => n21709, B2 => 
                           n21446, ZN => n7034);
   U16977 : OAI22_X1 port map( A1 => n21453, A2 => n14408, B1 => n21712, B2 => 
                           n21446, ZN => n7035);
   U16978 : OAI22_X1 port map( A1 => n21453, A2 => n14406, B1 => n21715, B2 => 
                           n21446, ZN => n7036);
   U16979 : OAI22_X1 port map( A1 => n21505, A2 => n14144, B1 => n21706, B2 => 
                           n21498, ZN => n7289);
   U16980 : OAI22_X1 port map( A1 => n21505, A2 => n14143, B1 => n21709, B2 => 
                           n21498, ZN => n7290);
   U16981 : OAI22_X1 port map( A1 => n21505, A2 => n14142, B1 => n21712, B2 => 
                           n21498, ZN => n7291);
   U16982 : OAI22_X1 port map( A1 => n21505, A2 => n14140, B1 => n21715, B2 => 
                           n21498, ZN => n7292);
   U16983 : AOI22_X1 port map( A1 => n20724, A2 => n19810, B1 => n20718, B2 => 
                           n19811, ZN => n18537);
   U16984 : AOI22_X1 port map( A1 => n20724, A2 => n19790, B1 => n20718, B2 => 
                           n19791, ZN => n18504);
   U16985 : AOI22_X1 port map( A1 => n20724, A2 => n19770, B1 => n20718, B2 => 
                           n19771, ZN => n18486);
   U16986 : AOI22_X1 port map( A1 => n20724, A2 => n19750, B1 => n20718, B2 => 
                           n19751, ZN => n18468);
   U16987 : AOI22_X1 port map( A1 => n20724, A2 => n19730, B1 => n20718, B2 => 
                           n19731, ZN => n18450);
   U16988 : AOI22_X1 port map( A1 => n20724, A2 => n19710, B1 => n20718, B2 => 
                           n19711, ZN => n18432);
   U16989 : AOI22_X1 port map( A1 => n20724, A2 => n19690, B1 => n20718, B2 => 
                           n19691, ZN => n18414);
   U16990 : AOI22_X1 port map( A1 => n20724, A2 => n19670, B1 => n20718, B2 => 
                           n19671, ZN => n18396);
   U16991 : AOI22_X1 port map( A1 => n20724, A2 => n19650, B1 => n20718, B2 => 
                           n19651, ZN => n18378);
   U16992 : AOI22_X1 port map( A1 => n20724, A2 => n19630, B1 => n20718, B2 => 
                           n19631, ZN => n18360);
   U16993 : AOI22_X1 port map( A1 => n20724, A2 => n19610, B1 => n20718, B2 => 
                           n19611, ZN => n18342);
   U16994 : AOI22_X1 port map( A1 => n20724, A2 => n19590, B1 => n20718, B2 => 
                           n19591, ZN => n18324);
   U16995 : AOI22_X1 port map( A1 => n20725, A2 => n19570, B1 => n20719, B2 => 
                           n19571, ZN => n18306);
   U16996 : AOI22_X1 port map( A1 => n20725, A2 => n19550, B1 => n20719, B2 => 
                           n19551, ZN => n18288);
   U16997 : AOI22_X1 port map( A1 => n20725, A2 => n19530, B1 => n20719, B2 => 
                           n19531, ZN => n18270);
   U16998 : AOI22_X1 port map( A1 => n20725, A2 => n19510, B1 => n20719, B2 => 
                           n19511, ZN => n18252);
   U16999 : AOI22_X1 port map( A1 => n20725, A2 => n19490, B1 => n20719, B2 => 
                           n19491, ZN => n18234);
   U17000 : AOI22_X1 port map( A1 => n20725, A2 => n19470, B1 => n20719, B2 => 
                           n19471, ZN => n18216);
   U17001 : AOI22_X1 port map( A1 => n20725, A2 => n19450, B1 => n20719, B2 => 
                           n19451, ZN => n18198);
   U17002 : AOI22_X1 port map( A1 => n20725, A2 => n19430, B1 => n20719, B2 => 
                           n19431, ZN => n18180);
   U17003 : AOI22_X1 port map( A1 => n20725, A2 => n19410, B1 => n20719, B2 => 
                           n19411, ZN => n18162);
   U17004 : AOI22_X1 port map( A1 => n20725, A2 => n19390, B1 => n20719, B2 => 
                           n19391, ZN => n18144);
   U17005 : AOI22_X1 port map( A1 => n20725, A2 => n19370, B1 => n20719, B2 => 
                           n19371, ZN => n18126);
   U17006 : AOI22_X1 port map( A1 => n20725, A2 => n19350, B1 => n20719, B2 => 
                           n19351, ZN => n18108);
   U17007 : AOI22_X1 port map( A1 => n20726, A2 => n19330, B1 => n20720, B2 => 
                           n19331, ZN => n18090);
   U17008 : AOI22_X1 port map( A1 => n20726, A2 => n19310, B1 => n20720, B2 => 
                           n19311, ZN => n18072);
   U17009 : AOI22_X1 port map( A1 => n20726, A2 => n19290, B1 => n20720, B2 => 
                           n19291, ZN => n18054);
   U17010 : AOI22_X1 port map( A1 => n20726, A2 => n19270, B1 => n20720, B2 => 
                           n19271, ZN => n18036);
   U17011 : AOI22_X1 port map( A1 => n20726, A2 => n19250, B1 => n20720, B2 => 
                           n19251, ZN => n18018);
   U17012 : AOI22_X1 port map( A1 => n20726, A2 => n19230, B1 => n20720, B2 => 
                           n19231, ZN => n18000);
   U17013 : AOI22_X1 port map( A1 => n20726, A2 => n19210, B1 => n20720, B2 => 
                           n19211, ZN => n17982);
   U17014 : AOI22_X1 port map( A1 => n20726, A2 => n19190, B1 => n20720, B2 => 
                           n19191, ZN => n17964);
   U17015 : AOI22_X1 port map( A1 => n20726, A2 => n19170, B1 => n20720, B2 => 
                           n19171, ZN => n17946);
   U17016 : AOI22_X1 port map( A1 => n20726, A2 => n19150, B1 => n20720, B2 => 
                           n19151, ZN => n17928);
   U17017 : AOI22_X1 port map( A1 => n20726, A2 => n19130, B1 => n20720, B2 => 
                           n19131, ZN => n17910);
   U17018 : AOI22_X1 port map( A1 => n20726, A2 => n19110, B1 => n20720, B2 => 
                           n19111, ZN => n17892);
   U17019 : AOI22_X1 port map( A1 => n20727, A2 => n19090, B1 => n20721, B2 => 
                           n19091, ZN => n17874);
   U17020 : AOI22_X1 port map( A1 => n20727, A2 => n19070, B1 => n20721, B2 => 
                           n19071, ZN => n17856);
   U17021 : AOI22_X1 port map( A1 => n20727, A2 => n19050, B1 => n20721, B2 => 
                           n19051, ZN => n17838);
   U17022 : AOI22_X1 port map( A1 => n20727, A2 => n19030, B1 => n20721, B2 => 
                           n19031, ZN => n17820);
   U17023 : AOI22_X1 port map( A1 => n20727, A2 => n19010, B1 => n20721, B2 => 
                           n19011, ZN => n17802);
   U17024 : AOI22_X1 port map( A1 => n20727, A2 => n18990, B1 => n20721, B2 => 
                           n18991, ZN => n17784);
   U17025 : AOI22_X1 port map( A1 => n20727, A2 => n18970, B1 => n20721, B2 => 
                           n18971, ZN => n17766);
   U17026 : AOI22_X1 port map( A1 => n20727, A2 => n18950, B1 => n20721, B2 => 
                           n18951, ZN => n17748);
   U17027 : AOI22_X1 port map( A1 => n20727, A2 => n18930, B1 => n20721, B2 => 
                           n18931, ZN => n17730);
   U17028 : AOI22_X1 port map( A1 => n20727, A2 => n18910, B1 => n20721, B2 => 
                           n18911, ZN => n17712);
   U17029 : AOI22_X1 port map( A1 => n20727, A2 => n18890, B1 => n20721, B2 => 
                           n18891, ZN => n17694);
   U17030 : AOI22_X1 port map( A1 => n20727, A2 => n18870, B1 => n20721, B2 => 
                           n18871, ZN => n17676);
   U17031 : AOI22_X1 port map( A1 => n20728, A2 => n18850, B1 => n20722, B2 => 
                           n18851, ZN => n17658);
   U17032 : AOI22_X1 port map( A1 => n20728, A2 => n18830, B1 => n20722, B2 => 
                           n18831, ZN => n17640);
   U17033 : AOI22_X1 port map( A1 => n20728, A2 => n18810, B1 => n20722, B2 => 
                           n18811, ZN => n17622);
   U17034 : AOI22_X1 port map( A1 => n20728, A2 => n18790, B1 => n20722, B2 => 
                           n18791, ZN => n17604);
   U17035 : AOI22_X1 port map( A1 => n20728, A2 => n18770, B1 => n20722, B2 => 
                           n18771, ZN => n17586);
   U17036 : AOI22_X1 port map( A1 => n20728, A2 => n18750, B1 => n20722, B2 => 
                           n18751, ZN => n17568);
   U17037 : AOI22_X1 port map( A1 => n20728, A2 => n18730, B1 => n20722, B2 => 
                           n18731, ZN => n17550);
   U17038 : AOI22_X1 port map( A1 => n20728, A2 => n18710, B1 => n20722, B2 => 
                           n18711, ZN => n17532);
   U17039 : AOI22_X1 port map( A1 => n20728, A2 => n18690, B1 => n20722, B2 => 
                           n18691, ZN => n17514);
   U17040 : AOI22_X1 port map( A1 => n20728, A2 => n18670, B1 => n20722, B2 => 
                           n18671, ZN => n17496);
   U17041 : AOI22_X1 port map( A1 => n20728, A2 => n18650, B1 => n20722, B2 => 
                           n18651, ZN => n17478);
   U17042 : AOI22_X1 port map( A1 => n20728, A2 => n18630, B1 => n20722, B2 => 
                           n18631, ZN => n17460);
   U17043 : AOI22_X1 port map( A1 => n20729, A2 => n18610, B1 => n20723, B2 => 
                           n18611, ZN => n17442);
   U17044 : AOI22_X1 port map( A1 => n20729, A2 => n18590, B1 => n20723, B2 => 
                           n18591, ZN => n17424);
   U17045 : AOI22_X1 port map( A1 => n20729, A2 => n18570, B1 => n20723, B2 => 
                           n18571, ZN => n17406);
   U17046 : AOI22_X1 port map( A1 => n20729, A2 => n18550, B1 => n20723, B2 => 
                           n18551, ZN => n17386);
   U17047 : AOI22_X1 port map( A1 => n20916, A2 => n19810, B1 => n20910, B2 => 
                           n19811, ZN => n17336);
   U17048 : AOI22_X1 port map( A1 => n20916, A2 => n19790, B1 => n20910, B2 => 
                           n19791, ZN => n17301);
   U17049 : AOI22_X1 port map( A1 => n20916, A2 => n19770, B1 => n20910, B2 => 
                           n19771, ZN => n17282);
   U17050 : AOI22_X1 port map( A1 => n20916, A2 => n19750, B1 => n20910, B2 => 
                           n19751, ZN => n17263);
   U17051 : AOI22_X1 port map( A1 => n20916, A2 => n19730, B1 => n20910, B2 => 
                           n19731, ZN => n17244);
   U17052 : AOI22_X1 port map( A1 => n20916, A2 => n19710, B1 => n20910, B2 => 
                           n19711, ZN => n17225);
   U17053 : AOI22_X1 port map( A1 => n20916, A2 => n19690, B1 => n20910, B2 => 
                           n19691, ZN => n17206);
   U17054 : AOI22_X1 port map( A1 => n20916, A2 => n19670, B1 => n20910, B2 => 
                           n19671, ZN => n17187);
   U17055 : AOI22_X1 port map( A1 => n20916, A2 => n19650, B1 => n20910, B2 => 
                           n19651, ZN => n17168);
   U17056 : AOI22_X1 port map( A1 => n20916, A2 => n19630, B1 => n20910, B2 => 
                           n19631, ZN => n17149);
   U17057 : AOI22_X1 port map( A1 => n20916, A2 => n19610, B1 => n20910, B2 => 
                           n19611, ZN => n17130);
   U17058 : AOI22_X1 port map( A1 => n20916, A2 => n19590, B1 => n20910, B2 => 
                           n19591, ZN => n17111);
   U17059 : AOI22_X1 port map( A1 => n20917, A2 => n19570, B1 => n20911, B2 => 
                           n19571, ZN => n17092);
   U17060 : AOI22_X1 port map( A1 => n20917, A2 => n19550, B1 => n20911, B2 => 
                           n19551, ZN => n17073);
   U17061 : AOI22_X1 port map( A1 => n20917, A2 => n19530, B1 => n20911, B2 => 
                           n19531, ZN => n17054);
   U17062 : AOI22_X1 port map( A1 => n20917, A2 => n19510, B1 => n20911, B2 => 
                           n19511, ZN => n17035);
   U17063 : AOI22_X1 port map( A1 => n20917, A2 => n19490, B1 => n20911, B2 => 
                           n19491, ZN => n17016);
   U17064 : AOI22_X1 port map( A1 => n20917, A2 => n19470, B1 => n20911, B2 => 
                           n19471, ZN => n16997);
   U17065 : AOI22_X1 port map( A1 => n20917, A2 => n19450, B1 => n20911, B2 => 
                           n19451, ZN => n16978);
   U17066 : AOI22_X1 port map( A1 => n20917, A2 => n19430, B1 => n20911, B2 => 
                           n19431, ZN => n16959);
   U17067 : AOI22_X1 port map( A1 => n20917, A2 => n19410, B1 => n20911, B2 => 
                           n19411, ZN => n16940);
   U17068 : AOI22_X1 port map( A1 => n20917, A2 => n19390, B1 => n20911, B2 => 
                           n19391, ZN => n16921);
   U17069 : AOI22_X1 port map( A1 => n20917, A2 => n19370, B1 => n20911, B2 => 
                           n19371, ZN => n16902);
   U17070 : AOI22_X1 port map( A1 => n20917, A2 => n19350, B1 => n20911, B2 => 
                           n19351, ZN => n16883);
   U17071 : AOI22_X1 port map( A1 => n20918, A2 => n19330, B1 => n20912, B2 => 
                           n19331, ZN => n16864);
   U17072 : AOI22_X1 port map( A1 => n20918, A2 => n19310, B1 => n20912, B2 => 
                           n19311, ZN => n16845);
   U17073 : AOI22_X1 port map( A1 => n20918, A2 => n19290, B1 => n20912, B2 => 
                           n19291, ZN => n16826);
   U17074 : AOI22_X1 port map( A1 => n20918, A2 => n19270, B1 => n20912, B2 => 
                           n19271, ZN => n16807);
   U17075 : AOI22_X1 port map( A1 => n20918, A2 => n19250, B1 => n20912, B2 => 
                           n19251, ZN => n16788);
   U17076 : AOI22_X1 port map( A1 => n20918, A2 => n19230, B1 => n20912, B2 => 
                           n19231, ZN => n16769);
   U17077 : AOI22_X1 port map( A1 => n20918, A2 => n19210, B1 => n20912, B2 => 
                           n19211, ZN => n16750);
   U17078 : AOI22_X1 port map( A1 => n20918, A2 => n19190, B1 => n20912, B2 => 
                           n19191, ZN => n16731);
   U17079 : AOI22_X1 port map( A1 => n20918, A2 => n19170, B1 => n20912, B2 => 
                           n19171, ZN => n16712);
   U17080 : AOI22_X1 port map( A1 => n20918, A2 => n19150, B1 => n20912, B2 => 
                           n19151, ZN => n16693);
   U17081 : AOI22_X1 port map( A1 => n20918, A2 => n19130, B1 => n20912, B2 => 
                           n19131, ZN => n16674);
   U17082 : AOI22_X1 port map( A1 => n20918, A2 => n19110, B1 => n20912, B2 => 
                           n19111, ZN => n16655);
   U17083 : AOI22_X1 port map( A1 => n20919, A2 => n19090, B1 => n20913, B2 => 
                           n19091, ZN => n16636);
   U17084 : AOI22_X1 port map( A1 => n20919, A2 => n19070, B1 => n20913, B2 => 
                           n19071, ZN => n16617);
   U17085 : AOI22_X1 port map( A1 => n20919, A2 => n19050, B1 => n20913, B2 => 
                           n19051, ZN => n16598);
   U17086 : AOI22_X1 port map( A1 => n20919, A2 => n19030, B1 => n20913, B2 => 
                           n19031, ZN => n16579);
   U17087 : AOI22_X1 port map( A1 => n20919, A2 => n19010, B1 => n20913, B2 => 
                           n19011, ZN => n16560);
   U17088 : AOI22_X1 port map( A1 => n20919, A2 => n18990, B1 => n20913, B2 => 
                           n18991, ZN => n16541);
   U17089 : AOI22_X1 port map( A1 => n20919, A2 => n18970, B1 => n20913, B2 => 
                           n18971, ZN => n16522);
   U17090 : AOI22_X1 port map( A1 => n20919, A2 => n18950, B1 => n20913, B2 => 
                           n18951, ZN => n16503);
   U17091 : AOI22_X1 port map( A1 => n20919, A2 => n18930, B1 => n20913, B2 => 
                           n18931, ZN => n16484);
   U17092 : AOI22_X1 port map( A1 => n20919, A2 => n18910, B1 => n20913, B2 => 
                           n18911, ZN => n16465);
   U17093 : AOI22_X1 port map( A1 => n20919, A2 => n18890, B1 => n20913, B2 => 
                           n18891, ZN => n16446);
   U17094 : AOI22_X1 port map( A1 => n20919, A2 => n18870, B1 => n20913, B2 => 
                           n18871, ZN => n16427);
   U17095 : AOI22_X1 port map( A1 => n20920, A2 => n18850, B1 => n20914, B2 => 
                           n18851, ZN => n16408);
   U17096 : AOI22_X1 port map( A1 => n20920, A2 => n18830, B1 => n20914, B2 => 
                           n18831, ZN => n16389);
   U17097 : AOI22_X1 port map( A1 => n20920, A2 => n18810, B1 => n20914, B2 => 
                           n18811, ZN => n16370);
   U17098 : AOI22_X1 port map( A1 => n20920, A2 => n18790, B1 => n20914, B2 => 
                           n18791, ZN => n16351);
   U17099 : AOI22_X1 port map( A1 => n20920, A2 => n18770, B1 => n20914, B2 => 
                           n18771, ZN => n16332);
   U17100 : AOI22_X1 port map( A1 => n20920, A2 => n18750, B1 => n20914, B2 => 
                           n18751, ZN => n16313);
   U17101 : AOI22_X1 port map( A1 => n20920, A2 => n18730, B1 => n20914, B2 => 
                           n18731, ZN => n16294);
   U17102 : AOI22_X1 port map( A1 => n20920, A2 => n18710, B1 => n20914, B2 => 
                           n18711, ZN => n16275);
   U17103 : AOI22_X1 port map( A1 => n20920, A2 => n18690, B1 => n20914, B2 => 
                           n18691, ZN => n16256);
   U17104 : AOI22_X1 port map( A1 => n20920, A2 => n18670, B1 => n20914, B2 => 
                           n18671, ZN => n16237);
   U17105 : AOI22_X1 port map( A1 => n20920, A2 => n18650, B1 => n20914, B2 => 
                           n18651, ZN => n16218);
   U17106 : AOI22_X1 port map( A1 => n20920, A2 => n18630, B1 => n20914, B2 => 
                           n18631, ZN => n16199);
   U17107 : AOI22_X1 port map( A1 => n20921, A2 => n18610, B1 => n20915, B2 => 
                           n18611, ZN => n16180);
   U17108 : AOI22_X1 port map( A1 => n20921, A2 => n18590, B1 => n20915, B2 => 
                           n18591, ZN => n16161);
   U17109 : AOI22_X1 port map( A1 => n20921, A2 => n18570, B1 => n20915, B2 => 
                           n18571, ZN => n16142);
   U17110 : AOI22_X1 port map( A1 => n20921, A2 => n18550, B1 => n20915, B2 => 
                           n18551, ZN => n16121);
   U17111 : OAI221_X1 port map( B1 => n14404, B2 => n20904, C1 => n14872, C2 =>
                           n20898, A => n18511, ZN => n18510);
   U17112 : AOI22_X1 port map( A1 => n20892, A2 => n19808, B1 => n20886, B2 => 
                           n19809, ZN => n18511);
   U17113 : OAI221_X1 port map( B1 => n17302, B2 => n20880, C1 => n14337, C2 =>
                           n20874, A => n18518, ZN => n18509);
   U17114 : AOI22_X1 port map( A1 => n20868, A2 => n9212, B1 => n20862, B2 => 
                           n8828, ZN => n18518);
   U17115 : OAI221_X1 port map( B1 => n14271, B2 => n20760, C1 => n15337, C2 =>
                           n20754, A => n18536, ZN => n18527);
   U17116 : AOI22_X1 port map( A1 => n20748, A2 => n19814, B1 => n20742, B2 => 
                           n19815, ZN => n18536);
   U17117 : OAI221_X1 port map( B1 => n15804, B2 => n20784, C1 => n14806, C2 =>
                           n20778, A => n18533, ZN => n18528);
   U17118 : AOI22_X1 port map( A1 => n20772, A2 => n8955, B1 => n20766, B2 => 
                           n19819, ZN => n18533);
   U17119 : OAI221_X1 port map( B1 => n14403, B2 => n20904, C1 => n14871, C2 =>
                           n20898, A => n18493, ZN => n18492);
   U17120 : AOI22_X1 port map( A1 => n20892, A2 => n19788, B1 => n20886, B2 => 
                           n19789, ZN => n18493);
   U17121 : OAI221_X1 port map( B1 => n17283, B2 => n20880, C1 => n14336, C2 =>
                           n20874, A => n18494, ZN => n18491);
   U17122 : AOI22_X1 port map( A1 => n20868, A2 => n9208, B1 => n20862, B2 => 
                           n8824, ZN => n18494);
   U17123 : OAI221_X1 port map( B1 => n14270, B2 => n20760, C1 => n15336, C2 =>
                           n20754, A => n18503, ZN => n18498);
   U17124 : AOI22_X1 port map( A1 => n20748, A2 => n19794, B1 => n20742, B2 => 
                           n19795, ZN => n18503);
   U17125 : OAI221_X1 port map( B1 => n15803, B2 => n20784, C1 => n14805, C2 =>
                           n20778, A => n18502, ZN => n18499);
   U17126 : AOI22_X1 port map( A1 => n20772, A2 => n8953, B1 => n20766, B2 => 
                           n19799, ZN => n18502);
   U17127 : OAI221_X1 port map( B1 => n14402, B2 => n20904, C1 => n14870, C2 =>
                           n20898, A => n18475, ZN => n18474);
   U17128 : AOI22_X1 port map( A1 => n20892, A2 => n19768, B1 => n20886, B2 => 
                           n19769, ZN => n18475);
   U17129 : OAI221_X1 port map( B1 => n17264, B2 => n20880, C1 => n14335, C2 =>
                           n20874, A => n18476, ZN => n18473);
   U17130 : AOI22_X1 port map( A1 => n20868, A2 => n9204, B1 => n20862, B2 => 
                           n8820, ZN => n18476);
   U17131 : OAI221_X1 port map( B1 => n14269, B2 => n20760, C1 => n15335, C2 =>
                           n20754, A => n18485, ZN => n18480);
   U17132 : AOI22_X1 port map( A1 => n20748, A2 => n19774, B1 => n20742, B2 => 
                           n19775, ZN => n18485);
   U17133 : OAI221_X1 port map( B1 => n15802, B2 => n20784, C1 => n14804, C2 =>
                           n20778, A => n18484, ZN => n18481);
   U17134 : AOI22_X1 port map( A1 => n20772, A2 => n8951, B1 => n20766, B2 => 
                           n19779, ZN => n18484);
   U17135 : OAI221_X1 port map( B1 => n14401, B2 => n20904, C1 => n14869, C2 =>
                           n20898, A => n18457, ZN => n18456);
   U17136 : AOI22_X1 port map( A1 => n20892, A2 => n19748, B1 => n20886, B2 => 
                           n19749, ZN => n18457);
   U17137 : OAI221_X1 port map( B1 => n17245, B2 => n20880, C1 => n14334, C2 =>
                           n20874, A => n18458, ZN => n18455);
   U17138 : AOI22_X1 port map( A1 => n20868, A2 => n9200, B1 => n20862, B2 => 
                           n8816, ZN => n18458);
   U17139 : OAI221_X1 port map( B1 => n14268, B2 => n20760, C1 => n15334, C2 =>
                           n20754, A => n18467, ZN => n18462);
   U17140 : AOI22_X1 port map( A1 => n20748, A2 => n19754, B1 => n20742, B2 => 
                           n19755, ZN => n18467);
   U17141 : OAI221_X1 port map( B1 => n15801, B2 => n20784, C1 => n14803, C2 =>
                           n20778, A => n18466, ZN => n18463);
   U17142 : AOI22_X1 port map( A1 => n20772, A2 => n8949, B1 => n20766, B2 => 
                           n19759, ZN => n18466);
   U17143 : OAI221_X1 port map( B1 => n14400, B2 => n20904, C1 => n14868, C2 =>
                           n20898, A => n18439, ZN => n18438);
   U17144 : AOI22_X1 port map( A1 => n20892, A2 => n19728, B1 => n20886, B2 => 
                           n19729, ZN => n18439);
   U17145 : OAI221_X1 port map( B1 => n17226, B2 => n20880, C1 => n14333, C2 =>
                           n20874, A => n18440, ZN => n18437);
   U17146 : AOI22_X1 port map( A1 => n20868, A2 => n9196, B1 => n20862, B2 => 
                           n8812, ZN => n18440);
   U17147 : OAI221_X1 port map( B1 => n14267, B2 => n20760, C1 => n15333, C2 =>
                           n20754, A => n18449, ZN => n18444);
   U17148 : AOI22_X1 port map( A1 => n20748, A2 => n19734, B1 => n20742, B2 => 
                           n19735, ZN => n18449);
   U17149 : OAI221_X1 port map( B1 => n15800, B2 => n20784, C1 => n14802, C2 =>
                           n20778, A => n18448, ZN => n18445);
   U17150 : AOI22_X1 port map( A1 => n20772, A2 => n8947, B1 => n20766, B2 => 
                           n19739, ZN => n18448);
   U17151 : OAI221_X1 port map( B1 => n14399, B2 => n20904, C1 => n14867, C2 =>
                           n20898, A => n18421, ZN => n18420);
   U17152 : AOI22_X1 port map( A1 => n20892, A2 => n19708, B1 => n20886, B2 => 
                           n19709, ZN => n18421);
   U17153 : OAI221_X1 port map( B1 => n17207, B2 => n20880, C1 => n14332, C2 =>
                           n20874, A => n18422, ZN => n18419);
   U17154 : AOI22_X1 port map( A1 => n20868, A2 => n9192, B1 => n20862, B2 => 
                           n8808, ZN => n18422);
   U17155 : OAI221_X1 port map( B1 => n14266, B2 => n20760, C1 => n15332, C2 =>
                           n20754, A => n18431, ZN => n18426);
   U17156 : AOI22_X1 port map( A1 => n20748, A2 => n19714, B1 => n20742, B2 => 
                           n19715, ZN => n18431);
   U17157 : OAI221_X1 port map( B1 => n15799, B2 => n20784, C1 => n14801, C2 =>
                           n20778, A => n18430, ZN => n18427);
   U17158 : AOI22_X1 port map( A1 => n20772, A2 => n8945, B1 => n20766, B2 => 
                           n19719, ZN => n18430);
   U17159 : OAI221_X1 port map( B1 => n14398, B2 => n20904, C1 => n14866, C2 =>
                           n20898, A => n18403, ZN => n18402);
   U17160 : AOI22_X1 port map( A1 => n20892, A2 => n19688, B1 => n20886, B2 => 
                           n19689, ZN => n18403);
   U17161 : OAI221_X1 port map( B1 => n17188, B2 => n20880, C1 => n14331, C2 =>
                           n20874, A => n18404, ZN => n18401);
   U17162 : AOI22_X1 port map( A1 => n20868, A2 => n9188, B1 => n20862, B2 => 
                           n8804, ZN => n18404);
   U17163 : OAI221_X1 port map( B1 => n14265, B2 => n20760, C1 => n15331, C2 =>
                           n20754, A => n18413, ZN => n18408);
   U17164 : AOI22_X1 port map( A1 => n20748, A2 => n19694, B1 => n20742, B2 => 
                           n19695, ZN => n18413);
   U17165 : OAI221_X1 port map( B1 => n15798, B2 => n20784, C1 => n14800, C2 =>
                           n20778, A => n18412, ZN => n18409);
   U17166 : AOI22_X1 port map( A1 => n20772, A2 => n8943, B1 => n20766, B2 => 
                           n19699, ZN => n18412);
   U17167 : OAI221_X1 port map( B1 => n14397, B2 => n20904, C1 => n14865, C2 =>
                           n20898, A => n18385, ZN => n18384);
   U17168 : AOI22_X1 port map( A1 => n20892, A2 => n19668, B1 => n20886, B2 => 
                           n19669, ZN => n18385);
   U17169 : OAI221_X1 port map( B1 => n17169, B2 => n20880, C1 => n14330, C2 =>
                           n20874, A => n18386, ZN => n18383);
   U17170 : AOI22_X1 port map( A1 => n20868, A2 => n9184, B1 => n20862, B2 => 
                           n8800, ZN => n18386);
   U17171 : OAI221_X1 port map( B1 => n14264, B2 => n20760, C1 => n15330, C2 =>
                           n20754, A => n18395, ZN => n18390);
   U17172 : AOI22_X1 port map( A1 => n20748, A2 => n19674, B1 => n20742, B2 => 
                           n19675, ZN => n18395);
   U17173 : OAI221_X1 port map( B1 => n15797, B2 => n20784, C1 => n14799, C2 =>
                           n20778, A => n18394, ZN => n18391);
   U17174 : AOI22_X1 port map( A1 => n20772, A2 => n8941, B1 => n20766, B2 => 
                           n19679, ZN => n18394);
   U17175 : OAI221_X1 port map( B1 => n14396, B2 => n20904, C1 => n14864, C2 =>
                           n20898, A => n18367, ZN => n18366);
   U17176 : AOI22_X1 port map( A1 => n20892, A2 => n19648, B1 => n20886, B2 => 
                           n19649, ZN => n18367);
   U17177 : OAI221_X1 port map( B1 => n17150, B2 => n20880, C1 => n14329, C2 =>
                           n20874, A => n18368, ZN => n18365);
   U17178 : AOI22_X1 port map( A1 => n20868, A2 => n9180, B1 => n20862, B2 => 
                           n8796, ZN => n18368);
   U17179 : OAI221_X1 port map( B1 => n14263, B2 => n20760, C1 => n15329, C2 =>
                           n20754, A => n18377, ZN => n18372);
   U17180 : AOI22_X1 port map( A1 => n20748, A2 => n19654, B1 => n20742, B2 => 
                           n19655, ZN => n18377);
   U17181 : OAI221_X1 port map( B1 => n15796, B2 => n20784, C1 => n14798, C2 =>
                           n20778, A => n18376, ZN => n18373);
   U17182 : AOI22_X1 port map( A1 => n20772, A2 => n8939, B1 => n20766, B2 => 
                           n19659, ZN => n18376);
   U17183 : OAI221_X1 port map( B1 => n14395, B2 => n20904, C1 => n14863, C2 =>
                           n20898, A => n18349, ZN => n18348);
   U17184 : AOI22_X1 port map( A1 => n20892, A2 => n19628, B1 => n20886, B2 => 
                           n19629, ZN => n18349);
   U17185 : OAI221_X1 port map( B1 => n17131, B2 => n20880, C1 => n14328, C2 =>
                           n20874, A => n18350, ZN => n18347);
   U17186 : AOI22_X1 port map( A1 => n20868, A2 => n9176, B1 => n20862, B2 => 
                           n8792, ZN => n18350);
   U17187 : OAI221_X1 port map( B1 => n14262, B2 => n20760, C1 => n15328, C2 =>
                           n20754, A => n18359, ZN => n18354);
   U17188 : AOI22_X1 port map( A1 => n20748, A2 => n19634, B1 => n20742, B2 => 
                           n19635, ZN => n18359);
   U17189 : OAI221_X1 port map( B1 => n15795, B2 => n20784, C1 => n14797, C2 =>
                           n20778, A => n18358, ZN => n18355);
   U17190 : AOI22_X1 port map( A1 => n20772, A2 => n8937, B1 => n20766, B2 => 
                           n19639, ZN => n18358);
   U17191 : OAI221_X1 port map( B1 => n14394, B2 => n20904, C1 => n14862, C2 =>
                           n20898, A => n18331, ZN => n18330);
   U17192 : AOI22_X1 port map( A1 => n20892, A2 => n19608, B1 => n20886, B2 => 
                           n19609, ZN => n18331);
   U17193 : OAI221_X1 port map( B1 => n17112, B2 => n20880, C1 => n14327, C2 =>
                           n20874, A => n18332, ZN => n18329);
   U17194 : AOI22_X1 port map( A1 => n20868, A2 => n9172, B1 => n20862, B2 => 
                           n8788, ZN => n18332);
   U17195 : OAI221_X1 port map( B1 => n14261, B2 => n20760, C1 => n15327, C2 =>
                           n20754, A => n18341, ZN => n18336);
   U17196 : AOI22_X1 port map( A1 => n20748, A2 => n19614, B1 => n20742, B2 => 
                           n19615, ZN => n18341);
   U17197 : OAI221_X1 port map( B1 => n15794, B2 => n20784, C1 => n14796, C2 =>
                           n20778, A => n18340, ZN => n18337);
   U17198 : AOI22_X1 port map( A1 => n20772, A2 => n8935, B1 => n20766, B2 => 
                           n19619, ZN => n18340);
   U17199 : OAI221_X1 port map( B1 => n14393, B2 => n20904, C1 => n14861, C2 =>
                           n20898, A => n18313, ZN => n18312);
   U17200 : AOI22_X1 port map( A1 => n20892, A2 => n19588, B1 => n20886, B2 => 
                           n19589, ZN => n18313);
   U17201 : OAI221_X1 port map( B1 => n17093, B2 => n20880, C1 => n14326, C2 =>
                           n20874, A => n18314, ZN => n18311);
   U17202 : AOI22_X1 port map( A1 => n20868, A2 => n9168, B1 => n20862, B2 => 
                           n8784, ZN => n18314);
   U17203 : OAI221_X1 port map( B1 => n14260, B2 => n20760, C1 => n15326, C2 =>
                           n20754, A => n18323, ZN => n18318);
   U17204 : AOI22_X1 port map( A1 => n20748, A2 => n19594, B1 => n20742, B2 => 
                           n19595, ZN => n18323);
   U17205 : OAI221_X1 port map( B1 => n15793, B2 => n20784, C1 => n14795, C2 =>
                           n20778, A => n18322, ZN => n18319);
   U17206 : AOI22_X1 port map( A1 => n20772, A2 => n8933, B1 => n20766, B2 => 
                           n19599, ZN => n18322);
   U17207 : OAI221_X1 port map( B1 => n14392, B2 => n20905, C1 => n14860, C2 =>
                           n20899, A => n18295, ZN => n18294);
   U17208 : AOI22_X1 port map( A1 => n20893, A2 => n19568, B1 => n20887, B2 => 
                           n19569, ZN => n18295);
   U17209 : OAI221_X1 port map( B1 => n15792, B2 => n20785, C1 => n14794, C2 =>
                           n20779, A => n18304, ZN => n18301);
   U17210 : AOI22_X1 port map( A1 => n20773, A2 => n8931, B1 => n20767, B2 => 
                           n19579, ZN => n18304);
   U17211 : OAI221_X1 port map( B1 => n14391, B2 => n20905, C1 => n14859, C2 =>
                           n20899, A => n18277, ZN => n18276);
   U17212 : AOI22_X1 port map( A1 => n20893, A2 => n19548, B1 => n20887, B2 => 
                           n19549, ZN => n18277);
   U17213 : OAI221_X1 port map( B1 => n15791, B2 => n20785, C1 => n14793, C2 =>
                           n20779, A => n18286, ZN => n18283);
   U17214 : AOI22_X1 port map( A1 => n20773, A2 => n8929, B1 => n20767, B2 => 
                           n19559, ZN => n18286);
   U17215 : OAI221_X1 port map( B1 => n14390, B2 => n20905, C1 => n14858, C2 =>
                           n20899, A => n18259, ZN => n18258);
   U17216 : AOI22_X1 port map( A1 => n20893, A2 => n19528, B1 => n20887, B2 => 
                           n19529, ZN => n18259);
   U17217 : OAI221_X1 port map( B1 => n15790, B2 => n20785, C1 => n14792, C2 =>
                           n20779, A => n18268, ZN => n18265);
   U17218 : AOI22_X1 port map( A1 => n20773, A2 => n8927, B1 => n20767, B2 => 
                           n19539, ZN => n18268);
   U17219 : OAI221_X1 port map( B1 => n14389, B2 => n20905, C1 => n14857, C2 =>
                           n20899, A => n18241, ZN => n18240);
   U17220 : AOI22_X1 port map( A1 => n20893, A2 => n19508, B1 => n20887, B2 => 
                           n19509, ZN => n18241);
   U17221 : OAI221_X1 port map( B1 => n15789, B2 => n20785, C1 => n14791, C2 =>
                           n20779, A => n18250, ZN => n18247);
   U17222 : AOI22_X1 port map( A1 => n20773, A2 => n8925, B1 => n20767, B2 => 
                           n19519, ZN => n18250);
   U17223 : OAI221_X1 port map( B1 => n14388, B2 => n20905, C1 => n14856, C2 =>
                           n20899, A => n18223, ZN => n18222);
   U17224 : AOI22_X1 port map( A1 => n20893, A2 => n19488, B1 => n20887, B2 => 
                           n19489, ZN => n18223);
   U17225 : OAI221_X1 port map( B1 => n15788, B2 => n20785, C1 => n14790, C2 =>
                           n20779, A => n18232, ZN => n18229);
   U17226 : AOI22_X1 port map( A1 => n20773, A2 => n8923, B1 => n20767, B2 => 
                           n19499, ZN => n18232);
   U17227 : OAI221_X1 port map( B1 => n14387, B2 => n20905, C1 => n14855, C2 =>
                           n20899, A => n18205, ZN => n18204);
   U17228 : AOI22_X1 port map( A1 => n20893, A2 => n19468, B1 => n20887, B2 => 
                           n19469, ZN => n18205);
   U17229 : OAI221_X1 port map( B1 => n15787, B2 => n20785, C1 => n14789, C2 =>
                           n20779, A => n18214, ZN => n18211);
   U17230 : AOI22_X1 port map( A1 => n20773, A2 => n8921, B1 => n20767, B2 => 
                           n19479, ZN => n18214);
   U17231 : OAI221_X1 port map( B1 => n14386, B2 => n20905, C1 => n14854, C2 =>
                           n20899, A => n18187, ZN => n18186);
   U17232 : AOI22_X1 port map( A1 => n20893, A2 => n19448, B1 => n20887, B2 => 
                           n19449, ZN => n18187);
   U17233 : OAI221_X1 port map( B1 => n15786, B2 => n20785, C1 => n14788, C2 =>
                           n20779, A => n18196, ZN => n18193);
   U17234 : AOI22_X1 port map( A1 => n20773, A2 => n8919, B1 => n20767, B2 => 
                           n19459, ZN => n18196);
   U17235 : OAI221_X1 port map( B1 => n14385, B2 => n20905, C1 => n14853, C2 =>
                           n20899, A => n18169, ZN => n18168);
   U17236 : AOI22_X1 port map( A1 => n20893, A2 => n19428, B1 => n20887, B2 => 
                           n19429, ZN => n18169);
   U17237 : OAI221_X1 port map( B1 => n15785, B2 => n20785, C1 => n14787, C2 =>
                           n20779, A => n18178, ZN => n18175);
   U17238 : AOI22_X1 port map( A1 => n20773, A2 => n8917, B1 => n20767, B2 => 
                           n19439, ZN => n18178);
   U17239 : OAI221_X1 port map( B1 => n14384, B2 => n20905, C1 => n14852, C2 =>
                           n20899, A => n18151, ZN => n18150);
   U17240 : AOI22_X1 port map( A1 => n20893, A2 => n19408, B1 => n20887, B2 => 
                           n19409, ZN => n18151);
   U17241 : OAI221_X1 port map( B1 => n15784, B2 => n20785, C1 => n14786, C2 =>
                           n20779, A => n18160, ZN => n18157);
   U17242 : AOI22_X1 port map( A1 => n20773, A2 => n8915, B1 => n20767, B2 => 
                           n19419, ZN => n18160);
   U17243 : OAI221_X1 port map( B1 => n14383, B2 => n20905, C1 => n14851, C2 =>
                           n20899, A => n18133, ZN => n18132);
   U17244 : AOI22_X1 port map( A1 => n20893, A2 => n19388, B1 => n20887, B2 => 
                           n19389, ZN => n18133);
   U17245 : OAI221_X1 port map( B1 => n15783, B2 => n20785, C1 => n14785, C2 =>
                           n20779, A => n18142, ZN => n18139);
   U17246 : AOI22_X1 port map( A1 => n20773, A2 => n8913, B1 => n20767, B2 => 
                           n19399, ZN => n18142);
   U17247 : OAI221_X1 port map( B1 => n14382, B2 => n20905, C1 => n14850, C2 =>
                           n20899, A => n18115, ZN => n18114);
   U17248 : AOI22_X1 port map( A1 => n20893, A2 => n19368, B1 => n20887, B2 => 
                           n19369, ZN => n18115);
   U17249 : OAI221_X1 port map( B1 => n15782, B2 => n20785, C1 => n14784, C2 =>
                           n20779, A => n18124, ZN => n18121);
   U17250 : AOI22_X1 port map( A1 => n20773, A2 => n8911, B1 => n20767, B2 => 
                           n19379, ZN => n18124);
   U17251 : OAI221_X1 port map( B1 => n14381, B2 => n20905, C1 => n14849, C2 =>
                           n20899, A => n18097, ZN => n18096);
   U17252 : AOI22_X1 port map( A1 => n20893, A2 => n19348, B1 => n20887, B2 => 
                           n19349, ZN => n18097);
   U17253 : OAI221_X1 port map( B1 => n15781, B2 => n20785, C1 => n14783, C2 =>
                           n20779, A => n18106, ZN => n18103);
   U17254 : AOI22_X1 port map( A1 => n20773, A2 => n8909, B1 => n20767, B2 => 
                           n19359, ZN => n18106);
   U17255 : OAI221_X1 port map( B1 => n14380, B2 => n20906, C1 => n14848, C2 =>
                           n20900, A => n18079, ZN => n18078);
   U17256 : AOI22_X1 port map( A1 => n20894, A2 => n19328, B1 => n20888, B2 => 
                           n19329, ZN => n18079);
   U17257 : OAI221_X1 port map( B1 => n15780, B2 => n20786, C1 => n14782, C2 =>
                           n20780, A => n18088, ZN => n18085);
   U17258 : AOI22_X1 port map( A1 => n20774, A2 => n8907, B1 => n20768, B2 => 
                           n19339, ZN => n18088);
   U17259 : OAI221_X1 port map( B1 => n14379, B2 => n20906, C1 => n14847, C2 =>
                           n20900, A => n18061, ZN => n18060);
   U17260 : AOI22_X1 port map( A1 => n20894, A2 => n19308, B1 => n20888, B2 => 
                           n19309, ZN => n18061);
   U17261 : OAI221_X1 port map( B1 => n15779, B2 => n20786, C1 => n14781, C2 =>
                           n20780, A => n18070, ZN => n18067);
   U17262 : AOI22_X1 port map( A1 => n20774, A2 => n8905, B1 => n20768, B2 => 
                           n19319, ZN => n18070);
   U17263 : OAI221_X1 port map( B1 => n14378, B2 => n20906, C1 => n14846, C2 =>
                           n20900, A => n18043, ZN => n18042);
   U17264 : AOI22_X1 port map( A1 => n20894, A2 => n19288, B1 => n20888, B2 => 
                           n19289, ZN => n18043);
   U17265 : OAI221_X1 port map( B1 => n15778, B2 => n20786, C1 => n14780, C2 =>
                           n20780, A => n18052, ZN => n18049);
   U17266 : AOI22_X1 port map( A1 => n20774, A2 => n8903, B1 => n20768, B2 => 
                           n19299, ZN => n18052);
   U17267 : OAI221_X1 port map( B1 => n14377, B2 => n20906, C1 => n14845, C2 =>
                           n20900, A => n18025, ZN => n18024);
   U17268 : AOI22_X1 port map( A1 => n20894, A2 => n19268, B1 => n20888, B2 => 
                           n19269, ZN => n18025);
   U17269 : OAI221_X1 port map( B1 => n15777, B2 => n20786, C1 => n14779, C2 =>
                           n20780, A => n18034, ZN => n18031);
   U17270 : AOI22_X1 port map( A1 => n20774, A2 => n8901, B1 => n20768, B2 => 
                           n19279, ZN => n18034);
   U17271 : OAI221_X1 port map( B1 => n14376, B2 => n20906, C1 => n14844, C2 =>
                           n20900, A => n18007, ZN => n18006);
   U17272 : AOI22_X1 port map( A1 => n20894, A2 => n19248, B1 => n20888, B2 => 
                           n19249, ZN => n18007);
   U17273 : OAI221_X1 port map( B1 => n15776, B2 => n20786, C1 => n14778, C2 =>
                           n20780, A => n18016, ZN => n18013);
   U17274 : AOI22_X1 port map( A1 => n20774, A2 => n8899, B1 => n20768, B2 => 
                           n19259, ZN => n18016);
   U17275 : OAI221_X1 port map( B1 => n14375, B2 => n20906, C1 => n14843, C2 =>
                           n20900, A => n17989, ZN => n17988);
   U17276 : AOI22_X1 port map( A1 => n20894, A2 => n19228, B1 => n20888, B2 => 
                           n19229, ZN => n17989);
   U17277 : OAI221_X1 port map( B1 => n15775, B2 => n20786, C1 => n14777, C2 =>
                           n20780, A => n17998, ZN => n17995);
   U17278 : AOI22_X1 port map( A1 => n20774, A2 => n8897, B1 => n20768, B2 => 
                           n19239, ZN => n17998);
   U17279 : OAI221_X1 port map( B1 => n14374, B2 => n20906, C1 => n14842, C2 =>
                           n20900, A => n17971, ZN => n17970);
   U17280 : AOI22_X1 port map( A1 => n20894, A2 => n19208, B1 => n20888, B2 => 
                           n19209, ZN => n17971);
   U17281 : OAI221_X1 port map( B1 => n15774, B2 => n20786, C1 => n14776, C2 =>
                           n20780, A => n17980, ZN => n17977);
   U17282 : AOI22_X1 port map( A1 => n20774, A2 => n8895, B1 => n20768, B2 => 
                           n19219, ZN => n17980);
   U17283 : OAI221_X1 port map( B1 => n14373, B2 => n20906, C1 => n14841, C2 =>
                           n20900, A => n17953, ZN => n17952);
   U17284 : AOI22_X1 port map( A1 => n20894, A2 => n19188, B1 => n20888, B2 => 
                           n19189, ZN => n17953);
   U17285 : OAI221_X1 port map( B1 => n15773, B2 => n20786, C1 => n14775, C2 =>
                           n20780, A => n17962, ZN => n17959);
   U17286 : AOI22_X1 port map( A1 => n20774, A2 => n8893, B1 => n20768, B2 => 
                           n19199, ZN => n17962);
   U17287 : OAI221_X1 port map( B1 => n14372, B2 => n20906, C1 => n14840, C2 =>
                           n20900, A => n17935, ZN => n17934);
   U17288 : AOI22_X1 port map( A1 => n20894, A2 => n19168, B1 => n20888, B2 => 
                           n19169, ZN => n17935);
   U17289 : OAI221_X1 port map( B1 => n15772, B2 => n20786, C1 => n14774, C2 =>
                           n20780, A => n17944, ZN => n17941);
   U17290 : AOI22_X1 port map( A1 => n20774, A2 => n8891, B1 => n20768, B2 => 
                           n19179, ZN => n17944);
   U17291 : OAI221_X1 port map( B1 => n14371, B2 => n20906, C1 => n14839, C2 =>
                           n20900, A => n17917, ZN => n17916);
   U17292 : AOI22_X1 port map( A1 => n20894, A2 => n19148, B1 => n20888, B2 => 
                           n19149, ZN => n17917);
   U17293 : OAI221_X1 port map( B1 => n15771, B2 => n20786, C1 => n14773, C2 =>
                           n20780, A => n17926, ZN => n17923);
   U17294 : AOI22_X1 port map( A1 => n20774, A2 => n8889, B1 => n20768, B2 => 
                           n19159, ZN => n17926);
   U17295 : OAI221_X1 port map( B1 => n14370, B2 => n20906, C1 => n14838, C2 =>
                           n20900, A => n17899, ZN => n17898);
   U17296 : AOI22_X1 port map( A1 => n20894, A2 => n19128, B1 => n20888, B2 => 
                           n19129, ZN => n17899);
   U17297 : OAI221_X1 port map( B1 => n15770, B2 => n20786, C1 => n14772, C2 =>
                           n20780, A => n17908, ZN => n17905);
   U17298 : AOI22_X1 port map( A1 => n20774, A2 => n8887, B1 => n20768, B2 => 
                           n19139, ZN => n17908);
   U17299 : OAI221_X1 port map( B1 => n14369, B2 => n20906, C1 => n14837, C2 =>
                           n20900, A => n17881, ZN => n17880);
   U17300 : AOI22_X1 port map( A1 => n20894, A2 => n19108, B1 => n20888, B2 => 
                           n19109, ZN => n17881);
   U17301 : OAI221_X1 port map( B1 => n15769, B2 => n20786, C1 => n14771, C2 =>
                           n20780, A => n17890, ZN => n17887);
   U17302 : AOI22_X1 port map( A1 => n20774, A2 => n8885, B1 => n20768, B2 => 
                           n19119, ZN => n17890);
   U17303 : OAI221_X1 port map( B1 => n14368, B2 => n20907, C1 => n14836, C2 =>
                           n20901, A => n17863, ZN => n17862);
   U17304 : AOI22_X1 port map( A1 => n20895, A2 => n19088, B1 => n20889, B2 => 
                           n19089, ZN => n17863);
   U17305 : OAI221_X1 port map( B1 => n15768, B2 => n20787, C1 => n14770, C2 =>
                           n20781, A => n17872, ZN => n17869);
   U17306 : AOI22_X1 port map( A1 => n20775, A2 => n8883, B1 => n20769, B2 => 
                           n19099, ZN => n17872);
   U17307 : OAI221_X1 port map( B1 => n14367, B2 => n20907, C1 => n14835, C2 =>
                           n20901, A => n17845, ZN => n17844);
   U17308 : AOI22_X1 port map( A1 => n20895, A2 => n19068, B1 => n20889, B2 => 
                           n19069, ZN => n17845);
   U17309 : OAI221_X1 port map( B1 => n15767, B2 => n20787, C1 => n14769, C2 =>
                           n20781, A => n17854, ZN => n17851);
   U17310 : AOI22_X1 port map( A1 => n20775, A2 => n8881, B1 => n20769, B2 => 
                           n19079, ZN => n17854);
   U17311 : OAI221_X1 port map( B1 => n14366, B2 => n20907, C1 => n14834, C2 =>
                           n20901, A => n17827, ZN => n17826);
   U17312 : AOI22_X1 port map( A1 => n20895, A2 => n19048, B1 => n20889, B2 => 
                           n19049, ZN => n17827);
   U17313 : OAI221_X1 port map( B1 => n15766, B2 => n20787, C1 => n14768, C2 =>
                           n20781, A => n17836, ZN => n17833);
   U17314 : AOI22_X1 port map( A1 => n20775, A2 => n8879, B1 => n20769, B2 => 
                           n19059, ZN => n17836);
   U17315 : OAI221_X1 port map( B1 => n14365, B2 => n20907, C1 => n14833, C2 =>
                           n20901, A => n17809, ZN => n17808);
   U17316 : AOI22_X1 port map( A1 => n20895, A2 => n19028, B1 => n20889, B2 => 
                           n19029, ZN => n17809);
   U17317 : OAI221_X1 port map( B1 => n15765, B2 => n20787, C1 => n14767, C2 =>
                           n20781, A => n17818, ZN => n17815);
   U17318 : AOI22_X1 port map( A1 => n20775, A2 => n8877, B1 => n20769, B2 => 
                           n19039, ZN => n17818);
   U17319 : OAI221_X1 port map( B1 => n14364, B2 => n20907, C1 => n14832, C2 =>
                           n20901, A => n17791, ZN => n17790);
   U17320 : AOI22_X1 port map( A1 => n20895, A2 => n19008, B1 => n20889, B2 => 
                           n19009, ZN => n17791);
   U17321 : OAI221_X1 port map( B1 => n15764, B2 => n20787, C1 => n14766, C2 =>
                           n20781, A => n17800, ZN => n17797);
   U17322 : AOI22_X1 port map( A1 => n20775, A2 => n8875, B1 => n20769, B2 => 
                           n19019, ZN => n17800);
   U17323 : OAI221_X1 port map( B1 => n14363, B2 => n20907, C1 => n14831, C2 =>
                           n20901, A => n17773, ZN => n17772);
   U17324 : AOI22_X1 port map( A1 => n20895, A2 => n18988, B1 => n20889, B2 => 
                           n18989, ZN => n17773);
   U17325 : OAI221_X1 port map( B1 => n15763, B2 => n20787, C1 => n14765, C2 =>
                           n20781, A => n17782, ZN => n17779);
   U17326 : AOI22_X1 port map( A1 => n20775, A2 => n8873, B1 => n20769, B2 => 
                           n18999, ZN => n17782);
   U17327 : OAI221_X1 port map( B1 => n14362, B2 => n20907, C1 => n14830, C2 =>
                           n20901, A => n17755, ZN => n17754);
   U17328 : AOI22_X1 port map( A1 => n20895, A2 => n18968, B1 => n20889, B2 => 
                           n18969, ZN => n17755);
   U17329 : OAI221_X1 port map( B1 => n15762, B2 => n20787, C1 => n14764, C2 =>
                           n20781, A => n17764, ZN => n17761);
   U17330 : AOI22_X1 port map( A1 => n20775, A2 => n8871, B1 => n20769, B2 => 
                           n18979, ZN => n17764);
   U17331 : OAI221_X1 port map( B1 => n14361, B2 => n20907, C1 => n14829, C2 =>
                           n20901, A => n17737, ZN => n17736);
   U17332 : AOI22_X1 port map( A1 => n20895, A2 => n18948, B1 => n20889, B2 => 
                           n18949, ZN => n17737);
   U17333 : OAI221_X1 port map( B1 => n15761, B2 => n20787, C1 => n14763, C2 =>
                           n20781, A => n17746, ZN => n17743);
   U17334 : AOI22_X1 port map( A1 => n20775, A2 => n8869, B1 => n20769, B2 => 
                           n18959, ZN => n17746);
   U17335 : OAI221_X1 port map( B1 => n14360, B2 => n20907, C1 => n14828, C2 =>
                           n20901, A => n17719, ZN => n17718);
   U17336 : AOI22_X1 port map( A1 => n20895, A2 => n18928, B1 => n20889, B2 => 
                           n18929, ZN => n17719);
   U17337 : OAI221_X1 port map( B1 => n15760, B2 => n20787, C1 => n14762, C2 =>
                           n20781, A => n17728, ZN => n17725);
   U17338 : AOI22_X1 port map( A1 => n20775, A2 => n8867, B1 => n20769, B2 => 
                           n18939, ZN => n17728);
   U17339 : OAI221_X1 port map( B1 => n14359, B2 => n20907, C1 => n14827, C2 =>
                           n20901, A => n17701, ZN => n17700);
   U17340 : AOI22_X1 port map( A1 => n20895, A2 => n18908, B1 => n20889, B2 => 
                           n18909, ZN => n17701);
   U17341 : OAI221_X1 port map( B1 => n15759, B2 => n20787, C1 => n14761, C2 =>
                           n20781, A => n17710, ZN => n17707);
   U17342 : AOI22_X1 port map( A1 => n20775, A2 => n8865, B1 => n20769, B2 => 
                           n18919, ZN => n17710);
   U17343 : OAI221_X1 port map( B1 => n14358, B2 => n20907, C1 => n14826, C2 =>
                           n20901, A => n17683, ZN => n17682);
   U17344 : AOI22_X1 port map( A1 => n20895, A2 => n18888, B1 => n20889, B2 => 
                           n18889, ZN => n17683);
   U17345 : OAI221_X1 port map( B1 => n15758, B2 => n20787, C1 => n14760, C2 =>
                           n20781, A => n17692, ZN => n17689);
   U17346 : AOI22_X1 port map( A1 => n20775, A2 => n8863, B1 => n20769, B2 => 
                           n18899, ZN => n17692);
   U17347 : OAI221_X1 port map( B1 => n14357, B2 => n20907, C1 => n14825, C2 =>
                           n20901, A => n17665, ZN => n17664);
   U17348 : AOI22_X1 port map( A1 => n20895, A2 => n18868, B1 => n20889, B2 => 
                           n18869, ZN => n17665);
   U17349 : OAI221_X1 port map( B1 => n15757, B2 => n20787, C1 => n14759, C2 =>
                           n20781, A => n17674, ZN => n17671);
   U17350 : AOI22_X1 port map( A1 => n20775, A2 => n8861, B1 => n20769, B2 => 
                           n18879, ZN => n17674);
   U17351 : OAI221_X1 port map( B1 => n14356, B2 => n20908, C1 => n14824, C2 =>
                           n20902, A => n17647, ZN => n17646);
   U17352 : AOI22_X1 port map( A1 => n20896, A2 => n18848, B1 => n20890, B2 => 
                           n18849, ZN => n17647);
   U17353 : OAI221_X1 port map( B1 => n15756, B2 => n20788, C1 => n14758, C2 =>
                           n20782, A => n17656, ZN => n17653);
   U17354 : AOI22_X1 port map( A1 => n20776, A2 => n8859, B1 => n20770, B2 => 
                           n18859, ZN => n17656);
   U17355 : OAI221_X1 port map( B1 => n14355, B2 => n20908, C1 => n14823, C2 =>
                           n20902, A => n17629, ZN => n17628);
   U17356 : AOI22_X1 port map( A1 => n20896, A2 => n18828, B1 => n20890, B2 => 
                           n18829, ZN => n17629);
   U17357 : OAI221_X1 port map( B1 => n15755, B2 => n20788, C1 => n14757, C2 =>
                           n20782, A => n17638, ZN => n17635);
   U17358 : AOI22_X1 port map( A1 => n20776, A2 => n8857, B1 => n20770, B2 => 
                           n18839, ZN => n17638);
   U17359 : OAI221_X1 port map( B1 => n14354, B2 => n20908, C1 => n14822, C2 =>
                           n20902, A => n17611, ZN => n17610);
   U17360 : AOI22_X1 port map( A1 => n20896, A2 => n18808, B1 => n20890, B2 => 
                           n18809, ZN => n17611);
   U17361 : OAI221_X1 port map( B1 => n15754, B2 => n20788, C1 => n14756, C2 =>
                           n20782, A => n17620, ZN => n17617);
   U17362 : AOI22_X1 port map( A1 => n20776, A2 => n8855, B1 => n20770, B2 => 
                           n18819, ZN => n17620);
   U17363 : OAI221_X1 port map( B1 => n14353, B2 => n20908, C1 => n14821, C2 =>
                           n20902, A => n17593, ZN => n17592);
   U17364 : AOI22_X1 port map( A1 => n20896, A2 => n18788, B1 => n20890, B2 => 
                           n18789, ZN => n17593);
   U17365 : OAI221_X1 port map( B1 => n15753, B2 => n20788, C1 => n14755, C2 =>
                           n20782, A => n17602, ZN => n17599);
   U17366 : AOI22_X1 port map( A1 => n20776, A2 => n8853, B1 => n20770, B2 => 
                           n18799, ZN => n17602);
   U17367 : OAI221_X1 port map( B1 => n14352, B2 => n20908, C1 => n14820, C2 =>
                           n20902, A => n17575, ZN => n17574);
   U17368 : AOI22_X1 port map( A1 => n20896, A2 => n18768, B1 => n20890, B2 => 
                           n18769, ZN => n17575);
   U17369 : OAI221_X1 port map( B1 => n15752, B2 => n20788, C1 => n14754, C2 =>
                           n20782, A => n17584, ZN => n17581);
   U17370 : AOI22_X1 port map( A1 => n20776, A2 => n8851, B1 => n20770, B2 => 
                           n18779, ZN => n17584);
   U17371 : OAI221_X1 port map( B1 => n14351, B2 => n20908, C1 => n14819, C2 =>
                           n20902, A => n17557, ZN => n17556);
   U17372 : AOI22_X1 port map( A1 => n20896, A2 => n18748, B1 => n20890, B2 => 
                           n18749, ZN => n17557);
   U17373 : OAI221_X1 port map( B1 => n15751, B2 => n20788, C1 => n14753, C2 =>
                           n20782, A => n17566, ZN => n17563);
   U17374 : AOI22_X1 port map( A1 => n20776, A2 => n8849, B1 => n20770, B2 => 
                           n18759, ZN => n17566);
   U17375 : OAI221_X1 port map( B1 => n14350, B2 => n20908, C1 => n14818, C2 =>
                           n20902, A => n17539, ZN => n17538);
   U17376 : AOI22_X1 port map( A1 => n20896, A2 => n18728, B1 => n20890, B2 => 
                           n18729, ZN => n17539);
   U17377 : OAI221_X1 port map( B1 => n15750, B2 => n20788, C1 => n14752, C2 =>
                           n20782, A => n17548, ZN => n17545);
   U17378 : AOI22_X1 port map( A1 => n20776, A2 => n8847, B1 => n20770, B2 => 
                           n18739, ZN => n17548);
   U17379 : OAI221_X1 port map( B1 => n14349, B2 => n20908, C1 => n14817, C2 =>
                           n20902, A => n17521, ZN => n17520);
   U17380 : AOI22_X1 port map( A1 => n20896, A2 => n18708, B1 => n20890, B2 => 
                           n18709, ZN => n17521);
   U17381 : OAI221_X1 port map( B1 => n15749, B2 => n20788, C1 => n14751, C2 =>
                           n20782, A => n17530, ZN => n17527);
   U17382 : AOI22_X1 port map( A1 => n20776, A2 => n8845, B1 => n20770, B2 => 
                           n18719, ZN => n17530);
   U17383 : OAI221_X1 port map( B1 => n14348, B2 => n20908, C1 => n14816, C2 =>
                           n20902, A => n17503, ZN => n17502);
   U17384 : AOI22_X1 port map( A1 => n20896, A2 => n18688, B1 => n20890, B2 => 
                           n18689, ZN => n17503);
   U17385 : OAI221_X1 port map( B1 => n15748, B2 => n20788, C1 => n14750, C2 =>
                           n20782, A => n17512, ZN => n17509);
   U17386 : AOI22_X1 port map( A1 => n20776, A2 => n8843, B1 => n20770, B2 => 
                           n18699, ZN => n17512);
   U17387 : OAI221_X1 port map( B1 => n14347, B2 => n20908, C1 => n14815, C2 =>
                           n20902, A => n17485, ZN => n17484);
   U17388 : AOI22_X1 port map( A1 => n20896, A2 => n18668, B1 => n20890, B2 => 
                           n18669, ZN => n17485);
   U17389 : OAI221_X1 port map( B1 => n15747, B2 => n20788, C1 => n14749, C2 =>
                           n20782, A => n17494, ZN => n17491);
   U17390 : AOI22_X1 port map( A1 => n20776, A2 => n8841, B1 => n20770, B2 => 
                           n18679, ZN => n17494);
   U17391 : OAI221_X1 port map( B1 => n14346, B2 => n20908, C1 => n14814, C2 =>
                           n20902, A => n17467, ZN => n17466);
   U17392 : AOI22_X1 port map( A1 => n20896, A2 => n18648, B1 => n20890, B2 => 
                           n18649, ZN => n17467);
   U17393 : OAI221_X1 port map( B1 => n15746, B2 => n20788, C1 => n14748, C2 =>
                           n20782, A => n17476, ZN => n17473);
   U17394 : AOI22_X1 port map( A1 => n20776, A2 => n8839, B1 => n20770, B2 => 
                           n18659, ZN => n17476);
   U17395 : OAI221_X1 port map( B1 => n14345, B2 => n20908, C1 => n14813, C2 =>
                           n20902, A => n17449, ZN => n17448);
   U17396 : AOI22_X1 port map( A1 => n20896, A2 => n18628, B1 => n20890, B2 => 
                           n18629, ZN => n17449);
   U17397 : OAI221_X1 port map( B1 => n15745, B2 => n20788, C1 => n14747, C2 =>
                           n20782, A => n17458, ZN => n17455);
   U17398 : AOI22_X1 port map( A1 => n20776, A2 => n8837, B1 => n20770, B2 => 
                           n18639, ZN => n17458);
   U17399 : OAI221_X1 port map( B1 => n14404, B2 => n21110, C1 => n14872, C2 =>
                           n21104, A => n17310, ZN => n17309);
   U17400 : AOI22_X1 port map( A1 => n21098, A2 => n19808, B1 => n21092, B2 => 
                           n19809, ZN => n17310);
   U17401 : OAI221_X1 port map( B1 => n15469, B2 => n21061, C1 => n16068, C2 =>
                           n21055, A => n17321, ZN => n17307);
   U17402 : AOI22_X1 port map( A1 => n21049, A2 => n9211, B1 => n21043, B2 => 
                           n8827, ZN => n17321);
   U17403 : OAI221_X1 port map( B1 => n14271, B2 => n20952, C1 => n15337, C2 =>
                           n20946, A => n17335, ZN => n17326);
   U17404 : AOI22_X1 port map( A1 => n20940, A2 => n19814, B1 => n20934, B2 => 
                           n19815, ZN => n17335);
   U17405 : OAI221_X1 port map( B1 => n15804, B2 => n20976, C1 => n14806, C2 =>
                           n20970, A => n17332, ZN => n17327);
   U17406 : AOI22_X1 port map( A1 => n20964, A2 => n8955, B1 => n20958, B2 => 
                           n19819, ZN => n17332);
   U17407 : OAI221_X1 port map( B1 => n14403, B2 => n21110, C1 => n14871, C2 =>
                           n21104, A => n17290, ZN => n17289);
   U17408 : AOI22_X1 port map( A1 => n21098, A2 => n19788, B1 => n21092, B2 => 
                           n19789, ZN => n17290);
   U17409 : OAI221_X1 port map( B1 => n15468, B2 => n21061, C1 => n16067, C2 =>
                           n21055, A => n17292, ZN => n17287);
   U17410 : AOI22_X1 port map( A1 => n21049, A2 => n9207, B1 => n21043, B2 => 
                           n8823, ZN => n17292);
   U17411 : OAI221_X1 port map( B1 => n14270, B2 => n20952, C1 => n15336, C2 =>
                           n20946, A => n17300, ZN => n17295);
   U17412 : AOI22_X1 port map( A1 => n20940, A2 => n19794, B1 => n20934, B2 => 
                           n19795, ZN => n17300);
   U17413 : OAI221_X1 port map( B1 => n15803, B2 => n20976, C1 => n14805, C2 =>
                           n20970, A => n17299, ZN => n17296);
   U17414 : AOI22_X1 port map( A1 => n20964, A2 => n8953, B1 => n20958, B2 => 
                           n19799, ZN => n17299);
   U17415 : OAI221_X1 port map( B1 => n14402, B2 => n21110, C1 => n14870, C2 =>
                           n21104, A => n17271, ZN => n17270);
   U17416 : AOI22_X1 port map( A1 => n21098, A2 => n19768, B1 => n21092, B2 => 
                           n19769, ZN => n17271);
   U17417 : OAI221_X1 port map( B1 => n15467, B2 => n21061, C1 => n16066, C2 =>
                           n21055, A => n17273, ZN => n17268);
   U17418 : AOI22_X1 port map( A1 => n21049, A2 => n9203, B1 => n21043, B2 => 
                           n8819, ZN => n17273);
   U17419 : OAI221_X1 port map( B1 => n14269, B2 => n20952, C1 => n15335, C2 =>
                           n20946, A => n17281, ZN => n17276);
   U17420 : AOI22_X1 port map( A1 => n20940, A2 => n19774, B1 => n20934, B2 => 
                           n19775, ZN => n17281);
   U17421 : OAI221_X1 port map( B1 => n15802, B2 => n20976, C1 => n14804, C2 =>
                           n20970, A => n17280, ZN => n17277);
   U17422 : AOI22_X1 port map( A1 => n20964, A2 => n8951, B1 => n20958, B2 => 
                           n19779, ZN => n17280);
   U17423 : OAI221_X1 port map( B1 => n14401, B2 => n21110, C1 => n14869, C2 =>
                           n21104, A => n17252, ZN => n17251);
   U17424 : AOI22_X1 port map( A1 => n21098, A2 => n19748, B1 => n21092, B2 => 
                           n19749, ZN => n17252);
   U17425 : OAI221_X1 port map( B1 => n15466, B2 => n21061, C1 => n16065, C2 =>
                           n21055, A => n17254, ZN => n17249);
   U17426 : AOI22_X1 port map( A1 => n21049, A2 => n9199, B1 => n21043, B2 => 
                           n8815, ZN => n17254);
   U17427 : OAI221_X1 port map( B1 => n14268, B2 => n20952, C1 => n15334, C2 =>
                           n20946, A => n17262, ZN => n17257);
   U17428 : AOI22_X1 port map( A1 => n20940, A2 => n19754, B1 => n20934, B2 => 
                           n19755, ZN => n17262);
   U17429 : OAI221_X1 port map( B1 => n15801, B2 => n20976, C1 => n14803, C2 =>
                           n20970, A => n17261, ZN => n17258);
   U17430 : AOI22_X1 port map( A1 => n20964, A2 => n8949, B1 => n20958, B2 => 
                           n19759, ZN => n17261);
   U17431 : OAI221_X1 port map( B1 => n14602, B2 => n21077, C1 => n14934, C2 =>
                           n21067, A => n17234, ZN => n17231);
   U17432 : AOI22_X1 port map( A1 => n19724, A2 => n21086, B1 => n21085, B2 => 
                           n19725, ZN => n17234);
   U17433 : OAI221_X1 port map( B1 => n14400, B2 => n21110, C1 => n14868, C2 =>
                           n21104, A => n17233, ZN => n17232);
   U17434 : AOI22_X1 port map( A1 => n21098, A2 => n19728, B1 => n21092, B2 => 
                           n19729, ZN => n17233);
   U17435 : OAI221_X1 port map( B1 => n15465, B2 => n21061, C1 => n16064, C2 =>
                           n21055, A => n17235, ZN => n17230);
   U17436 : AOI22_X1 port map( A1 => n21049, A2 => n9195, B1 => n21043, B2 => 
                           n8811, ZN => n17235);
   U17437 : OAI221_X1 port map( B1 => n14267, B2 => n20952, C1 => n15333, C2 =>
                           n20946, A => n17243, ZN => n17238);
   U17438 : AOI22_X1 port map( A1 => n20940, A2 => n19734, B1 => n20934, B2 => 
                           n19735, ZN => n17243);
   U17439 : OAI221_X1 port map( B1 => n15800, B2 => n20976, C1 => n14802, C2 =>
                           n20970, A => n17242, ZN => n17239);
   U17440 : AOI22_X1 port map( A1 => n20964, A2 => n8947, B1 => n20958, B2 => 
                           n19739, ZN => n17242);
   U17441 : OAI221_X1 port map( B1 => n14601, B2 => n21077, C1 => n14933, C2 =>
                           n21067, A => n17215, ZN => n17212);
   U17442 : AOI22_X1 port map( A1 => n19704, A2 => n21086, B1 => n21085, B2 => 
                           n19705, ZN => n17215);
   U17443 : OAI221_X1 port map( B1 => n14399, B2 => n21110, C1 => n14867, C2 =>
                           n21104, A => n17214, ZN => n17213);
   U17444 : AOI22_X1 port map( A1 => n21098, A2 => n19708, B1 => n21092, B2 => 
                           n19709, ZN => n17214);
   U17445 : OAI221_X1 port map( B1 => n15464, B2 => n21061, C1 => n16063, C2 =>
                           n21055, A => n17216, ZN => n17211);
   U17446 : AOI22_X1 port map( A1 => n21049, A2 => n9191, B1 => n21043, B2 => 
                           n8807, ZN => n17216);
   U17447 : OAI221_X1 port map( B1 => n14266, B2 => n20952, C1 => n15332, C2 =>
                           n20946, A => n17224, ZN => n17219);
   U17448 : AOI22_X1 port map( A1 => n20940, A2 => n19714, B1 => n20934, B2 => 
                           n19715, ZN => n17224);
   U17449 : OAI221_X1 port map( B1 => n15799, B2 => n20976, C1 => n14801, C2 =>
                           n20970, A => n17223, ZN => n17220);
   U17450 : AOI22_X1 port map( A1 => n20964, A2 => n8945, B1 => n20958, B2 => 
                           n19719, ZN => n17223);
   U17451 : OAI221_X1 port map( B1 => n14600, B2 => n21077, C1 => n14932, C2 =>
                           n21067, A => n17196, ZN => n17193);
   U17452 : AOI22_X1 port map( A1 => n19684, A2 => n21086, B1 => n21085, B2 => 
                           n19685, ZN => n17196);
   U17453 : OAI221_X1 port map( B1 => n14398, B2 => n21110, C1 => n14866, C2 =>
                           n21104, A => n17195, ZN => n17194);
   U17454 : AOI22_X1 port map( A1 => n21098, A2 => n19688, B1 => n21092, B2 => 
                           n19689, ZN => n17195);
   U17455 : OAI221_X1 port map( B1 => n15463, B2 => n21061, C1 => n16062, C2 =>
                           n21055, A => n17197, ZN => n17192);
   U17456 : AOI22_X1 port map( A1 => n21049, A2 => n9187, B1 => n21043, B2 => 
                           n8803, ZN => n17197);
   U17457 : OAI221_X1 port map( B1 => n14265, B2 => n20952, C1 => n15331, C2 =>
                           n20946, A => n17205, ZN => n17200);
   U17458 : AOI22_X1 port map( A1 => n20940, A2 => n19694, B1 => n20934, B2 => 
                           n19695, ZN => n17205);
   U17459 : OAI221_X1 port map( B1 => n15798, B2 => n20976, C1 => n14800, C2 =>
                           n20970, A => n17204, ZN => n17201);
   U17460 : AOI22_X1 port map( A1 => n20964, A2 => n8943, B1 => n20958, B2 => 
                           n19699, ZN => n17204);
   U17461 : OAI221_X1 port map( B1 => n14599, B2 => n21077, C1 => n14931, C2 =>
                           n21067, A => n17177, ZN => n17174);
   U17462 : AOI22_X1 port map( A1 => n19664, A2 => n21086, B1 => n21085, B2 => 
                           n19665, ZN => n17177);
   U17463 : OAI221_X1 port map( B1 => n14397, B2 => n21110, C1 => n14865, C2 =>
                           n21104, A => n17176, ZN => n17175);
   U17464 : AOI22_X1 port map( A1 => n21098, A2 => n19668, B1 => n21092, B2 => 
                           n19669, ZN => n17176);
   U17465 : OAI221_X1 port map( B1 => n15462, B2 => n21061, C1 => n16061, C2 =>
                           n21055, A => n17178, ZN => n17173);
   U17466 : AOI22_X1 port map( A1 => n21049, A2 => n9183, B1 => n21043, B2 => 
                           n8799, ZN => n17178);
   U17467 : OAI221_X1 port map( B1 => n14264, B2 => n20952, C1 => n15330, C2 =>
                           n20946, A => n17186, ZN => n17181);
   U17468 : AOI22_X1 port map( A1 => n20940, A2 => n19674, B1 => n20934, B2 => 
                           n19675, ZN => n17186);
   U17469 : OAI221_X1 port map( B1 => n15797, B2 => n20976, C1 => n14799, C2 =>
                           n20970, A => n17185, ZN => n17182);
   U17470 : AOI22_X1 port map( A1 => n20964, A2 => n8941, B1 => n20958, B2 => 
                           n19679, ZN => n17185);
   U17471 : OAI221_X1 port map( B1 => n14598, B2 => n21077, C1 => n14930, C2 =>
                           n21067, A => n17158, ZN => n17155);
   U17472 : AOI22_X1 port map( A1 => n19644, A2 => n21086, B1 => n21085, B2 => 
                           n19645, ZN => n17158);
   U17473 : OAI221_X1 port map( B1 => n14396, B2 => n21110, C1 => n14864, C2 =>
                           n21104, A => n17157, ZN => n17156);
   U17474 : AOI22_X1 port map( A1 => n21098, A2 => n19648, B1 => n21092, B2 => 
                           n19649, ZN => n17157);
   U17475 : OAI221_X1 port map( B1 => n15461, B2 => n21061, C1 => n16060, C2 =>
                           n21055, A => n17159, ZN => n17154);
   U17476 : AOI22_X1 port map( A1 => n21049, A2 => n9179, B1 => n21043, B2 => 
                           n8795, ZN => n17159);
   U17477 : OAI221_X1 port map( B1 => n14263, B2 => n20952, C1 => n15329, C2 =>
                           n20946, A => n17167, ZN => n17162);
   U17478 : AOI22_X1 port map( A1 => n20940, A2 => n19654, B1 => n20934, B2 => 
                           n19655, ZN => n17167);
   U17479 : OAI221_X1 port map( B1 => n15796, B2 => n20976, C1 => n14798, C2 =>
                           n20970, A => n17166, ZN => n17163);
   U17480 : AOI22_X1 port map( A1 => n20964, A2 => n8939, B1 => n20958, B2 => 
                           n19659, ZN => n17166);
   U17481 : OAI221_X1 port map( B1 => n14395, B2 => n21110, C1 => n14863, C2 =>
                           n21104, A => n17138, ZN => n17137);
   U17482 : AOI22_X1 port map( A1 => n21098, A2 => n19628, B1 => n21092, B2 => 
                           n19629, ZN => n17138);
   U17483 : OAI221_X1 port map( B1 => n15460, B2 => n21061, C1 => n16059, C2 =>
                           n21055, A => n17140, ZN => n17135);
   U17484 : AOI22_X1 port map( A1 => n21049, A2 => n9175, B1 => n21043, B2 => 
                           n8791, ZN => n17140);
   U17485 : OAI221_X1 port map( B1 => n14262, B2 => n20952, C1 => n15328, C2 =>
                           n20946, A => n17148, ZN => n17143);
   U17486 : AOI22_X1 port map( A1 => n20940, A2 => n19634, B1 => n20934, B2 => 
                           n19635, ZN => n17148);
   U17487 : OAI221_X1 port map( B1 => n15795, B2 => n20976, C1 => n14797, C2 =>
                           n20970, A => n17147, ZN => n17144);
   U17488 : AOI22_X1 port map( A1 => n20964, A2 => n8937, B1 => n20958, B2 => 
                           n19639, ZN => n17147);
   U17489 : OAI221_X1 port map( B1 => n14394, B2 => n21110, C1 => n14862, C2 =>
                           n21104, A => n17119, ZN => n17118);
   U17490 : AOI22_X1 port map( A1 => n21098, A2 => n19608, B1 => n21092, B2 => 
                           n19609, ZN => n17119);
   U17491 : OAI221_X1 port map( B1 => n15459, B2 => n21061, C1 => n16058, C2 =>
                           n21055, A => n17121, ZN => n17116);
   U17492 : AOI22_X1 port map( A1 => n21049, A2 => n9171, B1 => n21043, B2 => 
                           n8787, ZN => n17121);
   U17493 : OAI221_X1 port map( B1 => n14261, B2 => n20952, C1 => n15327, C2 =>
                           n20946, A => n17129, ZN => n17124);
   U17494 : AOI22_X1 port map( A1 => n20940, A2 => n19614, B1 => n20934, B2 => 
                           n19615, ZN => n17129);
   U17495 : OAI221_X1 port map( B1 => n15794, B2 => n20976, C1 => n14796, C2 =>
                           n20970, A => n17128, ZN => n17125);
   U17496 : AOI22_X1 port map( A1 => n20964, A2 => n8935, B1 => n20958, B2 => 
                           n19619, ZN => n17128);
   U17497 : OAI221_X1 port map( B1 => n14393, B2 => n21110, C1 => n14861, C2 =>
                           n21104, A => n17100, ZN => n17099);
   U17498 : AOI22_X1 port map( A1 => n21098, A2 => n19588, B1 => n21092, B2 => 
                           n19589, ZN => n17100);
   U17499 : OAI221_X1 port map( B1 => n15458, B2 => n21061, C1 => n16057, C2 =>
                           n21055, A => n17102, ZN => n17097);
   U17500 : AOI22_X1 port map( A1 => n21049, A2 => n9167, B1 => n21043, B2 => 
                           n8783, ZN => n17102);
   U17501 : OAI221_X1 port map( B1 => n14260, B2 => n20952, C1 => n15326, C2 =>
                           n20946, A => n17110, ZN => n17105);
   U17502 : AOI22_X1 port map( A1 => n20940, A2 => n19594, B1 => n20934, B2 => 
                           n19595, ZN => n17110);
   U17503 : OAI221_X1 port map( B1 => n15793, B2 => n20976, C1 => n14795, C2 =>
                           n20970, A => n17109, ZN => n17106);
   U17504 : AOI22_X1 port map( A1 => n20964, A2 => n8933, B1 => n20958, B2 => 
                           n19599, ZN => n17109);
   U17505 : OAI221_X1 port map( B1 => n14392, B2 => n21111, C1 => n14860, C2 =>
                           n21105, A => n17081, ZN => n17080);
   U17506 : AOI22_X1 port map( A1 => n21099, A2 => n19568, B1 => n21093, B2 => 
                           n19569, ZN => n17081);
   U17507 : OAI221_X1 port map( B1 => n15457, B2 => n21062, C1 => n16056, C2 =>
                           n21056, A => n17083, ZN => n17078);
   U17508 : AOI22_X1 port map( A1 => n21050, A2 => n9163, B1 => n21044, B2 => 
                           n8779, ZN => n17083);
   U17509 : OAI221_X1 port map( B1 => n15792, B2 => n20977, C1 => n14794, C2 =>
                           n20971, A => n17090, ZN => n17087);
   U17510 : AOI22_X1 port map( A1 => n20965, A2 => n8931, B1 => n20959, B2 => 
                           n19579, ZN => n17090);
   U17511 : OAI221_X1 port map( B1 => n14391, B2 => n21111, C1 => n14859, C2 =>
                           n21105, A => n17062, ZN => n17061);
   U17512 : AOI22_X1 port map( A1 => n21099, A2 => n19548, B1 => n21093, B2 => 
                           n19549, ZN => n17062);
   U17513 : OAI221_X1 port map( B1 => n15456, B2 => n21062, C1 => n16055, C2 =>
                           n21056, A => n17064, ZN => n17059);
   U17514 : AOI22_X1 port map( A1 => n21050, A2 => n9159, B1 => n21044, B2 => 
                           n8775, ZN => n17064);
   U17515 : OAI221_X1 port map( B1 => n15791, B2 => n20977, C1 => n14793, C2 =>
                           n20971, A => n17071, ZN => n17068);
   U17516 : AOI22_X1 port map( A1 => n20965, A2 => n8929, B1 => n20959, B2 => 
                           n19559, ZN => n17071);
   U17517 : OAI221_X1 port map( B1 => n14390, B2 => n21111, C1 => n14858, C2 =>
                           n21105, A => n17043, ZN => n17042);
   U17518 : AOI22_X1 port map( A1 => n21099, A2 => n19528, B1 => n21093, B2 => 
                           n19529, ZN => n17043);
   U17519 : OAI221_X1 port map( B1 => n15455, B2 => n21062, C1 => n16054, C2 =>
                           n21056, A => n17045, ZN => n17040);
   U17520 : AOI22_X1 port map( A1 => n21050, A2 => n9155, B1 => n21044, B2 => 
                           n8771, ZN => n17045);
   U17521 : OAI221_X1 port map( B1 => n15790, B2 => n20977, C1 => n14792, C2 =>
                           n20971, A => n17052, ZN => n17049);
   U17522 : AOI22_X1 port map( A1 => n20965, A2 => n8927, B1 => n20959, B2 => 
                           n19539, ZN => n17052);
   U17523 : OAI221_X1 port map( B1 => n14389, B2 => n21111, C1 => n14857, C2 =>
                           n21105, A => n17024, ZN => n17023);
   U17524 : AOI22_X1 port map( A1 => n21099, A2 => n19508, B1 => n21093, B2 => 
                           n19509, ZN => n17024);
   U17525 : OAI221_X1 port map( B1 => n15454, B2 => n21062, C1 => n16053, C2 =>
                           n21056, A => n17026, ZN => n17021);
   U17526 : AOI22_X1 port map( A1 => n21050, A2 => n9151, B1 => n21044, B2 => 
                           n8767, ZN => n17026);
   U17527 : OAI221_X1 port map( B1 => n15789, B2 => n20977, C1 => n14791, C2 =>
                           n20971, A => n17033, ZN => n17030);
   U17528 : AOI22_X1 port map( A1 => n20965, A2 => n8925, B1 => n20959, B2 => 
                           n19519, ZN => n17033);
   U17529 : OAI221_X1 port map( B1 => n14388, B2 => n21111, C1 => n14856, C2 =>
                           n21105, A => n17005, ZN => n17004);
   U17530 : AOI22_X1 port map( A1 => n21099, A2 => n19488, B1 => n21093, B2 => 
                           n19489, ZN => n17005);
   U17531 : OAI221_X1 port map( B1 => n15453, B2 => n21062, C1 => n16052, C2 =>
                           n21056, A => n17007, ZN => n17002);
   U17532 : AOI22_X1 port map( A1 => n21050, A2 => n9147, B1 => n21044, B2 => 
                           n8763, ZN => n17007);
   U17533 : OAI221_X1 port map( B1 => n15788, B2 => n20977, C1 => n14790, C2 =>
                           n20971, A => n17014, ZN => n17011);
   U17534 : AOI22_X1 port map( A1 => n20965, A2 => n8923, B1 => n20959, B2 => 
                           n19499, ZN => n17014);
   U17535 : OAI221_X1 port map( B1 => n14387, B2 => n21111, C1 => n14855, C2 =>
                           n21105, A => n16986, ZN => n16985);
   U17536 : AOI22_X1 port map( A1 => n21099, A2 => n19468, B1 => n21093, B2 => 
                           n19469, ZN => n16986);
   U17537 : OAI221_X1 port map( B1 => n15452, B2 => n21062, C1 => n16051, C2 =>
                           n21056, A => n16988, ZN => n16983);
   U17538 : AOI22_X1 port map( A1 => n21050, A2 => n9143, B1 => n21044, B2 => 
                           n8759, ZN => n16988);
   U17539 : OAI221_X1 port map( B1 => n15787, B2 => n20977, C1 => n14789, C2 =>
                           n20971, A => n16995, ZN => n16992);
   U17540 : AOI22_X1 port map( A1 => n20965, A2 => n8921, B1 => n20959, B2 => 
                           n19479, ZN => n16995);
   U17541 : OAI221_X1 port map( B1 => n14386, B2 => n21111, C1 => n14854, C2 =>
                           n21105, A => n16967, ZN => n16966);
   U17542 : AOI22_X1 port map( A1 => n21099, A2 => n19448, B1 => n21093, B2 => 
                           n19449, ZN => n16967);
   U17543 : OAI221_X1 port map( B1 => n15451, B2 => n21062, C1 => n16050, C2 =>
                           n21056, A => n16969, ZN => n16964);
   U17544 : AOI22_X1 port map( A1 => n21050, A2 => n9139, B1 => n21044, B2 => 
                           n8755, ZN => n16969);
   U17545 : OAI221_X1 port map( B1 => n15786, B2 => n20977, C1 => n14788, C2 =>
                           n20971, A => n16976, ZN => n16973);
   U17546 : AOI22_X1 port map( A1 => n20965, A2 => n8919, B1 => n20959, B2 => 
                           n19459, ZN => n16976);
   U17547 : OAI221_X1 port map( B1 => n14385, B2 => n21111, C1 => n14853, C2 =>
                           n21105, A => n16948, ZN => n16947);
   U17548 : AOI22_X1 port map( A1 => n21099, A2 => n19428, B1 => n21093, B2 => 
                           n19429, ZN => n16948);
   U17549 : OAI221_X1 port map( B1 => n15450, B2 => n21062, C1 => n16049, C2 =>
                           n21056, A => n16950, ZN => n16945);
   U17550 : AOI22_X1 port map( A1 => n21050, A2 => n9135, B1 => n21044, B2 => 
                           n8751, ZN => n16950);
   U17551 : OAI221_X1 port map( B1 => n15785, B2 => n20977, C1 => n14787, C2 =>
                           n20971, A => n16957, ZN => n16954);
   U17552 : AOI22_X1 port map( A1 => n20965, A2 => n8917, B1 => n20959, B2 => 
                           n19439, ZN => n16957);
   U17553 : OAI221_X1 port map( B1 => n14384, B2 => n21111, C1 => n14852, C2 =>
                           n21105, A => n16929, ZN => n16928);
   U17554 : AOI22_X1 port map( A1 => n21099, A2 => n19408, B1 => n21093, B2 => 
                           n19409, ZN => n16929);
   U17555 : OAI221_X1 port map( B1 => n15449, B2 => n21062, C1 => n16048, C2 =>
                           n21056, A => n16931, ZN => n16926);
   U17556 : AOI22_X1 port map( A1 => n21050, A2 => n9131, B1 => n21044, B2 => 
                           n8747, ZN => n16931);
   U17557 : OAI221_X1 port map( B1 => n15784, B2 => n20977, C1 => n14786, C2 =>
                           n20971, A => n16938, ZN => n16935);
   U17558 : AOI22_X1 port map( A1 => n20965, A2 => n8915, B1 => n20959, B2 => 
                           n19419, ZN => n16938);
   U17559 : OAI221_X1 port map( B1 => n14383, B2 => n21111, C1 => n14851, C2 =>
                           n21105, A => n16910, ZN => n16909);
   U17560 : AOI22_X1 port map( A1 => n21099, A2 => n19388, B1 => n21093, B2 => 
                           n19389, ZN => n16910);
   U17561 : OAI221_X1 port map( B1 => n15448, B2 => n21062, C1 => n16047, C2 =>
                           n21056, A => n16912, ZN => n16907);
   U17562 : AOI22_X1 port map( A1 => n21050, A2 => n9127, B1 => n21044, B2 => 
                           n8743, ZN => n16912);
   U17563 : OAI221_X1 port map( B1 => n15783, B2 => n20977, C1 => n14785, C2 =>
                           n20971, A => n16919, ZN => n16916);
   U17564 : AOI22_X1 port map( A1 => n20965, A2 => n8913, B1 => n20959, B2 => 
                           n19399, ZN => n16919);
   U17565 : OAI221_X1 port map( B1 => n14382, B2 => n21111, C1 => n14850, C2 =>
                           n21105, A => n16891, ZN => n16890);
   U17566 : AOI22_X1 port map( A1 => n21099, A2 => n19368, B1 => n21093, B2 => 
                           n19369, ZN => n16891);
   U17567 : OAI221_X1 port map( B1 => n15447, B2 => n21062, C1 => n16046, C2 =>
                           n21056, A => n16893, ZN => n16888);
   U17568 : AOI22_X1 port map( A1 => n21050, A2 => n9123, B1 => n21044, B2 => 
                           n8739, ZN => n16893);
   U17569 : OAI221_X1 port map( B1 => n15782, B2 => n20977, C1 => n14784, C2 =>
                           n20971, A => n16900, ZN => n16897);
   U17570 : AOI22_X1 port map( A1 => n20965, A2 => n8911, B1 => n20959, B2 => 
                           n19379, ZN => n16900);
   U17571 : OAI221_X1 port map( B1 => n14381, B2 => n21111, C1 => n14849, C2 =>
                           n21105, A => n16872, ZN => n16871);
   U17572 : AOI22_X1 port map( A1 => n21099, A2 => n19348, B1 => n21093, B2 => 
                           n19349, ZN => n16872);
   U17573 : OAI221_X1 port map( B1 => n15446, B2 => n21062, C1 => n16045, C2 =>
                           n21056, A => n16874, ZN => n16869);
   U17574 : AOI22_X1 port map( A1 => n21050, A2 => n9119, B1 => n21044, B2 => 
                           n8735, ZN => n16874);
   U17575 : OAI221_X1 port map( B1 => n15781, B2 => n20977, C1 => n14783, C2 =>
                           n20971, A => n16881, ZN => n16878);
   U17576 : AOI22_X1 port map( A1 => n20965, A2 => n8909, B1 => n20959, B2 => 
                           n19359, ZN => n16881);
   U17577 : OAI221_X1 port map( B1 => n14380, B2 => n21112, C1 => n14848, C2 =>
                           n21106, A => n16853, ZN => n16852);
   U17578 : AOI22_X1 port map( A1 => n21100, A2 => n19328, B1 => n21094, B2 => 
                           n19329, ZN => n16853);
   U17579 : OAI221_X1 port map( B1 => n15445, B2 => n21063, C1 => n16044, C2 =>
                           n21057, A => n16855, ZN => n16850);
   U17580 : AOI22_X1 port map( A1 => n21051, A2 => n9115, B1 => n21045, B2 => 
                           n8731, ZN => n16855);
   U17581 : OAI221_X1 port map( B1 => n15780, B2 => n20978, C1 => n14782, C2 =>
                           n20972, A => n16862, ZN => n16859);
   U17582 : AOI22_X1 port map( A1 => n20966, A2 => n8907, B1 => n20960, B2 => 
                           n19339, ZN => n16862);
   U17583 : OAI221_X1 port map( B1 => n14379, B2 => n21112, C1 => n14847, C2 =>
                           n21106, A => n16834, ZN => n16833);
   U17584 : AOI22_X1 port map( A1 => n21100, A2 => n19308, B1 => n21094, B2 => 
                           n19309, ZN => n16834);
   U17585 : OAI221_X1 port map( B1 => n15444, B2 => n21063, C1 => n16043, C2 =>
                           n21057, A => n16836, ZN => n16831);
   U17586 : AOI22_X1 port map( A1 => n21051, A2 => n9111, B1 => n21045, B2 => 
                           n8727, ZN => n16836);
   U17587 : OAI221_X1 port map( B1 => n15779, B2 => n20978, C1 => n14781, C2 =>
                           n20972, A => n16843, ZN => n16840);
   U17588 : AOI22_X1 port map( A1 => n20966, A2 => n8905, B1 => n20960, B2 => 
                           n19319, ZN => n16843);
   U17589 : OAI221_X1 port map( B1 => n14378, B2 => n21112, C1 => n14846, C2 =>
                           n21106, A => n16815, ZN => n16814);
   U17590 : AOI22_X1 port map( A1 => n21100, A2 => n19288, B1 => n21094, B2 => 
                           n19289, ZN => n16815);
   U17591 : OAI221_X1 port map( B1 => n15443, B2 => n21063, C1 => n16042, C2 =>
                           n21057, A => n16817, ZN => n16812);
   U17592 : AOI22_X1 port map( A1 => n21051, A2 => n9107, B1 => n21045, B2 => 
                           n8723, ZN => n16817);
   U17593 : OAI221_X1 port map( B1 => n15778, B2 => n20978, C1 => n14780, C2 =>
                           n20972, A => n16824, ZN => n16821);
   U17594 : AOI22_X1 port map( A1 => n20966, A2 => n8903, B1 => n20960, B2 => 
                           n19299, ZN => n16824);
   U17595 : OAI221_X1 port map( B1 => n14377, B2 => n21112, C1 => n14845, C2 =>
                           n21106, A => n16796, ZN => n16795);
   U17596 : AOI22_X1 port map( A1 => n21100, A2 => n19268, B1 => n21094, B2 => 
                           n19269, ZN => n16796);
   U17597 : OAI221_X1 port map( B1 => n15442, B2 => n21063, C1 => n16041, C2 =>
                           n21057, A => n16798, ZN => n16793);
   U17598 : AOI22_X1 port map( A1 => n21051, A2 => n9103, B1 => n21045, B2 => 
                           n8719, ZN => n16798);
   U17599 : OAI221_X1 port map( B1 => n15777, B2 => n20978, C1 => n14779, C2 =>
                           n20972, A => n16805, ZN => n16802);
   U17600 : AOI22_X1 port map( A1 => n20966, A2 => n8901, B1 => n20960, B2 => 
                           n19279, ZN => n16805);
   U17601 : OAI221_X1 port map( B1 => n14376, B2 => n21112, C1 => n14844, C2 =>
                           n21106, A => n16777, ZN => n16776);
   U17602 : AOI22_X1 port map( A1 => n21100, A2 => n19248, B1 => n21094, B2 => 
                           n19249, ZN => n16777);
   U17603 : OAI221_X1 port map( B1 => n15441, B2 => n21063, C1 => n16040, C2 =>
                           n21057, A => n16779, ZN => n16774);
   U17604 : AOI22_X1 port map( A1 => n21051, A2 => n9099, B1 => n21045, B2 => 
                           n8715, ZN => n16779);
   U17605 : OAI221_X1 port map( B1 => n15776, B2 => n20978, C1 => n14778, C2 =>
                           n20972, A => n16786, ZN => n16783);
   U17606 : AOI22_X1 port map( A1 => n20966, A2 => n8899, B1 => n20960, B2 => 
                           n19259, ZN => n16786);
   U17607 : OAI221_X1 port map( B1 => n14375, B2 => n21112, C1 => n14843, C2 =>
                           n21106, A => n16758, ZN => n16757);
   U17608 : AOI22_X1 port map( A1 => n21100, A2 => n19228, B1 => n21094, B2 => 
                           n19229, ZN => n16758);
   U17609 : OAI221_X1 port map( B1 => n15440, B2 => n21063, C1 => n16039, C2 =>
                           n21057, A => n16760, ZN => n16755);
   U17610 : AOI22_X1 port map( A1 => n21051, A2 => n9095, B1 => n21045, B2 => 
                           n8711, ZN => n16760);
   U17611 : OAI221_X1 port map( B1 => n15775, B2 => n20978, C1 => n14777, C2 =>
                           n20972, A => n16767, ZN => n16764);
   U17612 : AOI22_X1 port map( A1 => n20966, A2 => n8897, B1 => n20960, B2 => 
                           n19239, ZN => n16767);
   U17613 : OAI221_X1 port map( B1 => n14374, B2 => n21112, C1 => n14842, C2 =>
                           n21106, A => n16739, ZN => n16738);
   U17614 : AOI22_X1 port map( A1 => n21100, A2 => n19208, B1 => n21094, B2 => 
                           n19209, ZN => n16739);
   U17615 : OAI221_X1 port map( B1 => n15439, B2 => n21063, C1 => n16038, C2 =>
                           n21057, A => n16741, ZN => n16736);
   U17616 : AOI22_X1 port map( A1 => n21051, A2 => n9091, B1 => n21045, B2 => 
                           n8707, ZN => n16741);
   U17617 : OAI221_X1 port map( B1 => n15774, B2 => n20978, C1 => n14776, C2 =>
                           n20972, A => n16748, ZN => n16745);
   U17618 : AOI22_X1 port map( A1 => n20966, A2 => n8895, B1 => n20960, B2 => 
                           n19219, ZN => n16748);
   U17619 : OAI221_X1 port map( B1 => n14373, B2 => n21112, C1 => n14841, C2 =>
                           n21106, A => n16720, ZN => n16719);
   U17620 : AOI22_X1 port map( A1 => n21100, A2 => n19188, B1 => n21094, B2 => 
                           n19189, ZN => n16720);
   U17621 : OAI221_X1 port map( B1 => n15438, B2 => n21063, C1 => n16037, C2 =>
                           n21057, A => n16722, ZN => n16717);
   U17622 : AOI22_X1 port map( A1 => n21051, A2 => n9087, B1 => n21045, B2 => 
                           n8703, ZN => n16722);
   U17623 : OAI221_X1 port map( B1 => n15773, B2 => n20978, C1 => n14775, C2 =>
                           n20972, A => n16729, ZN => n16726);
   U17624 : AOI22_X1 port map( A1 => n20966, A2 => n8893, B1 => n20960, B2 => 
                           n19199, ZN => n16729);
   U17625 : OAI221_X1 port map( B1 => n14372, B2 => n21112, C1 => n14840, C2 =>
                           n21106, A => n16701, ZN => n16700);
   U17626 : AOI22_X1 port map( A1 => n21100, A2 => n19168, B1 => n21094, B2 => 
                           n19169, ZN => n16701);
   U17627 : OAI221_X1 port map( B1 => n15437, B2 => n21063, C1 => n16036, C2 =>
                           n21057, A => n16703, ZN => n16698);
   U17628 : AOI22_X1 port map( A1 => n21051, A2 => n9083, B1 => n21045, B2 => 
                           n8699, ZN => n16703);
   U17629 : OAI221_X1 port map( B1 => n15772, B2 => n20978, C1 => n14774, C2 =>
                           n20972, A => n16710, ZN => n16707);
   U17630 : AOI22_X1 port map( A1 => n20966, A2 => n8891, B1 => n20960, B2 => 
                           n19179, ZN => n16710);
   U17631 : OAI221_X1 port map( B1 => n14371, B2 => n21112, C1 => n14839, C2 =>
                           n21106, A => n16682, ZN => n16681);
   U17632 : AOI22_X1 port map( A1 => n21100, A2 => n19148, B1 => n21094, B2 => 
                           n19149, ZN => n16682);
   U17633 : OAI221_X1 port map( B1 => n15436, B2 => n21063, C1 => n16035, C2 =>
                           n21057, A => n16684, ZN => n16679);
   U17634 : AOI22_X1 port map( A1 => n21051, A2 => n9079, B1 => n21045, B2 => 
                           n8695, ZN => n16684);
   U17635 : OAI221_X1 port map( B1 => n15771, B2 => n20978, C1 => n14773, C2 =>
                           n20972, A => n16691, ZN => n16688);
   U17636 : AOI22_X1 port map( A1 => n20966, A2 => n8889, B1 => n20960, B2 => 
                           n19159, ZN => n16691);
   U17637 : OAI221_X1 port map( B1 => n14370, B2 => n21112, C1 => n14838, C2 =>
                           n21106, A => n16663, ZN => n16662);
   U17638 : AOI22_X1 port map( A1 => n21100, A2 => n19128, B1 => n21094, B2 => 
                           n19129, ZN => n16663);
   U17639 : OAI221_X1 port map( B1 => n15435, B2 => n21063, C1 => n16034, C2 =>
                           n21057, A => n16665, ZN => n16660);
   U17640 : AOI22_X1 port map( A1 => n21051, A2 => n9075, B1 => n21045, B2 => 
                           n8691, ZN => n16665);
   U17641 : OAI221_X1 port map( B1 => n15770, B2 => n20978, C1 => n14772, C2 =>
                           n20972, A => n16672, ZN => n16669);
   U17642 : AOI22_X1 port map( A1 => n20966, A2 => n8887, B1 => n20960, B2 => 
                           n19139, ZN => n16672);
   U17643 : OAI221_X1 port map( B1 => n14369, B2 => n21112, C1 => n14837, C2 =>
                           n21106, A => n16644, ZN => n16643);
   U17644 : AOI22_X1 port map( A1 => n21100, A2 => n19108, B1 => n21094, B2 => 
                           n19109, ZN => n16644);
   U17645 : OAI221_X1 port map( B1 => n15434, B2 => n21063, C1 => n16033, C2 =>
                           n21057, A => n16646, ZN => n16641);
   U17646 : AOI22_X1 port map( A1 => n21051, A2 => n9071, B1 => n21045, B2 => 
                           n8687, ZN => n16646);
   U17647 : OAI221_X1 port map( B1 => n15769, B2 => n20978, C1 => n14771, C2 =>
                           n20972, A => n16653, ZN => n16650);
   U17648 : AOI22_X1 port map( A1 => n20966, A2 => n8885, B1 => n20960, B2 => 
                           n19119, ZN => n16653);
   U17649 : OAI221_X1 port map( B1 => n14368, B2 => n21113, C1 => n14836, C2 =>
                           n21107, A => n16625, ZN => n16624);
   U17650 : AOI22_X1 port map( A1 => n21101, A2 => n19088, B1 => n21095, B2 => 
                           n19089, ZN => n16625);
   U17651 : OAI221_X1 port map( B1 => n15433, B2 => n21064, C1 => n16032, C2 =>
                           n21058, A => n16627, ZN => n16622);
   U17652 : AOI22_X1 port map( A1 => n21052, A2 => n9067, B1 => n21046, B2 => 
                           n8683, ZN => n16627);
   U17653 : OAI221_X1 port map( B1 => n15768, B2 => n20979, C1 => n14770, C2 =>
                           n20973, A => n16634, ZN => n16631);
   U17654 : AOI22_X1 port map( A1 => n20967, A2 => n8883, B1 => n20961, B2 => 
                           n19099, ZN => n16634);
   U17655 : OAI221_X1 port map( B1 => n14367, B2 => n21113, C1 => n14835, C2 =>
                           n21107, A => n16606, ZN => n16605);
   U17656 : AOI22_X1 port map( A1 => n21101, A2 => n19068, B1 => n21095, B2 => 
                           n19069, ZN => n16606);
   U17657 : OAI221_X1 port map( B1 => n15432, B2 => n21064, C1 => n16031, C2 =>
                           n21058, A => n16608, ZN => n16603);
   U17658 : AOI22_X1 port map( A1 => n21052, A2 => n9063, B1 => n21046, B2 => 
                           n8679, ZN => n16608);
   U17659 : OAI221_X1 port map( B1 => n15767, B2 => n20979, C1 => n14769, C2 =>
                           n20973, A => n16615, ZN => n16612);
   U17660 : AOI22_X1 port map( A1 => n20967, A2 => n8881, B1 => n20961, B2 => 
                           n19079, ZN => n16615);
   U17661 : OAI221_X1 port map( B1 => n14366, B2 => n21113, C1 => n14834, C2 =>
                           n21107, A => n16587, ZN => n16586);
   U17662 : AOI22_X1 port map( A1 => n21101, A2 => n19048, B1 => n21095, B2 => 
                           n19049, ZN => n16587);
   U17663 : OAI221_X1 port map( B1 => n15431, B2 => n21064, C1 => n16030, C2 =>
                           n21058, A => n16589, ZN => n16584);
   U17664 : AOI22_X1 port map( A1 => n21052, A2 => n9059, B1 => n21046, B2 => 
                           n8675, ZN => n16589);
   U17665 : OAI221_X1 port map( B1 => n15766, B2 => n20979, C1 => n14768, C2 =>
                           n20973, A => n16596, ZN => n16593);
   U17666 : AOI22_X1 port map( A1 => n20967, A2 => n8879, B1 => n20961, B2 => 
                           n19059, ZN => n16596);
   U17667 : OAI221_X1 port map( B1 => n14365, B2 => n21113, C1 => n14833, C2 =>
                           n21107, A => n16568, ZN => n16567);
   U17668 : AOI22_X1 port map( A1 => n21101, A2 => n19028, B1 => n21095, B2 => 
                           n19029, ZN => n16568);
   U17669 : OAI221_X1 port map( B1 => n15430, B2 => n21064, C1 => n16029, C2 =>
                           n21058, A => n16570, ZN => n16565);
   U17670 : AOI22_X1 port map( A1 => n21052, A2 => n9055, B1 => n21046, B2 => 
                           n8671, ZN => n16570);
   U17671 : OAI221_X1 port map( B1 => n15765, B2 => n20979, C1 => n14767, C2 =>
                           n20973, A => n16577, ZN => n16574);
   U17672 : AOI22_X1 port map( A1 => n20967, A2 => n8877, B1 => n20961, B2 => 
                           n19039, ZN => n16577);
   U17673 : OAI221_X1 port map( B1 => n14364, B2 => n21113, C1 => n14832, C2 =>
                           n21107, A => n16549, ZN => n16548);
   U17674 : AOI22_X1 port map( A1 => n21101, A2 => n19008, B1 => n21095, B2 => 
                           n19009, ZN => n16549);
   U17675 : OAI221_X1 port map( B1 => n15429, B2 => n21064, C1 => n16028, C2 =>
                           n21058, A => n16551, ZN => n16546);
   U17676 : AOI22_X1 port map( A1 => n21052, A2 => n9051, B1 => n21046, B2 => 
                           n8667, ZN => n16551);
   U17677 : OAI221_X1 port map( B1 => n15764, B2 => n20979, C1 => n14766, C2 =>
                           n20973, A => n16558, ZN => n16555);
   U17678 : AOI22_X1 port map( A1 => n20967, A2 => n8875, B1 => n20961, B2 => 
                           n19019, ZN => n16558);
   U17679 : OAI221_X1 port map( B1 => n14363, B2 => n21113, C1 => n14831, C2 =>
                           n21107, A => n16530, ZN => n16529);
   U17680 : AOI22_X1 port map( A1 => n21101, A2 => n18988, B1 => n21095, B2 => 
                           n18989, ZN => n16530);
   U17681 : OAI221_X1 port map( B1 => n15428, B2 => n21064, C1 => n16027, C2 =>
                           n21058, A => n16532, ZN => n16527);
   U17682 : AOI22_X1 port map( A1 => n21052, A2 => n9047, B1 => n21046, B2 => 
                           n8663, ZN => n16532);
   U17683 : OAI221_X1 port map( B1 => n15763, B2 => n20979, C1 => n14765, C2 =>
                           n20973, A => n16539, ZN => n16536);
   U17684 : AOI22_X1 port map( A1 => n20967, A2 => n8873, B1 => n20961, B2 => 
                           n18999, ZN => n16539);
   U17685 : OAI221_X1 port map( B1 => n14362, B2 => n21113, C1 => n14830, C2 =>
                           n21107, A => n16511, ZN => n16510);
   U17686 : AOI22_X1 port map( A1 => n21101, A2 => n18968, B1 => n21095, B2 => 
                           n18969, ZN => n16511);
   U17687 : OAI221_X1 port map( B1 => n15427, B2 => n21064, C1 => n16026, C2 =>
                           n21058, A => n16513, ZN => n16508);
   U17688 : AOI22_X1 port map( A1 => n21052, A2 => n9043, B1 => n21046, B2 => 
                           n8659, ZN => n16513);
   U17689 : OAI221_X1 port map( B1 => n15762, B2 => n20979, C1 => n14764, C2 =>
                           n20973, A => n16520, ZN => n16517);
   U17690 : AOI22_X1 port map( A1 => n20967, A2 => n8871, B1 => n20961, B2 => 
                           n18979, ZN => n16520);
   U17691 : OAI221_X1 port map( B1 => n14361, B2 => n21113, C1 => n14829, C2 =>
                           n21107, A => n16492, ZN => n16491);
   U17692 : AOI22_X1 port map( A1 => n21101, A2 => n18948, B1 => n21095, B2 => 
                           n18949, ZN => n16492);
   U17693 : OAI221_X1 port map( B1 => n15426, B2 => n21064, C1 => n16025, C2 =>
                           n21058, A => n16494, ZN => n16489);
   U17694 : AOI22_X1 port map( A1 => n21052, A2 => n9039, B1 => n21046, B2 => 
                           n8655, ZN => n16494);
   U17695 : OAI221_X1 port map( B1 => n15761, B2 => n20979, C1 => n14763, C2 =>
                           n20973, A => n16501, ZN => n16498);
   U17696 : AOI22_X1 port map( A1 => n20967, A2 => n8869, B1 => n20961, B2 => 
                           n18959, ZN => n16501);
   U17697 : OAI221_X1 port map( B1 => n14360, B2 => n21113, C1 => n14828, C2 =>
                           n21107, A => n16473, ZN => n16472);
   U17698 : AOI22_X1 port map( A1 => n21101, A2 => n18928, B1 => n21095, B2 => 
                           n18929, ZN => n16473);
   U17699 : OAI221_X1 port map( B1 => n15425, B2 => n21064, C1 => n16024, C2 =>
                           n21058, A => n16475, ZN => n16470);
   U17700 : AOI22_X1 port map( A1 => n21052, A2 => n9035, B1 => n21046, B2 => 
                           n8651, ZN => n16475);
   U17701 : OAI221_X1 port map( B1 => n15760, B2 => n20979, C1 => n14762, C2 =>
                           n20973, A => n16482, ZN => n16479);
   U17702 : AOI22_X1 port map( A1 => n20967, A2 => n8867, B1 => n20961, B2 => 
                           n18939, ZN => n16482);
   U17703 : OAI221_X1 port map( B1 => n14359, B2 => n21113, C1 => n14827, C2 =>
                           n21107, A => n16454, ZN => n16453);
   U17704 : AOI22_X1 port map( A1 => n21101, A2 => n18908, B1 => n21095, B2 => 
                           n18909, ZN => n16454);
   U17705 : OAI221_X1 port map( B1 => n15424, B2 => n21064, C1 => n16023, C2 =>
                           n21058, A => n16456, ZN => n16451);
   U17706 : AOI22_X1 port map( A1 => n21052, A2 => n9031, B1 => n21046, B2 => 
                           n8647, ZN => n16456);
   U17707 : OAI221_X1 port map( B1 => n15759, B2 => n20979, C1 => n14761, C2 =>
                           n20973, A => n16463, ZN => n16460);
   U17708 : AOI22_X1 port map( A1 => n20967, A2 => n8865, B1 => n20961, B2 => 
                           n18919, ZN => n16463);
   U17709 : OAI221_X1 port map( B1 => n14358, B2 => n21113, C1 => n14826, C2 =>
                           n21107, A => n16435, ZN => n16434);
   U17710 : AOI22_X1 port map( A1 => n21101, A2 => n18888, B1 => n21095, B2 => 
                           n18889, ZN => n16435);
   U17711 : OAI221_X1 port map( B1 => n15423, B2 => n21064, C1 => n16022, C2 =>
                           n21058, A => n16437, ZN => n16432);
   U17712 : AOI22_X1 port map( A1 => n21052, A2 => n9027, B1 => n21046, B2 => 
                           n8643, ZN => n16437);
   U17713 : OAI221_X1 port map( B1 => n15758, B2 => n20979, C1 => n14760, C2 =>
                           n20973, A => n16444, ZN => n16441);
   U17714 : AOI22_X1 port map( A1 => n20967, A2 => n8863, B1 => n20961, B2 => 
                           n18899, ZN => n16444);
   U17715 : OAI221_X1 port map( B1 => n14357, B2 => n21113, C1 => n14825, C2 =>
                           n21107, A => n16416, ZN => n16415);
   U17716 : AOI22_X1 port map( A1 => n21101, A2 => n18868, B1 => n21095, B2 => 
                           n18869, ZN => n16416);
   U17717 : OAI221_X1 port map( B1 => n15422, B2 => n21064, C1 => n16021, C2 =>
                           n21058, A => n16418, ZN => n16413);
   U17718 : AOI22_X1 port map( A1 => n21052, A2 => n9023, B1 => n21046, B2 => 
                           n8639, ZN => n16418);
   U17719 : OAI221_X1 port map( B1 => n15757, B2 => n20979, C1 => n14759, C2 =>
                           n20973, A => n16425, ZN => n16422);
   U17720 : AOI22_X1 port map( A1 => n20967, A2 => n8861, B1 => n20961, B2 => 
                           n18879, ZN => n16425);
   U17721 : OAI221_X1 port map( B1 => n14356, B2 => n21114, C1 => n14824, C2 =>
                           n21108, A => n16397, ZN => n16396);
   U17722 : AOI22_X1 port map( A1 => n21102, A2 => n18848, B1 => n21096, B2 => 
                           n18849, ZN => n16397);
   U17723 : OAI221_X1 port map( B1 => n15421, B2 => n21065, C1 => n16020, C2 =>
                           n21059, A => n16399, ZN => n16394);
   U17724 : AOI22_X1 port map( A1 => n21053, A2 => n9019, B1 => n21047, B2 => 
                           n8635, ZN => n16399);
   U17725 : OAI221_X1 port map( B1 => n15756, B2 => n20980, C1 => n14758, C2 =>
                           n20974, A => n16406, ZN => n16403);
   U17726 : AOI22_X1 port map( A1 => n20968, A2 => n8859, B1 => n20962, B2 => 
                           n18859, ZN => n16406);
   U17727 : OAI221_X1 port map( B1 => n14355, B2 => n21114, C1 => n14823, C2 =>
                           n21108, A => n16378, ZN => n16377);
   U17728 : AOI22_X1 port map( A1 => n21102, A2 => n18828, B1 => n21096, B2 => 
                           n18829, ZN => n16378);
   U17729 : OAI221_X1 port map( B1 => n15420, B2 => n21065, C1 => n16019, C2 =>
                           n21059, A => n16380, ZN => n16375);
   U17730 : AOI22_X1 port map( A1 => n21053, A2 => n9015, B1 => n21047, B2 => 
                           n8631, ZN => n16380);
   U17731 : OAI221_X1 port map( B1 => n15755, B2 => n20980, C1 => n14757, C2 =>
                           n20974, A => n16387, ZN => n16384);
   U17732 : AOI22_X1 port map( A1 => n20968, A2 => n8857, B1 => n20962, B2 => 
                           n18839, ZN => n16387);
   U17733 : OAI221_X1 port map( B1 => n14354, B2 => n21114, C1 => n14822, C2 =>
                           n21108, A => n16359, ZN => n16358);
   U17734 : AOI22_X1 port map( A1 => n21102, A2 => n18808, B1 => n21096, B2 => 
                           n18809, ZN => n16359);
   U17735 : OAI221_X1 port map( B1 => n15419, B2 => n21065, C1 => n16018, C2 =>
                           n21059, A => n16361, ZN => n16356);
   U17736 : AOI22_X1 port map( A1 => n21053, A2 => n9011, B1 => n21047, B2 => 
                           n8627, ZN => n16361);
   U17737 : OAI221_X1 port map( B1 => n15754, B2 => n20980, C1 => n14756, C2 =>
                           n20974, A => n16368, ZN => n16365);
   U17738 : AOI22_X1 port map( A1 => n20968, A2 => n8855, B1 => n20962, B2 => 
                           n18819, ZN => n16368);
   U17739 : OAI221_X1 port map( B1 => n14353, B2 => n21114, C1 => n14821, C2 =>
                           n21108, A => n16340, ZN => n16339);
   U17740 : AOI22_X1 port map( A1 => n21102, A2 => n18788, B1 => n21096, B2 => 
                           n18789, ZN => n16340);
   U17741 : OAI221_X1 port map( B1 => n15418, B2 => n21065, C1 => n16017, C2 =>
                           n21059, A => n16342, ZN => n16337);
   U17742 : AOI22_X1 port map( A1 => n21053, A2 => n9007, B1 => n21047, B2 => 
                           n8623, ZN => n16342);
   U17743 : OAI221_X1 port map( B1 => n15753, B2 => n20980, C1 => n14755, C2 =>
                           n20974, A => n16349, ZN => n16346);
   U17744 : AOI22_X1 port map( A1 => n20968, A2 => n8853, B1 => n20962, B2 => 
                           n18799, ZN => n16349);
   U17745 : OAI221_X1 port map( B1 => n14554, B2 => n21073, C1 => n14886, C2 =>
                           n21071, A => n16322, ZN => n16319);
   U17746 : AOI22_X1 port map( A1 => n18764, A2 => n21090, B1 => n21081, B2 => 
                           n18765, ZN => n16322);
   U17747 : OAI221_X1 port map( B1 => n14352, B2 => n21114, C1 => n14820, C2 =>
                           n21108, A => n16321, ZN => n16320);
   U17748 : AOI22_X1 port map( A1 => n21102, A2 => n18768, B1 => n21096, B2 => 
                           n18769, ZN => n16321);
   U17749 : OAI221_X1 port map( B1 => n15417, B2 => n21065, C1 => n16016, C2 =>
                           n21059, A => n16323, ZN => n16318);
   U17750 : AOI22_X1 port map( A1 => n21053, A2 => n9003, B1 => n21047, B2 => 
                           n8619, ZN => n16323);
   U17751 : OAI221_X1 port map( B1 => n15752, B2 => n20980, C1 => n14754, C2 =>
                           n20974, A => n16330, ZN => n16327);
   U17752 : AOI22_X1 port map( A1 => n20968, A2 => n8851, B1 => n20962, B2 => 
                           n18779, ZN => n16330);
   U17753 : OAI221_X1 port map( B1 => n14553, B2 => n21073, C1 => n14885, C2 =>
                           n21071, A => n16303, ZN => n16300);
   U17754 : AOI22_X1 port map( A1 => n18744, A2 => n21090, B1 => n21081, B2 => 
                           n18745, ZN => n16303);
   U17755 : OAI221_X1 port map( B1 => n14351, B2 => n21114, C1 => n14819, C2 =>
                           n21108, A => n16302, ZN => n16301);
   U17756 : AOI22_X1 port map( A1 => n21102, A2 => n18748, B1 => n21096, B2 => 
                           n18749, ZN => n16302);
   U17757 : OAI221_X1 port map( B1 => n15416, B2 => n21065, C1 => n16015, C2 =>
                           n21059, A => n16304, ZN => n16299);
   U17758 : AOI22_X1 port map( A1 => n21053, A2 => n8999, B1 => n21047, B2 => 
                           n8615, ZN => n16304);
   U17759 : OAI221_X1 port map( B1 => n15751, B2 => n20980, C1 => n14753, C2 =>
                           n20974, A => n16311, ZN => n16308);
   U17760 : AOI22_X1 port map( A1 => n20968, A2 => n8849, B1 => n20962, B2 => 
                           n18759, ZN => n16311);
   U17761 : OAI221_X1 port map( B1 => n14552, B2 => n21073, C1 => n14884, C2 =>
                           n21071, A => n16284, ZN => n16281);
   U17762 : AOI22_X1 port map( A1 => n18724, A2 => n21090, B1 => n21081, B2 => 
                           n18725, ZN => n16284);
   U17763 : OAI221_X1 port map( B1 => n14350, B2 => n21114, C1 => n14818, C2 =>
                           n21108, A => n16283, ZN => n16282);
   U17764 : AOI22_X1 port map( A1 => n21102, A2 => n18728, B1 => n21096, B2 => 
                           n18729, ZN => n16283);
   U17765 : OAI221_X1 port map( B1 => n15415, B2 => n21065, C1 => n16014, C2 =>
                           n21059, A => n16285, ZN => n16280);
   U17766 : AOI22_X1 port map( A1 => n21053, A2 => n8995, B1 => n21047, B2 => 
                           n8611, ZN => n16285);
   U17767 : OAI221_X1 port map( B1 => n15750, B2 => n20980, C1 => n14752, C2 =>
                           n20974, A => n16292, ZN => n16289);
   U17768 : AOI22_X1 port map( A1 => n20968, A2 => n8847, B1 => n20962, B2 => 
                           n18739, ZN => n16292);
   U17769 : OAI221_X1 port map( B1 => n14551, B2 => n21073, C1 => n14883, C2 =>
                           n21071, A => n16265, ZN => n16262);
   U17770 : AOI22_X1 port map( A1 => n18704, A2 => n21090, B1 => n21081, B2 => 
                           n18705, ZN => n16265);
   U17771 : OAI221_X1 port map( B1 => n14349, B2 => n21114, C1 => n14817, C2 =>
                           n21108, A => n16264, ZN => n16263);
   U17772 : AOI22_X1 port map( A1 => n21102, A2 => n18708, B1 => n21096, B2 => 
                           n18709, ZN => n16264);
   U17773 : OAI221_X1 port map( B1 => n15414, B2 => n21065, C1 => n16013, C2 =>
                           n21059, A => n16266, ZN => n16261);
   U17774 : AOI22_X1 port map( A1 => n21053, A2 => n8991, B1 => n21047, B2 => 
                           n8607, ZN => n16266);
   U17775 : OAI221_X1 port map( B1 => n15749, B2 => n20980, C1 => n14751, C2 =>
                           n20974, A => n16273, ZN => n16270);
   U17776 : AOI22_X1 port map( A1 => n20968, A2 => n8845, B1 => n20962, B2 => 
                           n18719, ZN => n16273);
   U17777 : OAI221_X1 port map( B1 => n14550, B2 => n21073, C1 => n14882, C2 =>
                           n21071, A => n16246, ZN => n16243);
   U17778 : AOI22_X1 port map( A1 => n18684, A2 => n21090, B1 => n21081, B2 => 
                           n18685, ZN => n16246);
   U17779 : OAI221_X1 port map( B1 => n14348, B2 => n21114, C1 => n14816, C2 =>
                           n21108, A => n16245, ZN => n16244);
   U17780 : AOI22_X1 port map( A1 => n21102, A2 => n18688, B1 => n21096, B2 => 
                           n18689, ZN => n16245);
   U17781 : OAI221_X1 port map( B1 => n15413, B2 => n21065, C1 => n16012, C2 =>
                           n21059, A => n16247, ZN => n16242);
   U17782 : AOI22_X1 port map( A1 => n21053, A2 => n8987, B1 => n21047, B2 => 
                           n8603, ZN => n16247);
   U17783 : OAI221_X1 port map( B1 => n15748, B2 => n20980, C1 => n14750, C2 =>
                           n20974, A => n16254, ZN => n16251);
   U17784 : AOI22_X1 port map( A1 => n20968, A2 => n8843, B1 => n20962, B2 => 
                           n18699, ZN => n16254);
   U17785 : OAI221_X1 port map( B1 => n14549, B2 => n21073, C1 => n14881, C2 =>
                           n21071, A => n16227, ZN => n16224);
   U17786 : AOI22_X1 port map( A1 => n18664, A2 => n21090, B1 => n21081, B2 => 
                           n18665, ZN => n16227);
   U17787 : OAI221_X1 port map( B1 => n14347, B2 => n21114, C1 => n14815, C2 =>
                           n21108, A => n16226, ZN => n16225);
   U17788 : AOI22_X1 port map( A1 => n21102, A2 => n18668, B1 => n21096, B2 => 
                           n18669, ZN => n16226);
   U17789 : OAI221_X1 port map( B1 => n15412, B2 => n21065, C1 => n16011, C2 =>
                           n21059, A => n16228, ZN => n16223);
   U17790 : AOI22_X1 port map( A1 => n21053, A2 => n8983, B1 => n21047, B2 => 
                           n8599, ZN => n16228);
   U17791 : OAI221_X1 port map( B1 => n15747, B2 => n20980, C1 => n14749, C2 =>
                           n20974, A => n16235, ZN => n16232);
   U17792 : AOI22_X1 port map( A1 => n20968, A2 => n8841, B1 => n20962, B2 => 
                           n18679, ZN => n16235);
   U17793 : OAI221_X1 port map( B1 => n14548, B2 => n21073, C1 => n14880, C2 =>
                           n21071, A => n16208, ZN => n16205);
   U17794 : AOI22_X1 port map( A1 => n18644, A2 => n21090, B1 => n21081, B2 => 
                           n18645, ZN => n16208);
   U17795 : OAI221_X1 port map( B1 => n14346, B2 => n21114, C1 => n14814, C2 =>
                           n21108, A => n16207, ZN => n16206);
   U17796 : AOI22_X1 port map( A1 => n21102, A2 => n18648, B1 => n21096, B2 => 
                           n18649, ZN => n16207);
   U17797 : OAI221_X1 port map( B1 => n15411, B2 => n21065, C1 => n16010, C2 =>
                           n21059, A => n16209, ZN => n16204);
   U17798 : AOI22_X1 port map( A1 => n21053, A2 => n8979, B1 => n21047, B2 => 
                           n8595, ZN => n16209);
   U17799 : OAI221_X1 port map( B1 => n15746, B2 => n20980, C1 => n14748, C2 =>
                           n20974, A => n16216, ZN => n16213);
   U17800 : AOI22_X1 port map( A1 => n20968, A2 => n8839, B1 => n20962, B2 => 
                           n18659, ZN => n16216);
   U17801 : OAI221_X1 port map( B1 => n14547, B2 => n21073, C1 => n14879, C2 =>
                           n21071, A => n16189, ZN => n16186);
   U17802 : AOI22_X1 port map( A1 => n18624, A2 => n21090, B1 => n21081, B2 => 
                           n18625, ZN => n16189);
   U17803 : OAI221_X1 port map( B1 => n14345, B2 => n21114, C1 => n14813, C2 =>
                           n21108, A => n16188, ZN => n16187);
   U17804 : AOI22_X1 port map( A1 => n21102, A2 => n18628, B1 => n21096, B2 => 
                           n18629, ZN => n16188);
   U17805 : OAI221_X1 port map( B1 => n15410, B2 => n21065, C1 => n16009, C2 =>
                           n21059, A => n16190, ZN => n16185);
   U17806 : AOI22_X1 port map( A1 => n21053, A2 => n8975, B1 => n21047, B2 => 
                           n8591, ZN => n16190);
   U17807 : OAI221_X1 port map( B1 => n15745, B2 => n20980, C1 => n14747, C2 =>
                           n20974, A => n16197, ZN => n16194);
   U17808 : AOI22_X1 port map( A1 => n20968, A2 => n8837, B1 => n20962, B2 => 
                           n18639, ZN => n16197);
   U17809 : OAI221_X1 port map( B1 => n14344, B2 => n21115, C1 => n14812, C2 =>
                           n21109, A => n16169, ZN => n16168);
   U17810 : AOI22_X1 port map( A1 => n21103, A2 => n18608, B1 => n21097, B2 => 
                           n18609, ZN => n16169);
   U17811 : OAI221_X1 port map( B1 => n14343, B2 => n21115, C1 => n14811, C2 =>
                           n21109, A => n16150, ZN => n16149);
   U17812 : AOI22_X1 port map( A1 => n21103, A2 => n18588, B1 => n21097, B2 => 
                           n18589, ZN => n16150);
   U17813 : OAI221_X1 port map( B1 => n14342, B2 => n21115, C1 => n14810, C2 =>
                           n21109, A => n16131, ZN => n16130);
   U17814 : AOI22_X1 port map( A1 => n21103, A2 => n18568, B1 => n21097, B2 => 
                           n18569, ZN => n16131);
   U17815 : OAI22_X1 port map( A1 => n21150, A2 => n16002, B1 => n21528, B2 => 
                           n21142, ZN => n5501);
   U17816 : OAI22_X1 port map( A1 => n21150, A2 => n16001, B1 => n21531, B2 => 
                           n21142, ZN => n5502);
   U17817 : OAI22_X1 port map( A1 => n21150, A2 => n16000, B1 => n21534, B2 => 
                           n21142, ZN => n5503);
   U17818 : OAI22_X1 port map( A1 => n21150, A2 => n15999, B1 => n21537, B2 => 
                           n21142, ZN => n5504);
   U17819 : OAI22_X1 port map( A1 => n21150, A2 => n15998, B1 => n21540, B2 => 
                           n21142, ZN => n5505);
   U17820 : OAI22_X1 port map( A1 => n21150, A2 => n15997, B1 => n21543, B2 => 
                           n21142, ZN => n5506);
   U17821 : OAI22_X1 port map( A1 => n21150, A2 => n15996, B1 => n21546, B2 => 
                           n21142, ZN => n5507);
   U17822 : OAI22_X1 port map( A1 => n21150, A2 => n15995, B1 => n21549, B2 => 
                           n21142, ZN => n5508);
   U17823 : OAI22_X1 port map( A1 => n21150, A2 => n15994, B1 => n21552, B2 => 
                           n21142, ZN => n5509);
   U17824 : OAI22_X1 port map( A1 => n21150, A2 => n15993, B1 => n21555, B2 => 
                           n21142, ZN => n5510);
   U17825 : OAI22_X1 port map( A1 => n21150, A2 => n15992, B1 => n21558, B2 => 
                           n21142, ZN => n5511);
   U17826 : OAI22_X1 port map( A1 => n21150, A2 => n15991, B1 => n21561, B2 => 
                           n21142, ZN => n5512);
   U17827 : OAI22_X1 port map( A1 => n21151, A2 => n15990, B1 => n21564, B2 => 
                           n21143, ZN => n5513);
   U17828 : OAI22_X1 port map( A1 => n21151, A2 => n15989, B1 => n21567, B2 => 
                           n21143, ZN => n5514);
   U17829 : OAI22_X1 port map( A1 => n21151, A2 => n15988, B1 => n21570, B2 => 
                           n21143, ZN => n5515);
   U17830 : OAI22_X1 port map( A1 => n21151, A2 => n15987, B1 => n21573, B2 => 
                           n21143, ZN => n5516);
   U17831 : OAI22_X1 port map( A1 => n21151, A2 => n15986, B1 => n21576, B2 => 
                           n21143, ZN => n5517);
   U17832 : OAI22_X1 port map( A1 => n21151, A2 => n15985, B1 => n21579, B2 => 
                           n21143, ZN => n5518);
   U17833 : OAI22_X1 port map( A1 => n21151, A2 => n15984, B1 => n21582, B2 => 
                           n21143, ZN => n5519);
   U17834 : OAI22_X1 port map( A1 => n21151, A2 => n15983, B1 => n21585, B2 => 
                           n21143, ZN => n5520);
   U17835 : OAI22_X1 port map( A1 => n21151, A2 => n15982, B1 => n21588, B2 => 
                           n21143, ZN => n5521);
   U17836 : OAI22_X1 port map( A1 => n21151, A2 => n15981, B1 => n21591, B2 => 
                           n21143, ZN => n5522);
   U17837 : OAI22_X1 port map( A1 => n21151, A2 => n15980, B1 => n21594, B2 => 
                           n21143, ZN => n5523);
   U17838 : OAI22_X1 port map( A1 => n21151, A2 => n15979, B1 => n21597, B2 => 
                           n21143, ZN => n5524);
   U17839 : OAI22_X1 port map( A1 => n21151, A2 => n15978, B1 => n21600, B2 => 
                           n21144, ZN => n5525);
   U17840 : OAI22_X1 port map( A1 => n21152, A2 => n15977, B1 => n21603, B2 => 
                           n21144, ZN => n5526);
   U17841 : OAI22_X1 port map( A1 => n21152, A2 => n15976, B1 => n21606, B2 => 
                           n21144, ZN => n5527);
   U17842 : OAI22_X1 port map( A1 => n21152, A2 => n15975, B1 => n21609, B2 => 
                           n21144, ZN => n5528);
   U17843 : OAI22_X1 port map( A1 => n21152, A2 => n15974, B1 => n21612, B2 => 
                           n21144, ZN => n5529);
   U17844 : OAI22_X1 port map( A1 => n21152, A2 => n15973, B1 => n21615, B2 => 
                           n21144, ZN => n5530);
   U17845 : OAI22_X1 port map( A1 => n21152, A2 => n15972, B1 => n21618, B2 => 
                           n21144, ZN => n5531);
   U17846 : OAI22_X1 port map( A1 => n21152, A2 => n15971, B1 => n21621, B2 => 
                           n21144, ZN => n5532);
   U17847 : OAI22_X1 port map( A1 => n21152, A2 => n15970, B1 => n21624, B2 => 
                           n21144, ZN => n5533);
   U17848 : OAI22_X1 port map( A1 => n21152, A2 => n15969, B1 => n21627, B2 => 
                           n21144, ZN => n5534);
   U17849 : OAI22_X1 port map( A1 => n21152, A2 => n15968, B1 => n21630, B2 => 
                           n21144, ZN => n5535);
   U17850 : OAI22_X1 port map( A1 => n21152, A2 => n15967, B1 => n21633, B2 => 
                           n21144, ZN => n5536);
   U17851 : OAI22_X1 port map( A1 => n21152, A2 => n15966, B1 => n21636, B2 => 
                           n21145, ZN => n5537);
   U17852 : OAI22_X1 port map( A1 => n21152, A2 => n15965, B1 => n21639, B2 => 
                           n21145, ZN => n5538);
   U17853 : OAI22_X1 port map( A1 => n21153, A2 => n15964, B1 => n21642, B2 => 
                           n21145, ZN => n5539);
   U17854 : OAI22_X1 port map( A1 => n21153, A2 => n15963, B1 => n21645, B2 => 
                           n21145, ZN => n5540);
   U17855 : OAI22_X1 port map( A1 => n21153, A2 => n15962, B1 => n21648, B2 => 
                           n21145, ZN => n5541);
   U17856 : OAI22_X1 port map( A1 => n21153, A2 => n15961, B1 => n21651, B2 => 
                           n21145, ZN => n5542);
   U17857 : OAI22_X1 port map( A1 => n21153, A2 => n15960, B1 => n21654, B2 => 
                           n21145, ZN => n5543);
   U17858 : OAI22_X1 port map( A1 => n21153, A2 => n15959, B1 => n21657, B2 => 
                           n21145, ZN => n5544);
   U17859 : OAI22_X1 port map( A1 => n21153, A2 => n15958, B1 => n21660, B2 => 
                           n21145, ZN => n5545);
   U17860 : OAI22_X1 port map( A1 => n21153, A2 => n15957, B1 => n21663, B2 => 
                           n21145, ZN => n5546);
   U17861 : OAI22_X1 port map( A1 => n21153, A2 => n15956, B1 => n21666, B2 => 
                           n21145, ZN => n5547);
   U17862 : OAI22_X1 port map( A1 => n21153, A2 => n15955, B1 => n21669, B2 => 
                           n21145, ZN => n5548);
   U17863 : OAI22_X1 port map( A1 => n21153, A2 => n15954, B1 => n21672, B2 => 
                           n21146, ZN => n5549);
   U17864 : OAI22_X1 port map( A1 => n21153, A2 => n15953, B1 => n21675, B2 => 
                           n21146, ZN => n5550);
   U17865 : OAI22_X1 port map( A1 => n21153, A2 => n15952, B1 => n21678, B2 => 
                           n21146, ZN => n5551);
   U17866 : OAI22_X1 port map( A1 => n21154, A2 => n15951, B1 => n21681, B2 => 
                           n21146, ZN => n5552);
   U17867 : OAI22_X1 port map( A1 => n21154, A2 => n15950, B1 => n21684, B2 => 
                           n21146, ZN => n5553);
   U17868 : OAI22_X1 port map( A1 => n21154, A2 => n15949, B1 => n21687, B2 => 
                           n21146, ZN => n5554);
   U17869 : OAI22_X1 port map( A1 => n21154, A2 => n15948, B1 => n21690, B2 => 
                           n21146, ZN => n5555);
   U17870 : OAI22_X1 port map( A1 => n21154, A2 => n15947, B1 => n21693, B2 => 
                           n21146, ZN => n5556);
   U17871 : OAI22_X1 port map( A1 => n21154, A2 => n15946, B1 => n21696, B2 => 
                           n21146, ZN => n5557);
   U17872 : OAI22_X1 port map( A1 => n21154, A2 => n15945, B1 => n21699, B2 => 
                           n21146, ZN => n5558);
   U17873 : OAI22_X1 port map( A1 => n21154, A2 => n15944, B1 => n21702, B2 => 
                           n21146, ZN => n5559);
   U17874 : OAI22_X1 port map( A1 => n21154, A2 => n15943, B1 => n21705, B2 => 
                           n21146, ZN => n5560);
   U17875 : OAI22_X1 port map( A1 => n21176, A2 => n15870, B1 => n21528, B2 => 
                           n21168, ZN => n5629);
   U17876 : OAI22_X1 port map( A1 => n21176, A2 => n15869, B1 => n21531, B2 => 
                           n21168, ZN => n5630);
   U17877 : OAI22_X1 port map( A1 => n21176, A2 => n15868, B1 => n21534, B2 => 
                           n21168, ZN => n5631);
   U17878 : OAI22_X1 port map( A1 => n21176, A2 => n15867, B1 => n21537, B2 => 
                           n21168, ZN => n5632);
   U17879 : OAI22_X1 port map( A1 => n21176, A2 => n15866, B1 => n21540, B2 => 
                           n21168, ZN => n5633);
   U17880 : OAI22_X1 port map( A1 => n21176, A2 => n15865, B1 => n21543, B2 => 
                           n21168, ZN => n5634);
   U17881 : OAI22_X1 port map( A1 => n21176, A2 => n15864, B1 => n21546, B2 => 
                           n21168, ZN => n5635);
   U17882 : OAI22_X1 port map( A1 => n21176, A2 => n15863, B1 => n21549, B2 => 
                           n21168, ZN => n5636);
   U17883 : OAI22_X1 port map( A1 => n21176, A2 => n15862, B1 => n21552, B2 => 
                           n21168, ZN => n5637);
   U17884 : OAI22_X1 port map( A1 => n21176, A2 => n15861, B1 => n21555, B2 => 
                           n21168, ZN => n5638);
   U17885 : OAI22_X1 port map( A1 => n21176, A2 => n15860, B1 => n21558, B2 => 
                           n21168, ZN => n5639);
   U17886 : OAI22_X1 port map( A1 => n21176, A2 => n15859, B1 => n21561, B2 => 
                           n21168, ZN => n5640);
   U17887 : OAI22_X1 port map( A1 => n21177, A2 => n15858, B1 => n21564, B2 => 
                           n21169, ZN => n5641);
   U17888 : OAI22_X1 port map( A1 => n21177, A2 => n15857, B1 => n21567, B2 => 
                           n21169, ZN => n5642);
   U17889 : OAI22_X1 port map( A1 => n21177, A2 => n15856, B1 => n21570, B2 => 
                           n21169, ZN => n5643);
   U17890 : OAI22_X1 port map( A1 => n21177, A2 => n15855, B1 => n21573, B2 => 
                           n21169, ZN => n5644);
   U17891 : OAI22_X1 port map( A1 => n21177, A2 => n15854, B1 => n21576, B2 => 
                           n21169, ZN => n5645);
   U17892 : OAI22_X1 port map( A1 => n21177, A2 => n15853, B1 => n21579, B2 => 
                           n21169, ZN => n5646);
   U17893 : OAI22_X1 port map( A1 => n21177, A2 => n15852, B1 => n21582, B2 => 
                           n21169, ZN => n5647);
   U17894 : OAI22_X1 port map( A1 => n21177, A2 => n15851, B1 => n21585, B2 => 
                           n21169, ZN => n5648);
   U17895 : OAI22_X1 port map( A1 => n21177, A2 => n15850, B1 => n21588, B2 => 
                           n21169, ZN => n5649);
   U17896 : OAI22_X1 port map( A1 => n21177, A2 => n15849, B1 => n21591, B2 => 
                           n21169, ZN => n5650);
   U17897 : OAI22_X1 port map( A1 => n21177, A2 => n15848, B1 => n21594, B2 => 
                           n21169, ZN => n5651);
   U17898 : OAI22_X1 port map( A1 => n21177, A2 => n15847, B1 => n21597, B2 => 
                           n21169, ZN => n5652);
   U17899 : OAI22_X1 port map( A1 => n21177, A2 => n15846, B1 => n21600, B2 => 
                           n21170, ZN => n5653);
   U17900 : OAI22_X1 port map( A1 => n21178, A2 => n15845, B1 => n21603, B2 => 
                           n21170, ZN => n5654);
   U17901 : OAI22_X1 port map( A1 => n21178, A2 => n15844, B1 => n21606, B2 => 
                           n21170, ZN => n5655);
   U17902 : OAI22_X1 port map( A1 => n21178, A2 => n15843, B1 => n21609, B2 => 
                           n21170, ZN => n5656);
   U17903 : OAI22_X1 port map( A1 => n21178, A2 => n15842, B1 => n21612, B2 => 
                           n21170, ZN => n5657);
   U17904 : OAI22_X1 port map( A1 => n21178, A2 => n15841, B1 => n21615, B2 => 
                           n21170, ZN => n5658);
   U17905 : OAI22_X1 port map( A1 => n21178, A2 => n15840, B1 => n21618, B2 => 
                           n21170, ZN => n5659);
   U17906 : OAI22_X1 port map( A1 => n21178, A2 => n15839, B1 => n21621, B2 => 
                           n21170, ZN => n5660);
   U17907 : OAI22_X1 port map( A1 => n21178, A2 => n15838, B1 => n21624, B2 => 
                           n21170, ZN => n5661);
   U17908 : OAI22_X1 port map( A1 => n21178, A2 => n15837, B1 => n21627, B2 => 
                           n21170, ZN => n5662);
   U17909 : OAI22_X1 port map( A1 => n21178, A2 => n15836, B1 => n21630, B2 => 
                           n21170, ZN => n5663);
   U17910 : OAI22_X1 port map( A1 => n21178, A2 => n15835, B1 => n21633, B2 => 
                           n21170, ZN => n5664);
   U17911 : OAI22_X1 port map( A1 => n21178, A2 => n15834, B1 => n21636, B2 => 
                           n21171, ZN => n5665);
   U17912 : OAI22_X1 port map( A1 => n21178, A2 => n15833, B1 => n21639, B2 => 
                           n21171, ZN => n5666);
   U17913 : OAI22_X1 port map( A1 => n21179, A2 => n15832, B1 => n21642, B2 => 
                           n21171, ZN => n5667);
   U17914 : OAI22_X1 port map( A1 => n21179, A2 => n15831, B1 => n21645, B2 => 
                           n21171, ZN => n5668);
   U17915 : OAI22_X1 port map( A1 => n21179, A2 => n15830, B1 => n21648, B2 => 
                           n21171, ZN => n5669);
   U17916 : OAI22_X1 port map( A1 => n21179, A2 => n15829, B1 => n21651, B2 => 
                           n21171, ZN => n5670);
   U17917 : OAI22_X1 port map( A1 => n21179, A2 => n15828, B1 => n21654, B2 => 
                           n21171, ZN => n5671);
   U17918 : OAI22_X1 port map( A1 => n21179, A2 => n15827, B1 => n21657, B2 => 
                           n21171, ZN => n5672);
   U17919 : OAI22_X1 port map( A1 => n21179, A2 => n15826, B1 => n21660, B2 => 
                           n21171, ZN => n5673);
   U17920 : OAI22_X1 port map( A1 => n21179, A2 => n15825, B1 => n21663, B2 => 
                           n21171, ZN => n5674);
   U17921 : OAI22_X1 port map( A1 => n21179, A2 => n15824, B1 => n21666, B2 => 
                           n21171, ZN => n5675);
   U17922 : OAI22_X1 port map( A1 => n21179, A2 => n15823, B1 => n21669, B2 => 
                           n21171, ZN => n5676);
   U17923 : OAI22_X1 port map( A1 => n21179, A2 => n15822, B1 => n21672, B2 => 
                           n21172, ZN => n5677);
   U17924 : OAI22_X1 port map( A1 => n21179, A2 => n15821, B1 => n21675, B2 => 
                           n21172, ZN => n5678);
   U17925 : OAI22_X1 port map( A1 => n21179, A2 => n15820, B1 => n21678, B2 => 
                           n21172, ZN => n5679);
   U17926 : OAI22_X1 port map( A1 => n21180, A2 => n15819, B1 => n21681, B2 => 
                           n21172, ZN => n5680);
   U17927 : OAI22_X1 port map( A1 => n21180, A2 => n15818, B1 => n21684, B2 => 
                           n21172, ZN => n5681);
   U17928 : OAI22_X1 port map( A1 => n21180, A2 => n15817, B1 => n21687, B2 => 
                           n21172, ZN => n5682);
   U17929 : OAI22_X1 port map( A1 => n21180, A2 => n15816, B1 => n21690, B2 => 
                           n21172, ZN => n5683);
   U17930 : OAI22_X1 port map( A1 => n21180, A2 => n15815, B1 => n21693, B2 => 
                           n21172, ZN => n5684);
   U17931 : OAI22_X1 port map( A1 => n21180, A2 => n15814, B1 => n21696, B2 => 
                           n21172, ZN => n5685);
   U17932 : OAI22_X1 port map( A1 => n21180, A2 => n15813, B1 => n21699, B2 => 
                           n21172, ZN => n5686);
   U17933 : OAI22_X1 port map( A1 => n21180, A2 => n15812, B1 => n21702, B2 => 
                           n21172, ZN => n5687);
   U17934 : OAI22_X1 port map( A1 => n21180, A2 => n15811, B1 => n21705, B2 => 
                           n21172, ZN => n5688);
   U17935 : OAI22_X1 port map( A1 => n21202, A2 => n15735, B1 => n21528, B2 => 
                           n21194, ZN => n5757);
   U17936 : OAI22_X1 port map( A1 => n21202, A2 => n15734, B1 => n21531, B2 => 
                           n21194, ZN => n5758);
   U17937 : OAI22_X1 port map( A1 => n21202, A2 => n15733, B1 => n21534, B2 => 
                           n21194, ZN => n5759);
   U17938 : OAI22_X1 port map( A1 => n21202, A2 => n15732, B1 => n21537, B2 => 
                           n21194, ZN => n5760);
   U17939 : OAI22_X1 port map( A1 => n21202, A2 => n15731, B1 => n21540, B2 => 
                           n21194, ZN => n5761);
   U17940 : OAI22_X1 port map( A1 => n21202, A2 => n15730, B1 => n21543, B2 => 
                           n21194, ZN => n5762);
   U17941 : OAI22_X1 port map( A1 => n21202, A2 => n15729, B1 => n21546, B2 => 
                           n21194, ZN => n5763);
   U17942 : OAI22_X1 port map( A1 => n21202, A2 => n15728, B1 => n21549, B2 => 
                           n21194, ZN => n5764);
   U17943 : OAI22_X1 port map( A1 => n21202, A2 => n15727, B1 => n21552, B2 => 
                           n21194, ZN => n5765);
   U17944 : OAI22_X1 port map( A1 => n21202, A2 => n15726, B1 => n21555, B2 => 
                           n21194, ZN => n5766);
   U17945 : OAI22_X1 port map( A1 => n21202, A2 => n15725, B1 => n21558, B2 => 
                           n21194, ZN => n5767);
   U17946 : OAI22_X1 port map( A1 => n21202, A2 => n15724, B1 => n21561, B2 => 
                           n21194, ZN => n5768);
   U17947 : OAI22_X1 port map( A1 => n21203, A2 => n15723, B1 => n21564, B2 => 
                           n21195, ZN => n5769);
   U17948 : OAI22_X1 port map( A1 => n21203, A2 => n15722, B1 => n21567, B2 => 
                           n21195, ZN => n5770);
   U17949 : OAI22_X1 port map( A1 => n21203, A2 => n15721, B1 => n21570, B2 => 
                           n21195, ZN => n5771);
   U17950 : OAI22_X1 port map( A1 => n21203, A2 => n15720, B1 => n21573, B2 => 
                           n21195, ZN => n5772);
   U17951 : OAI22_X1 port map( A1 => n21203, A2 => n15719, B1 => n21576, B2 => 
                           n21195, ZN => n5773);
   U17952 : OAI22_X1 port map( A1 => n21203, A2 => n15718, B1 => n21579, B2 => 
                           n21195, ZN => n5774);
   U17953 : OAI22_X1 port map( A1 => n21203, A2 => n15717, B1 => n21582, B2 => 
                           n21195, ZN => n5775);
   U17954 : OAI22_X1 port map( A1 => n21203, A2 => n15716, B1 => n21585, B2 => 
                           n21195, ZN => n5776);
   U17955 : OAI22_X1 port map( A1 => n21203, A2 => n15715, B1 => n21588, B2 => 
                           n21195, ZN => n5777);
   U17956 : OAI22_X1 port map( A1 => n21203, A2 => n15714, B1 => n21591, B2 => 
                           n21195, ZN => n5778);
   U17957 : OAI22_X1 port map( A1 => n21203, A2 => n15713, B1 => n21594, B2 => 
                           n21195, ZN => n5779);
   U17958 : OAI22_X1 port map( A1 => n21203, A2 => n15712, B1 => n21597, B2 => 
                           n21195, ZN => n5780);
   U17959 : OAI22_X1 port map( A1 => n21203, A2 => n15711, B1 => n21600, B2 => 
                           n21196, ZN => n5781);
   U17960 : OAI22_X1 port map( A1 => n21204, A2 => n15710, B1 => n21603, B2 => 
                           n21196, ZN => n5782);
   U17961 : OAI22_X1 port map( A1 => n21204, A2 => n15709, B1 => n21606, B2 => 
                           n21196, ZN => n5783);
   U17962 : OAI22_X1 port map( A1 => n21204, A2 => n15708, B1 => n21609, B2 => 
                           n21196, ZN => n5784);
   U17963 : OAI22_X1 port map( A1 => n21204, A2 => n15707, B1 => n21612, B2 => 
                           n21196, ZN => n5785);
   U17964 : OAI22_X1 port map( A1 => n21204, A2 => n15706, B1 => n21615, B2 => 
                           n21196, ZN => n5786);
   U17965 : OAI22_X1 port map( A1 => n21204, A2 => n15705, B1 => n21618, B2 => 
                           n21196, ZN => n5787);
   U17966 : OAI22_X1 port map( A1 => n21204, A2 => n15704, B1 => n21621, B2 => 
                           n21196, ZN => n5788);
   U17967 : OAI22_X1 port map( A1 => n21204, A2 => n15703, B1 => n21624, B2 => 
                           n21196, ZN => n5789);
   U17968 : OAI22_X1 port map( A1 => n21204, A2 => n15702, B1 => n21627, B2 => 
                           n21196, ZN => n5790);
   U17969 : OAI22_X1 port map( A1 => n21204, A2 => n15701, B1 => n21630, B2 => 
                           n21196, ZN => n5791);
   U17970 : OAI22_X1 port map( A1 => n21204, A2 => n15700, B1 => n21633, B2 => 
                           n21196, ZN => n5792);
   U17971 : OAI22_X1 port map( A1 => n21204, A2 => n15699, B1 => n21636, B2 => 
                           n21197, ZN => n5793);
   U17972 : OAI22_X1 port map( A1 => n21204, A2 => n15698, B1 => n21639, B2 => 
                           n21197, ZN => n5794);
   U17973 : OAI22_X1 port map( A1 => n21205, A2 => n15697, B1 => n21642, B2 => 
                           n21197, ZN => n5795);
   U17974 : OAI22_X1 port map( A1 => n21205, A2 => n15696, B1 => n21645, B2 => 
                           n21197, ZN => n5796);
   U17975 : OAI22_X1 port map( A1 => n21205, A2 => n15695, B1 => n21648, B2 => 
                           n21197, ZN => n5797);
   U17976 : OAI22_X1 port map( A1 => n21205, A2 => n15694, B1 => n21651, B2 => 
                           n21197, ZN => n5798);
   U17977 : OAI22_X1 port map( A1 => n21205, A2 => n15693, B1 => n21654, B2 => 
                           n21197, ZN => n5799);
   U17978 : OAI22_X1 port map( A1 => n21205, A2 => n15692, B1 => n21657, B2 => 
                           n21197, ZN => n5800);
   U17979 : OAI22_X1 port map( A1 => n21205, A2 => n15691, B1 => n21660, B2 => 
                           n21197, ZN => n5801);
   U17980 : OAI22_X1 port map( A1 => n21205, A2 => n15690, B1 => n21663, B2 => 
                           n21197, ZN => n5802);
   U17981 : OAI22_X1 port map( A1 => n21205, A2 => n15689, B1 => n21666, B2 => 
                           n21197, ZN => n5803);
   U17982 : OAI22_X1 port map( A1 => n21205, A2 => n15688, B1 => n21669, B2 => 
                           n21197, ZN => n5804);
   U17983 : OAI22_X1 port map( A1 => n21205, A2 => n15687, B1 => n21672, B2 => 
                           n21198, ZN => n5805);
   U17984 : OAI22_X1 port map( A1 => n21205, A2 => n15686, B1 => n21675, B2 => 
                           n21198, ZN => n5806);
   U17985 : OAI22_X1 port map( A1 => n21205, A2 => n15685, B1 => n21678, B2 => 
                           n21198, ZN => n5807);
   U17986 : OAI22_X1 port map( A1 => n21206, A2 => n15684, B1 => n21681, B2 => 
                           n21198, ZN => n5808);
   U17987 : OAI22_X1 port map( A1 => n21206, A2 => n15683, B1 => n21684, B2 => 
                           n21198, ZN => n5809);
   U17988 : OAI22_X1 port map( A1 => n21206, A2 => n15682, B1 => n21687, B2 => 
                           n21198, ZN => n5810);
   U17989 : OAI22_X1 port map( A1 => n21206, A2 => n15681, B1 => n21690, B2 => 
                           n21198, ZN => n5811);
   U17990 : OAI22_X1 port map( A1 => n21206, A2 => n15680, B1 => n21693, B2 => 
                           n21198, ZN => n5812);
   U17991 : OAI22_X1 port map( A1 => n21206, A2 => n15679, B1 => n21696, B2 => 
                           n21198, ZN => n5813);
   U17992 : OAI22_X1 port map( A1 => n21206, A2 => n15678, B1 => n21699, B2 => 
                           n21198, ZN => n5814);
   U17993 : OAI22_X1 port map( A1 => n21206, A2 => n15677, B1 => n21702, B2 => 
                           n21198, ZN => n5815);
   U17994 : OAI22_X1 port map( A1 => n21206, A2 => n15676, B1 => n21705, B2 => 
                           n21198, ZN => n5816);
   U17995 : OAI22_X1 port map( A1 => n21228, A2 => n15602, B1 => n21527, B2 => 
                           n21220, ZN => n5885);
   U17996 : OAI22_X1 port map( A1 => n21228, A2 => n15601, B1 => n21530, B2 => 
                           n21220, ZN => n5886);
   U17997 : OAI22_X1 port map( A1 => n21228, A2 => n15600, B1 => n21533, B2 => 
                           n21220, ZN => n5887);
   U17998 : OAI22_X1 port map( A1 => n21228, A2 => n15599, B1 => n21536, B2 => 
                           n21220, ZN => n5888);
   U17999 : OAI22_X1 port map( A1 => n21228, A2 => n15598, B1 => n21539, B2 => 
                           n21220, ZN => n5889);
   U18000 : OAI22_X1 port map( A1 => n21228, A2 => n15597, B1 => n21542, B2 => 
                           n21220, ZN => n5890);
   U18001 : OAI22_X1 port map( A1 => n21228, A2 => n15596, B1 => n21545, B2 => 
                           n21220, ZN => n5891);
   U18002 : OAI22_X1 port map( A1 => n21228, A2 => n15595, B1 => n21548, B2 => 
                           n21220, ZN => n5892);
   U18003 : OAI22_X1 port map( A1 => n21228, A2 => n15594, B1 => n21551, B2 => 
                           n21220, ZN => n5893);
   U18004 : OAI22_X1 port map( A1 => n21228, A2 => n15593, B1 => n21554, B2 => 
                           n21220, ZN => n5894);
   U18005 : OAI22_X1 port map( A1 => n21228, A2 => n15592, B1 => n21557, B2 => 
                           n21220, ZN => n5895);
   U18006 : OAI22_X1 port map( A1 => n21228, A2 => n15591, B1 => n21560, B2 => 
                           n21220, ZN => n5896);
   U18007 : OAI22_X1 port map( A1 => n21229, A2 => n15590, B1 => n21563, B2 => 
                           n21221, ZN => n5897);
   U18008 : OAI22_X1 port map( A1 => n21229, A2 => n15589, B1 => n21566, B2 => 
                           n21221, ZN => n5898);
   U18009 : OAI22_X1 port map( A1 => n21229, A2 => n15588, B1 => n21569, B2 => 
                           n21221, ZN => n5899);
   U18010 : OAI22_X1 port map( A1 => n21229, A2 => n15587, B1 => n21572, B2 => 
                           n21221, ZN => n5900);
   U18011 : OAI22_X1 port map( A1 => n21229, A2 => n15586, B1 => n21575, B2 => 
                           n21221, ZN => n5901);
   U18012 : OAI22_X1 port map( A1 => n21229, A2 => n15585, B1 => n21578, B2 => 
                           n21221, ZN => n5902);
   U18013 : OAI22_X1 port map( A1 => n21229, A2 => n15584, B1 => n21581, B2 => 
                           n21221, ZN => n5903);
   U18014 : OAI22_X1 port map( A1 => n21229, A2 => n15583, B1 => n21584, B2 => 
                           n21221, ZN => n5904);
   U18015 : OAI22_X1 port map( A1 => n21229, A2 => n15582, B1 => n21587, B2 => 
                           n21221, ZN => n5905);
   U18016 : OAI22_X1 port map( A1 => n21229, A2 => n15581, B1 => n21590, B2 => 
                           n21221, ZN => n5906);
   U18017 : OAI22_X1 port map( A1 => n21229, A2 => n15580, B1 => n21593, B2 => 
                           n21221, ZN => n5907);
   U18018 : OAI22_X1 port map( A1 => n21229, A2 => n15579, B1 => n21596, B2 => 
                           n21221, ZN => n5908);
   U18019 : OAI22_X1 port map( A1 => n21229, A2 => n15578, B1 => n21599, B2 => 
                           n21222, ZN => n5909);
   U18020 : OAI22_X1 port map( A1 => n21230, A2 => n15577, B1 => n21602, B2 => 
                           n21222, ZN => n5910);
   U18021 : OAI22_X1 port map( A1 => n21230, A2 => n15576, B1 => n21605, B2 => 
                           n21222, ZN => n5911);
   U18022 : OAI22_X1 port map( A1 => n21230, A2 => n15575, B1 => n21608, B2 => 
                           n21222, ZN => n5912);
   U18023 : OAI22_X1 port map( A1 => n21230, A2 => n15574, B1 => n21611, B2 => 
                           n21222, ZN => n5913);
   U18024 : OAI22_X1 port map( A1 => n21230, A2 => n15573, B1 => n21614, B2 => 
                           n21222, ZN => n5914);
   U18025 : OAI22_X1 port map( A1 => n21230, A2 => n15572, B1 => n21617, B2 => 
                           n21222, ZN => n5915);
   U18026 : OAI22_X1 port map( A1 => n21230, A2 => n15571, B1 => n21620, B2 => 
                           n21222, ZN => n5916);
   U18027 : OAI22_X1 port map( A1 => n21230, A2 => n15570, B1 => n21623, B2 => 
                           n21222, ZN => n5917);
   U18028 : OAI22_X1 port map( A1 => n21230, A2 => n15569, B1 => n21626, B2 => 
                           n21222, ZN => n5918);
   U18029 : OAI22_X1 port map( A1 => n21230, A2 => n15568, B1 => n21629, B2 => 
                           n21222, ZN => n5919);
   U18030 : OAI22_X1 port map( A1 => n21230, A2 => n15567, B1 => n21632, B2 => 
                           n21222, ZN => n5920);
   U18031 : OAI22_X1 port map( A1 => n21230, A2 => n15566, B1 => n21635, B2 => 
                           n21223, ZN => n5921);
   U18032 : OAI22_X1 port map( A1 => n21230, A2 => n15565, B1 => n21638, B2 => 
                           n21223, ZN => n5922);
   U18033 : OAI22_X1 port map( A1 => n21231, A2 => n15564, B1 => n21641, B2 => 
                           n21223, ZN => n5923);
   U18034 : OAI22_X1 port map( A1 => n21231, A2 => n15563, B1 => n21644, B2 => 
                           n21223, ZN => n5924);
   U18035 : OAI22_X1 port map( A1 => n21231, A2 => n15562, B1 => n21647, B2 => 
                           n21223, ZN => n5925);
   U18036 : OAI22_X1 port map( A1 => n21231, A2 => n15561, B1 => n21650, B2 => 
                           n21223, ZN => n5926);
   U18037 : OAI22_X1 port map( A1 => n21231, A2 => n15560, B1 => n21653, B2 => 
                           n21223, ZN => n5927);
   U18038 : OAI22_X1 port map( A1 => n21231, A2 => n15559, B1 => n21656, B2 => 
                           n21223, ZN => n5928);
   U18039 : OAI22_X1 port map( A1 => n21231, A2 => n15558, B1 => n21659, B2 => 
                           n21223, ZN => n5929);
   U18040 : OAI22_X1 port map( A1 => n21231, A2 => n15557, B1 => n21662, B2 => 
                           n21223, ZN => n5930);
   U18041 : OAI22_X1 port map( A1 => n21231, A2 => n15556, B1 => n21665, B2 => 
                           n21223, ZN => n5931);
   U18042 : OAI22_X1 port map( A1 => n21231, A2 => n15555, B1 => n21668, B2 => 
                           n21223, ZN => n5932);
   U18043 : OAI22_X1 port map( A1 => n21231, A2 => n15554, B1 => n21671, B2 => 
                           n21224, ZN => n5933);
   U18044 : OAI22_X1 port map( A1 => n21231, A2 => n15553, B1 => n21674, B2 => 
                           n21224, ZN => n5934);
   U18045 : OAI22_X1 port map( A1 => n21231, A2 => n15552, B1 => n21677, B2 => 
                           n21224, ZN => n5935);
   U18046 : OAI22_X1 port map( A1 => n21232, A2 => n15551, B1 => n21680, B2 => 
                           n21224, ZN => n5936);
   U18047 : OAI22_X1 port map( A1 => n21232, A2 => n15550, B1 => n21683, B2 => 
                           n21224, ZN => n5937);
   U18048 : OAI22_X1 port map( A1 => n21232, A2 => n15549, B1 => n21686, B2 => 
                           n21224, ZN => n5938);
   U18049 : OAI22_X1 port map( A1 => n21232, A2 => n15548, B1 => n21689, B2 => 
                           n21224, ZN => n5939);
   U18050 : OAI22_X1 port map( A1 => n21232, A2 => n15547, B1 => n21692, B2 => 
                           n21224, ZN => n5940);
   U18051 : OAI22_X1 port map( A1 => n21232, A2 => n15546, B1 => n21695, B2 => 
                           n21224, ZN => n5941);
   U18052 : OAI22_X1 port map( A1 => n21232, A2 => n15545, B1 => n21698, B2 => 
                           n21224, ZN => n5942);
   U18053 : OAI22_X1 port map( A1 => n21232, A2 => n15544, B1 => n21701, B2 => 
                           n21224, ZN => n5943);
   U18054 : OAI22_X1 port map( A1 => n21232, A2 => n15543, B1 => n21704, B2 => 
                           n21224, ZN => n5944);
   U18055 : OAI22_X1 port map( A1 => n21241, A2 => n15535, B1 => n21527, B2 => 
                           n21233, ZN => n5949);
   U18056 : OAI22_X1 port map( A1 => n21241, A2 => n15534, B1 => n21530, B2 => 
                           n21233, ZN => n5950);
   U18057 : OAI22_X1 port map( A1 => n21241, A2 => n15533, B1 => n21533, B2 => 
                           n21233, ZN => n5951);
   U18058 : OAI22_X1 port map( A1 => n21241, A2 => n15532, B1 => n21536, B2 => 
                           n21233, ZN => n5952);
   U18059 : OAI22_X1 port map( A1 => n21241, A2 => n15531, B1 => n21539, B2 => 
                           n21233, ZN => n5953);
   U18060 : OAI22_X1 port map( A1 => n21241, A2 => n15530, B1 => n21542, B2 => 
                           n21233, ZN => n5954);
   U18061 : OAI22_X1 port map( A1 => n21241, A2 => n15529, B1 => n21545, B2 => 
                           n21233, ZN => n5955);
   U18062 : OAI22_X1 port map( A1 => n21241, A2 => n15528, B1 => n21548, B2 => 
                           n21233, ZN => n5956);
   U18063 : OAI22_X1 port map( A1 => n21241, A2 => n15527, B1 => n21551, B2 => 
                           n21233, ZN => n5957);
   U18064 : OAI22_X1 port map( A1 => n21241, A2 => n15526, B1 => n21554, B2 => 
                           n21233, ZN => n5958);
   U18065 : OAI22_X1 port map( A1 => n21241, A2 => n15525, B1 => n21557, B2 => 
                           n21233, ZN => n5959);
   U18066 : OAI22_X1 port map( A1 => n21241, A2 => n15524, B1 => n21560, B2 => 
                           n21233, ZN => n5960);
   U18067 : OAI22_X1 port map( A1 => n21242, A2 => n15523, B1 => n21563, B2 => 
                           n21234, ZN => n5961);
   U18068 : OAI22_X1 port map( A1 => n21242, A2 => n15522, B1 => n21566, B2 => 
                           n21234, ZN => n5962);
   U18069 : OAI22_X1 port map( A1 => n21242, A2 => n15521, B1 => n21569, B2 => 
                           n21234, ZN => n5963);
   U18070 : OAI22_X1 port map( A1 => n21242, A2 => n15520, B1 => n21572, B2 => 
                           n21234, ZN => n5964);
   U18071 : OAI22_X1 port map( A1 => n21242, A2 => n15519, B1 => n21575, B2 => 
                           n21234, ZN => n5965);
   U18072 : OAI22_X1 port map( A1 => n21242, A2 => n15518, B1 => n21578, B2 => 
                           n21234, ZN => n5966);
   U18073 : OAI22_X1 port map( A1 => n21242, A2 => n15517, B1 => n21581, B2 => 
                           n21234, ZN => n5967);
   U18074 : OAI22_X1 port map( A1 => n21242, A2 => n15516, B1 => n21584, B2 => 
                           n21234, ZN => n5968);
   U18075 : OAI22_X1 port map( A1 => n21242, A2 => n15515, B1 => n21587, B2 => 
                           n21234, ZN => n5969);
   U18076 : OAI22_X1 port map( A1 => n21242, A2 => n15514, B1 => n21590, B2 => 
                           n21234, ZN => n5970);
   U18077 : OAI22_X1 port map( A1 => n21242, A2 => n15513, B1 => n21593, B2 => 
                           n21234, ZN => n5971);
   U18078 : OAI22_X1 port map( A1 => n21242, A2 => n15512, B1 => n21596, B2 => 
                           n21234, ZN => n5972);
   U18079 : OAI22_X1 port map( A1 => n21242, A2 => n15511, B1 => n21599, B2 => 
                           n21235, ZN => n5973);
   U18080 : OAI22_X1 port map( A1 => n21243, A2 => n15510, B1 => n21602, B2 => 
                           n21235, ZN => n5974);
   U18081 : OAI22_X1 port map( A1 => n21243, A2 => n15509, B1 => n21605, B2 => 
                           n21235, ZN => n5975);
   U18082 : OAI22_X1 port map( A1 => n21243, A2 => n15508, B1 => n21608, B2 => 
                           n21235, ZN => n5976);
   U18083 : OAI22_X1 port map( A1 => n21243, A2 => n15507, B1 => n21611, B2 => 
                           n21235, ZN => n5977);
   U18084 : OAI22_X1 port map( A1 => n21243, A2 => n15506, B1 => n21614, B2 => 
                           n21235, ZN => n5978);
   U18085 : OAI22_X1 port map( A1 => n21243, A2 => n15505, B1 => n21617, B2 => 
                           n21235, ZN => n5979);
   U18086 : OAI22_X1 port map( A1 => n21243, A2 => n15504, B1 => n21620, B2 => 
                           n21235, ZN => n5980);
   U18087 : OAI22_X1 port map( A1 => n21243, A2 => n15503, B1 => n21623, B2 => 
                           n21235, ZN => n5981);
   U18088 : OAI22_X1 port map( A1 => n21243, A2 => n15502, B1 => n21626, B2 => 
                           n21235, ZN => n5982);
   U18089 : OAI22_X1 port map( A1 => n21243, A2 => n15501, B1 => n21629, B2 => 
                           n21235, ZN => n5983);
   U18090 : OAI22_X1 port map( A1 => n21243, A2 => n15500, B1 => n21632, B2 => 
                           n21235, ZN => n5984);
   U18091 : OAI22_X1 port map( A1 => n21243, A2 => n15499, B1 => n21635, B2 => 
                           n21236, ZN => n5985);
   U18092 : OAI22_X1 port map( A1 => n21243, A2 => n15498, B1 => n21638, B2 => 
                           n21236, ZN => n5986);
   U18093 : OAI22_X1 port map( A1 => n21244, A2 => n15497, B1 => n21641, B2 => 
                           n21236, ZN => n5987);
   U18094 : OAI22_X1 port map( A1 => n21244, A2 => n15496, B1 => n21644, B2 => 
                           n21236, ZN => n5988);
   U18095 : OAI22_X1 port map( A1 => n21244, A2 => n15495, B1 => n21647, B2 => 
                           n21236, ZN => n5989);
   U18096 : OAI22_X1 port map( A1 => n21244, A2 => n15494, B1 => n21650, B2 => 
                           n21236, ZN => n5990);
   U18097 : OAI22_X1 port map( A1 => n21244, A2 => n15493, B1 => n21653, B2 => 
                           n21236, ZN => n5991);
   U18098 : OAI22_X1 port map( A1 => n21244, A2 => n15492, B1 => n21656, B2 => 
                           n21236, ZN => n5992);
   U18099 : OAI22_X1 port map( A1 => n21244, A2 => n15491, B1 => n21659, B2 => 
                           n21236, ZN => n5993);
   U18100 : OAI22_X1 port map( A1 => n21244, A2 => n15490, B1 => n21662, B2 => 
                           n21236, ZN => n5994);
   U18101 : OAI22_X1 port map( A1 => n21244, A2 => n15489, B1 => n21665, B2 => 
                           n21236, ZN => n5995);
   U18102 : OAI22_X1 port map( A1 => n21244, A2 => n15488, B1 => n21668, B2 => 
                           n21236, ZN => n5996);
   U18103 : OAI22_X1 port map( A1 => n21244, A2 => n15487, B1 => n21671, B2 => 
                           n21237, ZN => n5997);
   U18104 : OAI22_X1 port map( A1 => n21244, A2 => n15486, B1 => n21674, B2 => 
                           n21237, ZN => n5998);
   U18105 : OAI22_X1 port map( A1 => n21244, A2 => n15485, B1 => n21677, B2 => 
                           n21237, ZN => n5999);
   U18106 : OAI22_X1 port map( A1 => n21245, A2 => n15484, B1 => n21680, B2 => 
                           n21237, ZN => n6000);
   U18107 : OAI22_X1 port map( A1 => n21245, A2 => n15483, B1 => n21683, B2 => 
                           n21237, ZN => n6001);
   U18108 : OAI22_X1 port map( A1 => n21245, A2 => n15482, B1 => n21686, B2 => 
                           n21237, ZN => n6002);
   U18109 : OAI22_X1 port map( A1 => n21245, A2 => n15481, B1 => n21689, B2 => 
                           n21237, ZN => n6003);
   U18110 : OAI22_X1 port map( A1 => n21245, A2 => n15480, B1 => n21692, B2 => 
                           n21237, ZN => n6004);
   U18111 : OAI22_X1 port map( A1 => n21245, A2 => n15479, B1 => n21695, B2 => 
                           n21237, ZN => n6005);
   U18112 : OAI22_X1 port map( A1 => n21245, A2 => n15478, B1 => n21698, B2 => 
                           n21237, ZN => n6006);
   U18113 : OAI22_X1 port map( A1 => n21245, A2 => n15477, B1 => n21701, B2 => 
                           n21237, ZN => n6007);
   U18114 : OAI22_X1 port map( A1 => n21245, A2 => n15476, B1 => n21704, B2 => 
                           n21237, ZN => n6008);
   U18115 : OAI22_X1 port map( A1 => n21267, A2 => n15403, B1 => n21527, B2 => 
                           n21259, ZN => n6077);
   U18116 : OAI22_X1 port map( A1 => n21267, A2 => n15402, B1 => n21530, B2 => 
                           n21259, ZN => n6078);
   U18117 : OAI22_X1 port map( A1 => n21267, A2 => n15401, B1 => n21533, B2 => 
                           n21259, ZN => n6079);
   U18118 : OAI22_X1 port map( A1 => n21267, A2 => n15400, B1 => n21536, B2 => 
                           n21259, ZN => n6080);
   U18119 : OAI22_X1 port map( A1 => n21267, A2 => n15399, B1 => n21539, B2 => 
                           n21259, ZN => n6081);
   U18120 : OAI22_X1 port map( A1 => n21267, A2 => n15398, B1 => n21542, B2 => 
                           n21259, ZN => n6082);
   U18121 : OAI22_X1 port map( A1 => n21267, A2 => n15397, B1 => n21545, B2 => 
                           n21259, ZN => n6083);
   U18122 : OAI22_X1 port map( A1 => n21267, A2 => n15396, B1 => n21548, B2 => 
                           n21259, ZN => n6084);
   U18123 : OAI22_X1 port map( A1 => n21267, A2 => n15395, B1 => n21551, B2 => 
                           n21259, ZN => n6085);
   U18124 : OAI22_X1 port map( A1 => n21267, A2 => n15394, B1 => n21554, B2 => 
                           n21259, ZN => n6086);
   U18125 : OAI22_X1 port map( A1 => n21267, A2 => n15393, B1 => n21557, B2 => 
                           n21259, ZN => n6087);
   U18126 : OAI22_X1 port map( A1 => n21267, A2 => n15392, B1 => n21560, B2 => 
                           n21259, ZN => n6088);
   U18127 : OAI22_X1 port map( A1 => n21268, A2 => n15391, B1 => n21563, B2 => 
                           n21260, ZN => n6089);
   U18128 : OAI22_X1 port map( A1 => n21268, A2 => n15390, B1 => n21566, B2 => 
                           n21260, ZN => n6090);
   U18129 : OAI22_X1 port map( A1 => n21268, A2 => n15389, B1 => n21569, B2 => 
                           n21260, ZN => n6091);
   U18130 : OAI22_X1 port map( A1 => n21268, A2 => n15388, B1 => n21572, B2 => 
                           n21260, ZN => n6092);
   U18131 : OAI22_X1 port map( A1 => n21268, A2 => n15387, B1 => n21575, B2 => 
                           n21260, ZN => n6093);
   U18132 : OAI22_X1 port map( A1 => n21268, A2 => n15386, B1 => n21578, B2 => 
                           n21260, ZN => n6094);
   U18133 : OAI22_X1 port map( A1 => n21268, A2 => n15385, B1 => n21581, B2 => 
                           n21260, ZN => n6095);
   U18134 : OAI22_X1 port map( A1 => n21268, A2 => n15384, B1 => n21584, B2 => 
                           n21260, ZN => n6096);
   U18135 : OAI22_X1 port map( A1 => n21268, A2 => n15383, B1 => n21587, B2 => 
                           n21260, ZN => n6097);
   U18136 : OAI22_X1 port map( A1 => n21268, A2 => n15382, B1 => n21590, B2 => 
                           n21260, ZN => n6098);
   U18137 : OAI22_X1 port map( A1 => n21268, A2 => n15381, B1 => n21593, B2 => 
                           n21260, ZN => n6099);
   U18138 : OAI22_X1 port map( A1 => n21268, A2 => n15380, B1 => n21596, B2 => 
                           n21260, ZN => n6100);
   U18139 : OAI22_X1 port map( A1 => n21268, A2 => n15379, B1 => n21599, B2 => 
                           n21261, ZN => n6101);
   U18140 : OAI22_X1 port map( A1 => n21269, A2 => n15378, B1 => n21602, B2 => 
                           n21261, ZN => n6102);
   U18141 : OAI22_X1 port map( A1 => n21269, A2 => n15377, B1 => n21605, B2 => 
                           n21261, ZN => n6103);
   U18142 : OAI22_X1 port map( A1 => n21269, A2 => n15376, B1 => n21608, B2 => 
                           n21261, ZN => n6104);
   U18143 : OAI22_X1 port map( A1 => n21269, A2 => n15375, B1 => n21611, B2 => 
                           n21261, ZN => n6105);
   U18144 : OAI22_X1 port map( A1 => n21269, A2 => n15374, B1 => n21614, B2 => 
                           n21261, ZN => n6106);
   U18145 : OAI22_X1 port map( A1 => n21269, A2 => n15373, B1 => n21617, B2 => 
                           n21261, ZN => n6107);
   U18146 : OAI22_X1 port map( A1 => n21269, A2 => n15372, B1 => n21620, B2 => 
                           n21261, ZN => n6108);
   U18147 : OAI22_X1 port map( A1 => n21269, A2 => n15371, B1 => n21623, B2 => 
                           n21261, ZN => n6109);
   U18148 : OAI22_X1 port map( A1 => n21269, A2 => n15370, B1 => n21626, B2 => 
                           n21261, ZN => n6110);
   U18149 : OAI22_X1 port map( A1 => n21269, A2 => n15369, B1 => n21629, B2 => 
                           n21261, ZN => n6111);
   U18150 : OAI22_X1 port map( A1 => n21269, A2 => n15368, B1 => n21632, B2 => 
                           n21261, ZN => n6112);
   U18151 : OAI22_X1 port map( A1 => n21269, A2 => n15367, B1 => n21635, B2 => 
                           n21262, ZN => n6113);
   U18152 : OAI22_X1 port map( A1 => n21269, A2 => n15366, B1 => n21638, B2 => 
                           n21262, ZN => n6114);
   U18153 : OAI22_X1 port map( A1 => n21270, A2 => n15365, B1 => n21641, B2 => 
                           n21262, ZN => n6115);
   U18154 : OAI22_X1 port map( A1 => n21270, A2 => n15364, B1 => n21644, B2 => 
                           n21262, ZN => n6116);
   U18155 : OAI22_X1 port map( A1 => n21270, A2 => n15363, B1 => n21647, B2 => 
                           n21262, ZN => n6117);
   U18156 : OAI22_X1 port map( A1 => n21270, A2 => n15362, B1 => n21650, B2 => 
                           n21262, ZN => n6118);
   U18157 : OAI22_X1 port map( A1 => n21270, A2 => n15361, B1 => n21653, B2 => 
                           n21262, ZN => n6119);
   U18158 : OAI22_X1 port map( A1 => n21270, A2 => n15360, B1 => n21656, B2 => 
                           n21262, ZN => n6120);
   U18159 : OAI22_X1 port map( A1 => n21270, A2 => n15359, B1 => n21659, B2 => 
                           n21262, ZN => n6121);
   U18160 : OAI22_X1 port map( A1 => n21270, A2 => n15358, B1 => n21662, B2 => 
                           n21262, ZN => n6122);
   U18161 : OAI22_X1 port map( A1 => n21270, A2 => n15357, B1 => n21665, B2 => 
                           n21262, ZN => n6123);
   U18162 : OAI22_X1 port map( A1 => n21270, A2 => n15356, B1 => n21668, B2 => 
                           n21262, ZN => n6124);
   U18163 : OAI22_X1 port map( A1 => n21270, A2 => n15355, B1 => n21671, B2 => 
                           n21263, ZN => n6125);
   U18164 : OAI22_X1 port map( A1 => n21270, A2 => n15354, B1 => n21674, B2 => 
                           n21263, ZN => n6126);
   U18165 : OAI22_X1 port map( A1 => n21270, A2 => n15353, B1 => n21677, B2 => 
                           n21263, ZN => n6127);
   U18166 : OAI22_X1 port map( A1 => n21271, A2 => n15352, B1 => n21680, B2 => 
                           n21263, ZN => n6128);
   U18167 : OAI22_X1 port map( A1 => n21271, A2 => n15351, B1 => n21683, B2 => 
                           n21263, ZN => n6129);
   U18168 : OAI22_X1 port map( A1 => n21271, A2 => n15350, B1 => n21686, B2 => 
                           n21263, ZN => n6130);
   U18169 : OAI22_X1 port map( A1 => n21271, A2 => n15349, B1 => n21689, B2 => 
                           n21263, ZN => n6131);
   U18170 : OAI22_X1 port map( A1 => n21271, A2 => n15348, B1 => n21692, B2 => 
                           n21263, ZN => n6132);
   U18171 : OAI22_X1 port map( A1 => n21271, A2 => n15347, B1 => n21695, B2 => 
                           n21263, ZN => n6133);
   U18172 : OAI22_X1 port map( A1 => n21271, A2 => n15346, B1 => n21698, B2 => 
                           n21263, ZN => n6134);
   U18173 : OAI22_X1 port map( A1 => n21271, A2 => n15345, B1 => n21701, B2 => 
                           n21263, ZN => n6135);
   U18174 : OAI22_X1 port map( A1 => n21271, A2 => n15344, B1 => n21704, B2 => 
                           n21263, ZN => n6136);
   U18175 : OAI22_X1 port map( A1 => n21293, A2 => n15271, B1 => n21527, B2 => 
                           n21285, ZN => n6205);
   U18176 : OAI22_X1 port map( A1 => n21293, A2 => n15270, B1 => n21530, B2 => 
                           n21285, ZN => n6206);
   U18177 : OAI22_X1 port map( A1 => n21293, A2 => n15269, B1 => n21533, B2 => 
                           n21285, ZN => n6207);
   U18178 : OAI22_X1 port map( A1 => n21293, A2 => n15268, B1 => n21536, B2 => 
                           n21285, ZN => n6208);
   U18179 : OAI22_X1 port map( A1 => n21293, A2 => n15267, B1 => n21539, B2 => 
                           n21285, ZN => n6209);
   U18180 : OAI22_X1 port map( A1 => n21293, A2 => n15266, B1 => n21542, B2 => 
                           n21285, ZN => n6210);
   U18181 : OAI22_X1 port map( A1 => n21293, A2 => n15265, B1 => n21545, B2 => 
                           n21285, ZN => n6211);
   U18182 : OAI22_X1 port map( A1 => n21293, A2 => n15264, B1 => n21548, B2 => 
                           n21285, ZN => n6212);
   U18183 : OAI22_X1 port map( A1 => n21293, A2 => n15263, B1 => n21551, B2 => 
                           n21285, ZN => n6213);
   U18184 : OAI22_X1 port map( A1 => n21293, A2 => n15262, B1 => n21554, B2 => 
                           n21285, ZN => n6214);
   U18185 : OAI22_X1 port map( A1 => n21293, A2 => n15261, B1 => n21557, B2 => 
                           n21285, ZN => n6215);
   U18186 : OAI22_X1 port map( A1 => n21293, A2 => n15260, B1 => n21560, B2 => 
                           n21285, ZN => n6216);
   U18187 : OAI22_X1 port map( A1 => n21294, A2 => n15259, B1 => n21563, B2 => 
                           n21286, ZN => n6217);
   U18188 : OAI22_X1 port map( A1 => n21294, A2 => n15258, B1 => n21566, B2 => 
                           n21286, ZN => n6218);
   U18189 : OAI22_X1 port map( A1 => n21294, A2 => n15257, B1 => n21569, B2 => 
                           n21286, ZN => n6219);
   U18190 : OAI22_X1 port map( A1 => n21294, A2 => n15256, B1 => n21572, B2 => 
                           n21286, ZN => n6220);
   U18191 : OAI22_X1 port map( A1 => n21294, A2 => n15255, B1 => n21575, B2 => 
                           n21286, ZN => n6221);
   U18192 : OAI22_X1 port map( A1 => n21294, A2 => n15254, B1 => n21578, B2 => 
                           n21286, ZN => n6222);
   U18193 : OAI22_X1 port map( A1 => n21294, A2 => n15253, B1 => n21581, B2 => 
                           n21286, ZN => n6223);
   U18194 : OAI22_X1 port map( A1 => n21294, A2 => n15252, B1 => n21584, B2 => 
                           n21286, ZN => n6224);
   U18195 : OAI22_X1 port map( A1 => n21294, A2 => n15251, B1 => n21587, B2 => 
                           n21286, ZN => n6225);
   U18196 : OAI22_X1 port map( A1 => n21294, A2 => n15250, B1 => n21590, B2 => 
                           n21286, ZN => n6226);
   U18197 : OAI22_X1 port map( A1 => n21294, A2 => n15249, B1 => n21593, B2 => 
                           n21286, ZN => n6227);
   U18198 : OAI22_X1 port map( A1 => n21294, A2 => n15248, B1 => n21596, B2 => 
                           n21286, ZN => n6228);
   U18199 : OAI22_X1 port map( A1 => n21294, A2 => n15247, B1 => n21599, B2 => 
                           n21287, ZN => n6229);
   U18200 : OAI22_X1 port map( A1 => n21295, A2 => n15246, B1 => n21602, B2 => 
                           n21287, ZN => n6230);
   U18201 : OAI22_X1 port map( A1 => n21295, A2 => n15245, B1 => n21605, B2 => 
                           n21287, ZN => n6231);
   U18202 : OAI22_X1 port map( A1 => n21295, A2 => n15244, B1 => n21608, B2 => 
                           n21287, ZN => n6232);
   U18203 : OAI22_X1 port map( A1 => n21295, A2 => n15243, B1 => n21611, B2 => 
                           n21287, ZN => n6233);
   U18204 : OAI22_X1 port map( A1 => n21295, A2 => n15242, B1 => n21614, B2 => 
                           n21287, ZN => n6234);
   U18205 : OAI22_X1 port map( A1 => n21295, A2 => n15241, B1 => n21617, B2 => 
                           n21287, ZN => n6235);
   U18206 : OAI22_X1 port map( A1 => n21295, A2 => n15240, B1 => n21620, B2 => 
                           n21287, ZN => n6236);
   U18207 : OAI22_X1 port map( A1 => n21295, A2 => n15239, B1 => n21623, B2 => 
                           n21287, ZN => n6237);
   U18208 : OAI22_X1 port map( A1 => n21295, A2 => n15238, B1 => n21626, B2 => 
                           n21287, ZN => n6238);
   U18209 : OAI22_X1 port map( A1 => n21295, A2 => n15237, B1 => n21629, B2 => 
                           n21287, ZN => n6239);
   U18210 : OAI22_X1 port map( A1 => n21295, A2 => n15236, B1 => n21632, B2 => 
                           n21287, ZN => n6240);
   U18211 : OAI22_X1 port map( A1 => n21295, A2 => n15235, B1 => n21635, B2 => 
                           n21288, ZN => n6241);
   U18212 : OAI22_X1 port map( A1 => n21295, A2 => n15234, B1 => n21638, B2 => 
                           n21288, ZN => n6242);
   U18213 : OAI22_X1 port map( A1 => n21296, A2 => n15233, B1 => n21641, B2 => 
                           n21288, ZN => n6243);
   U18214 : OAI22_X1 port map( A1 => n21296, A2 => n15232, B1 => n21644, B2 => 
                           n21288, ZN => n6244);
   U18215 : OAI22_X1 port map( A1 => n21296, A2 => n15231, B1 => n21647, B2 => 
                           n21288, ZN => n6245);
   U18216 : OAI22_X1 port map( A1 => n21296, A2 => n15230, B1 => n21650, B2 => 
                           n21288, ZN => n6246);
   U18217 : OAI22_X1 port map( A1 => n21296, A2 => n15229, B1 => n21653, B2 => 
                           n21288, ZN => n6247);
   U18218 : OAI22_X1 port map( A1 => n21296, A2 => n15228, B1 => n21656, B2 => 
                           n21288, ZN => n6248);
   U18219 : OAI22_X1 port map( A1 => n21296, A2 => n15227, B1 => n21659, B2 => 
                           n21288, ZN => n6249);
   U18220 : OAI22_X1 port map( A1 => n21296, A2 => n15226, B1 => n21662, B2 => 
                           n21288, ZN => n6250);
   U18221 : OAI22_X1 port map( A1 => n21296, A2 => n15225, B1 => n21665, B2 => 
                           n21288, ZN => n6251);
   U18222 : OAI22_X1 port map( A1 => n21296, A2 => n15224, B1 => n21668, B2 => 
                           n21288, ZN => n6252);
   U18223 : OAI22_X1 port map( A1 => n21296, A2 => n15223, B1 => n21671, B2 => 
                           n21289, ZN => n6253);
   U18224 : OAI22_X1 port map( A1 => n21296, A2 => n15222, B1 => n21674, B2 => 
                           n21289, ZN => n6254);
   U18225 : OAI22_X1 port map( A1 => n21296, A2 => n15221, B1 => n21677, B2 => 
                           n21289, ZN => n6255);
   U18226 : OAI22_X1 port map( A1 => n21297, A2 => n15220, B1 => n21680, B2 => 
                           n21289, ZN => n6256);
   U18227 : OAI22_X1 port map( A1 => n21297, A2 => n15219, B1 => n21683, B2 => 
                           n21289, ZN => n6257);
   U18228 : OAI22_X1 port map( A1 => n21297, A2 => n15218, B1 => n21686, B2 => 
                           n21289, ZN => n6258);
   U18229 : OAI22_X1 port map( A1 => n21297, A2 => n15217, B1 => n21689, B2 => 
                           n21289, ZN => n6259);
   U18230 : OAI22_X1 port map( A1 => n21297, A2 => n15216, B1 => n21692, B2 => 
                           n21289, ZN => n6260);
   U18231 : OAI22_X1 port map( A1 => n21297, A2 => n15215, B1 => n21695, B2 => 
                           n21289, ZN => n6261);
   U18232 : OAI22_X1 port map( A1 => n21297, A2 => n15214, B1 => n21698, B2 => 
                           n21289, ZN => n6262);
   U18233 : OAI22_X1 port map( A1 => n21297, A2 => n15213, B1 => n21701, B2 => 
                           n21289, ZN => n6263);
   U18234 : OAI22_X1 port map( A1 => n21297, A2 => n15212, B1 => n21704, B2 => 
                           n21289, ZN => n6264);
   U18235 : OAI22_X1 port map( A1 => n21306, A2 => n15204, B1 => n21527, B2 => 
                           n21298, ZN => n6269);
   U18236 : OAI22_X1 port map( A1 => n21306, A2 => n15203, B1 => n21530, B2 => 
                           n21298, ZN => n6270);
   U18237 : OAI22_X1 port map( A1 => n21306, A2 => n15202, B1 => n21533, B2 => 
                           n21298, ZN => n6271);
   U18238 : OAI22_X1 port map( A1 => n21306, A2 => n15201, B1 => n21536, B2 => 
                           n21298, ZN => n6272);
   U18239 : OAI22_X1 port map( A1 => n21306, A2 => n15200, B1 => n21539, B2 => 
                           n21298, ZN => n6273);
   U18240 : OAI22_X1 port map( A1 => n21306, A2 => n15199, B1 => n21542, B2 => 
                           n21298, ZN => n6274);
   U18241 : OAI22_X1 port map( A1 => n21306, A2 => n15198, B1 => n21545, B2 => 
                           n21298, ZN => n6275);
   U18242 : OAI22_X1 port map( A1 => n21306, A2 => n15197, B1 => n21548, B2 => 
                           n21298, ZN => n6276);
   U18243 : OAI22_X1 port map( A1 => n21306, A2 => n15196, B1 => n21551, B2 => 
                           n21298, ZN => n6277);
   U18244 : OAI22_X1 port map( A1 => n21306, A2 => n15195, B1 => n21554, B2 => 
                           n21298, ZN => n6278);
   U18245 : OAI22_X1 port map( A1 => n21306, A2 => n15194, B1 => n21557, B2 => 
                           n21298, ZN => n6279);
   U18246 : OAI22_X1 port map( A1 => n21306, A2 => n15193, B1 => n21560, B2 => 
                           n21298, ZN => n6280);
   U18247 : OAI22_X1 port map( A1 => n21307, A2 => n15192, B1 => n21563, B2 => 
                           n21299, ZN => n6281);
   U18248 : OAI22_X1 port map( A1 => n21307, A2 => n15191, B1 => n21566, B2 => 
                           n21299, ZN => n6282);
   U18249 : OAI22_X1 port map( A1 => n21307, A2 => n15190, B1 => n21569, B2 => 
                           n21299, ZN => n6283);
   U18250 : OAI22_X1 port map( A1 => n21307, A2 => n15189, B1 => n21572, B2 => 
                           n21299, ZN => n6284);
   U18251 : OAI22_X1 port map( A1 => n21307, A2 => n15188, B1 => n21575, B2 => 
                           n21299, ZN => n6285);
   U18252 : OAI22_X1 port map( A1 => n21307, A2 => n15187, B1 => n21578, B2 => 
                           n21299, ZN => n6286);
   U18253 : OAI22_X1 port map( A1 => n21307, A2 => n15186, B1 => n21581, B2 => 
                           n21299, ZN => n6287);
   U18254 : OAI22_X1 port map( A1 => n21307, A2 => n15185, B1 => n21584, B2 => 
                           n21299, ZN => n6288);
   U18255 : OAI22_X1 port map( A1 => n21307, A2 => n15184, B1 => n21587, B2 => 
                           n21299, ZN => n6289);
   U18256 : OAI22_X1 port map( A1 => n21307, A2 => n15183, B1 => n21590, B2 => 
                           n21299, ZN => n6290);
   U18257 : OAI22_X1 port map( A1 => n21307, A2 => n15182, B1 => n21593, B2 => 
                           n21299, ZN => n6291);
   U18258 : OAI22_X1 port map( A1 => n21307, A2 => n15181, B1 => n21596, B2 => 
                           n21299, ZN => n6292);
   U18259 : OAI22_X1 port map( A1 => n21307, A2 => n15180, B1 => n21599, B2 => 
                           n21300, ZN => n6293);
   U18260 : OAI22_X1 port map( A1 => n21308, A2 => n15179, B1 => n21602, B2 => 
                           n21300, ZN => n6294);
   U18261 : OAI22_X1 port map( A1 => n21308, A2 => n15178, B1 => n21605, B2 => 
                           n21300, ZN => n6295);
   U18262 : OAI22_X1 port map( A1 => n21308, A2 => n15177, B1 => n21608, B2 => 
                           n21300, ZN => n6296);
   U18263 : OAI22_X1 port map( A1 => n21308, A2 => n15176, B1 => n21611, B2 => 
                           n21300, ZN => n6297);
   U18264 : OAI22_X1 port map( A1 => n21308, A2 => n15175, B1 => n21614, B2 => 
                           n21300, ZN => n6298);
   U18265 : OAI22_X1 port map( A1 => n21308, A2 => n15174, B1 => n21617, B2 => 
                           n21300, ZN => n6299);
   U18266 : OAI22_X1 port map( A1 => n21308, A2 => n15173, B1 => n21620, B2 => 
                           n21300, ZN => n6300);
   U18267 : OAI22_X1 port map( A1 => n21308, A2 => n15172, B1 => n21623, B2 => 
                           n21300, ZN => n6301);
   U18268 : OAI22_X1 port map( A1 => n21308, A2 => n15171, B1 => n21626, B2 => 
                           n21300, ZN => n6302);
   U18269 : OAI22_X1 port map( A1 => n21308, A2 => n15170, B1 => n21629, B2 => 
                           n21300, ZN => n6303);
   U18270 : OAI22_X1 port map( A1 => n21308, A2 => n15169, B1 => n21632, B2 => 
                           n21300, ZN => n6304);
   U18271 : OAI22_X1 port map( A1 => n21308, A2 => n15168, B1 => n21635, B2 => 
                           n21301, ZN => n6305);
   U18272 : OAI22_X1 port map( A1 => n21308, A2 => n15167, B1 => n21638, B2 => 
                           n21301, ZN => n6306);
   U18273 : OAI22_X1 port map( A1 => n21309, A2 => n15166, B1 => n21641, B2 => 
                           n21301, ZN => n6307);
   U18274 : OAI22_X1 port map( A1 => n21309, A2 => n15165, B1 => n21644, B2 => 
                           n21301, ZN => n6308);
   U18275 : OAI22_X1 port map( A1 => n21309, A2 => n15164, B1 => n21647, B2 => 
                           n21301, ZN => n6309);
   U18276 : OAI22_X1 port map( A1 => n21309, A2 => n15163, B1 => n21650, B2 => 
                           n21301, ZN => n6310);
   U18277 : OAI22_X1 port map( A1 => n21309, A2 => n15162, B1 => n21653, B2 => 
                           n21301, ZN => n6311);
   U18278 : OAI22_X1 port map( A1 => n21309, A2 => n15161, B1 => n21656, B2 => 
                           n21301, ZN => n6312);
   U18279 : OAI22_X1 port map( A1 => n21309, A2 => n15160, B1 => n21659, B2 => 
                           n21301, ZN => n6313);
   U18280 : OAI22_X1 port map( A1 => n21309, A2 => n15159, B1 => n21662, B2 => 
                           n21301, ZN => n6314);
   U18281 : OAI22_X1 port map( A1 => n21309, A2 => n15158, B1 => n21665, B2 => 
                           n21301, ZN => n6315);
   U18282 : OAI22_X1 port map( A1 => n21309, A2 => n15157, B1 => n21668, B2 => 
                           n21301, ZN => n6316);
   U18283 : OAI22_X1 port map( A1 => n21309, A2 => n15156, B1 => n21671, B2 => 
                           n21302, ZN => n6317);
   U18284 : OAI22_X1 port map( A1 => n21309, A2 => n15155, B1 => n21674, B2 => 
                           n21302, ZN => n6318);
   U18285 : OAI22_X1 port map( A1 => n21309, A2 => n15154, B1 => n21677, B2 => 
                           n21302, ZN => n6319);
   U18286 : OAI22_X1 port map( A1 => n21310, A2 => n15153, B1 => n21680, B2 => 
                           n21302, ZN => n6320);
   U18287 : OAI22_X1 port map( A1 => n21310, A2 => n15152, B1 => n21683, B2 => 
                           n21302, ZN => n6321);
   U18288 : OAI22_X1 port map( A1 => n21310, A2 => n15151, B1 => n21686, B2 => 
                           n21302, ZN => n6322);
   U18289 : OAI22_X1 port map( A1 => n21310, A2 => n15150, B1 => n21689, B2 => 
                           n21302, ZN => n6323);
   U18290 : OAI22_X1 port map( A1 => n21310, A2 => n15149, B1 => n21692, B2 => 
                           n21302, ZN => n6324);
   U18291 : OAI22_X1 port map( A1 => n21310, A2 => n15148, B1 => n21695, B2 => 
                           n21302, ZN => n6325);
   U18292 : OAI22_X1 port map( A1 => n21310, A2 => n15147, B1 => n21698, B2 => 
                           n21302, ZN => n6326);
   U18293 : OAI22_X1 port map( A1 => n21310, A2 => n15146, B1 => n21701, B2 => 
                           n21302, ZN => n6327);
   U18294 : OAI22_X1 port map( A1 => n21310, A2 => n15145, B1 => n21704, B2 => 
                           n21302, ZN => n6328);
   U18295 : OAI22_X1 port map( A1 => n21319, A2 => n15137, B1 => n21527, B2 => 
                           n21311, ZN => n6333);
   U18296 : OAI22_X1 port map( A1 => n21319, A2 => n15136, B1 => n21530, B2 => 
                           n21311, ZN => n6334);
   U18297 : OAI22_X1 port map( A1 => n21319, A2 => n15135, B1 => n21533, B2 => 
                           n21311, ZN => n6335);
   U18298 : OAI22_X1 port map( A1 => n21319, A2 => n15134, B1 => n21536, B2 => 
                           n21311, ZN => n6336);
   U18299 : OAI22_X1 port map( A1 => n21319, A2 => n15133, B1 => n21539, B2 => 
                           n21311, ZN => n6337);
   U18300 : OAI22_X1 port map( A1 => n21319, A2 => n15132, B1 => n21542, B2 => 
                           n21311, ZN => n6338);
   U18301 : OAI22_X1 port map( A1 => n21319, A2 => n15131, B1 => n21545, B2 => 
                           n21311, ZN => n6339);
   U18302 : OAI22_X1 port map( A1 => n21319, A2 => n15130, B1 => n21548, B2 => 
                           n21311, ZN => n6340);
   U18303 : OAI22_X1 port map( A1 => n21319, A2 => n15129, B1 => n21551, B2 => 
                           n21311, ZN => n6341);
   U18304 : OAI22_X1 port map( A1 => n21319, A2 => n15128, B1 => n21554, B2 => 
                           n21311, ZN => n6342);
   U18305 : OAI22_X1 port map( A1 => n21319, A2 => n15127, B1 => n21557, B2 => 
                           n21311, ZN => n6343);
   U18306 : OAI22_X1 port map( A1 => n21319, A2 => n15126, B1 => n21560, B2 => 
                           n21311, ZN => n6344);
   U18307 : OAI22_X1 port map( A1 => n21320, A2 => n15125, B1 => n21563, B2 => 
                           n21312, ZN => n6345);
   U18308 : OAI22_X1 port map( A1 => n21320, A2 => n15124, B1 => n21566, B2 => 
                           n21312, ZN => n6346);
   U18309 : OAI22_X1 port map( A1 => n21320, A2 => n15123, B1 => n21569, B2 => 
                           n21312, ZN => n6347);
   U18310 : OAI22_X1 port map( A1 => n21320, A2 => n15122, B1 => n21572, B2 => 
                           n21312, ZN => n6348);
   U18311 : OAI22_X1 port map( A1 => n21320, A2 => n15121, B1 => n21575, B2 => 
                           n21312, ZN => n6349);
   U18312 : OAI22_X1 port map( A1 => n21320, A2 => n15120, B1 => n21578, B2 => 
                           n21312, ZN => n6350);
   U18313 : OAI22_X1 port map( A1 => n21320, A2 => n15119, B1 => n21581, B2 => 
                           n21312, ZN => n6351);
   U18314 : OAI22_X1 port map( A1 => n21320, A2 => n15118, B1 => n21584, B2 => 
                           n21312, ZN => n6352);
   U18315 : OAI22_X1 port map( A1 => n21320, A2 => n15117, B1 => n21587, B2 => 
                           n21312, ZN => n6353);
   U18316 : OAI22_X1 port map( A1 => n21320, A2 => n15116, B1 => n21590, B2 => 
                           n21312, ZN => n6354);
   U18317 : OAI22_X1 port map( A1 => n21320, A2 => n15115, B1 => n21593, B2 => 
                           n21312, ZN => n6355);
   U18318 : OAI22_X1 port map( A1 => n21320, A2 => n15114, B1 => n21596, B2 => 
                           n21312, ZN => n6356);
   U18319 : OAI22_X1 port map( A1 => n21320, A2 => n15113, B1 => n21599, B2 => 
                           n21313, ZN => n6357);
   U18320 : OAI22_X1 port map( A1 => n21321, A2 => n15112, B1 => n21602, B2 => 
                           n21313, ZN => n6358);
   U18321 : OAI22_X1 port map( A1 => n21321, A2 => n15111, B1 => n21605, B2 => 
                           n21313, ZN => n6359);
   U18322 : OAI22_X1 port map( A1 => n21321, A2 => n15110, B1 => n21608, B2 => 
                           n21313, ZN => n6360);
   U18323 : OAI22_X1 port map( A1 => n21321, A2 => n15109, B1 => n21611, B2 => 
                           n21313, ZN => n6361);
   U18324 : OAI22_X1 port map( A1 => n21321, A2 => n15108, B1 => n21614, B2 => 
                           n21313, ZN => n6362);
   U18325 : OAI22_X1 port map( A1 => n21321, A2 => n15107, B1 => n21617, B2 => 
                           n21313, ZN => n6363);
   U18326 : OAI22_X1 port map( A1 => n21321, A2 => n15106, B1 => n21620, B2 => 
                           n21313, ZN => n6364);
   U18327 : OAI22_X1 port map( A1 => n21321, A2 => n15105, B1 => n21623, B2 => 
                           n21313, ZN => n6365);
   U18328 : OAI22_X1 port map( A1 => n21321, A2 => n15104, B1 => n21626, B2 => 
                           n21313, ZN => n6366);
   U18329 : OAI22_X1 port map( A1 => n21321, A2 => n15103, B1 => n21629, B2 => 
                           n21313, ZN => n6367);
   U18330 : OAI22_X1 port map( A1 => n21321, A2 => n15102, B1 => n21632, B2 => 
                           n21313, ZN => n6368);
   U18331 : OAI22_X1 port map( A1 => n21321, A2 => n15101, B1 => n21635, B2 => 
                           n21314, ZN => n6369);
   U18332 : OAI22_X1 port map( A1 => n21321, A2 => n15100, B1 => n21638, B2 => 
                           n21314, ZN => n6370);
   U18333 : OAI22_X1 port map( A1 => n21322, A2 => n15099, B1 => n21641, B2 => 
                           n21314, ZN => n6371);
   U18334 : OAI22_X1 port map( A1 => n21322, A2 => n15098, B1 => n21644, B2 => 
                           n21314, ZN => n6372);
   U18335 : OAI22_X1 port map( A1 => n21322, A2 => n15097, B1 => n21647, B2 => 
                           n21314, ZN => n6373);
   U18336 : OAI22_X1 port map( A1 => n21322, A2 => n15096, B1 => n21650, B2 => 
                           n21314, ZN => n6374);
   U18337 : OAI22_X1 port map( A1 => n21322, A2 => n15095, B1 => n21653, B2 => 
                           n21314, ZN => n6375);
   U18338 : OAI22_X1 port map( A1 => n21322, A2 => n15094, B1 => n21656, B2 => 
                           n21314, ZN => n6376);
   U18339 : OAI22_X1 port map( A1 => n21322, A2 => n15093, B1 => n21659, B2 => 
                           n21314, ZN => n6377);
   U18340 : OAI22_X1 port map( A1 => n21322, A2 => n15092, B1 => n21662, B2 => 
                           n21314, ZN => n6378);
   U18341 : OAI22_X1 port map( A1 => n21322, A2 => n15091, B1 => n21665, B2 => 
                           n21314, ZN => n6379);
   U18342 : OAI22_X1 port map( A1 => n21322, A2 => n15090, B1 => n21668, B2 => 
                           n21314, ZN => n6380);
   U18343 : OAI22_X1 port map( A1 => n21322, A2 => n15089, B1 => n21671, B2 => 
                           n21315, ZN => n6381);
   U18344 : OAI22_X1 port map( A1 => n21322, A2 => n15088, B1 => n21674, B2 => 
                           n21315, ZN => n6382);
   U18345 : OAI22_X1 port map( A1 => n21322, A2 => n15087, B1 => n21677, B2 => 
                           n21315, ZN => n6383);
   U18346 : OAI22_X1 port map( A1 => n21323, A2 => n15086, B1 => n21680, B2 => 
                           n21315, ZN => n6384);
   U18347 : OAI22_X1 port map( A1 => n21323, A2 => n15085, B1 => n21683, B2 => 
                           n21315, ZN => n6385);
   U18348 : OAI22_X1 port map( A1 => n21323, A2 => n15084, B1 => n21686, B2 => 
                           n21315, ZN => n6386);
   U18349 : OAI22_X1 port map( A1 => n21323, A2 => n15083, B1 => n21689, B2 => 
                           n21315, ZN => n6387);
   U18350 : OAI22_X1 port map( A1 => n21323, A2 => n15082, B1 => n21692, B2 => 
                           n21315, ZN => n6388);
   U18351 : OAI22_X1 port map( A1 => n21323, A2 => n15081, B1 => n21695, B2 => 
                           n21315, ZN => n6389);
   U18352 : OAI22_X1 port map( A1 => n21323, A2 => n15080, B1 => n21698, B2 => 
                           n21315, ZN => n6390);
   U18353 : OAI22_X1 port map( A1 => n21323, A2 => n15079, B1 => n21701, B2 => 
                           n21315, ZN => n6391);
   U18354 : OAI22_X1 port map( A1 => n21323, A2 => n15078, B1 => n21704, B2 => 
                           n21315, ZN => n6392);
   U18355 : OAI22_X1 port map( A1 => n21397, A2 => n14740, B1 => n21526, B2 => 
                           n21389, ZN => n6717);
   U18356 : OAI22_X1 port map( A1 => n21397, A2 => n14739, B1 => n21529, B2 => 
                           n21389, ZN => n6718);
   U18357 : OAI22_X1 port map( A1 => n21397, A2 => n14738, B1 => n21532, B2 => 
                           n21389, ZN => n6719);
   U18358 : OAI22_X1 port map( A1 => n21397, A2 => n14737, B1 => n21535, B2 => 
                           n21389, ZN => n6720);
   U18359 : OAI22_X1 port map( A1 => n21397, A2 => n14736, B1 => n21538, B2 => 
                           n21389, ZN => n6721);
   U18360 : OAI22_X1 port map( A1 => n21397, A2 => n14735, B1 => n21541, B2 => 
                           n21389, ZN => n6722);
   U18361 : OAI22_X1 port map( A1 => n21397, A2 => n14734, B1 => n21544, B2 => 
                           n21389, ZN => n6723);
   U18362 : OAI22_X1 port map( A1 => n21397, A2 => n14733, B1 => n21547, B2 => 
                           n21389, ZN => n6724);
   U18363 : OAI22_X1 port map( A1 => n21397, A2 => n14732, B1 => n21550, B2 => 
                           n21389, ZN => n6725);
   U18364 : OAI22_X1 port map( A1 => n21397, A2 => n14731, B1 => n21553, B2 => 
                           n21389, ZN => n6726);
   U18365 : OAI22_X1 port map( A1 => n21397, A2 => n14730, B1 => n21556, B2 => 
                           n21389, ZN => n6727);
   U18366 : OAI22_X1 port map( A1 => n21397, A2 => n14729, B1 => n21559, B2 => 
                           n21389, ZN => n6728);
   U18367 : OAI22_X1 port map( A1 => n21398, A2 => n14728, B1 => n21562, B2 => 
                           n21390, ZN => n6729);
   U18368 : OAI22_X1 port map( A1 => n21398, A2 => n14727, B1 => n21565, B2 => 
                           n21390, ZN => n6730);
   U18369 : OAI22_X1 port map( A1 => n21398, A2 => n14726, B1 => n21568, B2 => 
                           n21390, ZN => n6731);
   U18370 : OAI22_X1 port map( A1 => n21398, A2 => n14725, B1 => n21571, B2 => 
                           n21390, ZN => n6732);
   U18371 : OAI22_X1 port map( A1 => n21398, A2 => n14724, B1 => n21574, B2 => 
                           n21390, ZN => n6733);
   U18372 : OAI22_X1 port map( A1 => n21398, A2 => n14723, B1 => n21577, B2 => 
                           n21390, ZN => n6734);
   U18373 : OAI22_X1 port map( A1 => n21398, A2 => n14722, B1 => n21580, B2 => 
                           n21390, ZN => n6735);
   U18374 : OAI22_X1 port map( A1 => n21398, A2 => n14721, B1 => n21583, B2 => 
                           n21390, ZN => n6736);
   U18375 : OAI22_X1 port map( A1 => n21398, A2 => n14720, B1 => n21586, B2 => 
                           n21390, ZN => n6737);
   U18376 : OAI22_X1 port map( A1 => n21398, A2 => n14719, B1 => n21589, B2 => 
                           n21390, ZN => n6738);
   U18377 : OAI22_X1 port map( A1 => n21398, A2 => n14718, B1 => n21592, B2 => 
                           n21390, ZN => n6739);
   U18378 : OAI22_X1 port map( A1 => n21398, A2 => n14717, B1 => n21595, B2 => 
                           n21390, ZN => n6740);
   U18379 : OAI22_X1 port map( A1 => n21398, A2 => n14716, B1 => n21598, B2 => 
                           n21391, ZN => n6741);
   U18380 : OAI22_X1 port map( A1 => n21399, A2 => n14715, B1 => n21601, B2 => 
                           n21391, ZN => n6742);
   U18381 : OAI22_X1 port map( A1 => n21399, A2 => n14714, B1 => n21604, B2 => 
                           n21391, ZN => n6743);
   U18382 : OAI22_X1 port map( A1 => n21399, A2 => n14713, B1 => n21607, B2 => 
                           n21391, ZN => n6744);
   U18383 : OAI22_X1 port map( A1 => n21399, A2 => n14712, B1 => n21610, B2 => 
                           n21391, ZN => n6745);
   U18384 : OAI22_X1 port map( A1 => n21399, A2 => n14711, B1 => n21613, B2 => 
                           n21391, ZN => n6746);
   U18385 : OAI22_X1 port map( A1 => n21399, A2 => n14710, B1 => n21616, B2 => 
                           n21391, ZN => n6747);
   U18386 : OAI22_X1 port map( A1 => n21399, A2 => n14709, B1 => n21619, B2 => 
                           n21391, ZN => n6748);
   U18387 : OAI22_X1 port map( A1 => n21399, A2 => n14708, B1 => n21622, B2 => 
                           n21391, ZN => n6749);
   U18388 : OAI22_X1 port map( A1 => n21399, A2 => n14707, B1 => n21625, B2 => 
                           n21391, ZN => n6750);
   U18389 : OAI22_X1 port map( A1 => n21399, A2 => n14706, B1 => n21628, B2 => 
                           n21391, ZN => n6751);
   U18390 : OAI22_X1 port map( A1 => n21399, A2 => n14705, B1 => n21631, B2 => 
                           n21391, ZN => n6752);
   U18391 : OAI22_X1 port map( A1 => n21399, A2 => n14704, B1 => n21634, B2 => 
                           n21392, ZN => n6753);
   U18392 : OAI22_X1 port map( A1 => n21399, A2 => n14703, B1 => n21637, B2 => 
                           n21392, ZN => n6754);
   U18393 : OAI22_X1 port map( A1 => n21400, A2 => n14702, B1 => n21640, B2 => 
                           n21392, ZN => n6755);
   U18394 : OAI22_X1 port map( A1 => n21400, A2 => n14701, B1 => n21643, B2 => 
                           n21392, ZN => n6756);
   U18395 : OAI22_X1 port map( A1 => n21400, A2 => n14700, B1 => n21646, B2 => 
                           n21392, ZN => n6757);
   U18396 : OAI22_X1 port map( A1 => n21400, A2 => n14699, B1 => n21649, B2 => 
                           n21392, ZN => n6758);
   U18397 : OAI22_X1 port map( A1 => n21400, A2 => n14698, B1 => n21652, B2 => 
                           n21392, ZN => n6759);
   U18398 : OAI22_X1 port map( A1 => n21400, A2 => n14697, B1 => n21655, B2 => 
                           n21392, ZN => n6760);
   U18399 : OAI22_X1 port map( A1 => n21400, A2 => n14696, B1 => n21658, B2 => 
                           n21392, ZN => n6761);
   U18400 : OAI22_X1 port map( A1 => n21400, A2 => n14695, B1 => n21661, B2 => 
                           n21392, ZN => n6762);
   U18401 : OAI22_X1 port map( A1 => n21400, A2 => n14694, B1 => n21664, B2 => 
                           n21392, ZN => n6763);
   U18402 : OAI22_X1 port map( A1 => n21400, A2 => n14693, B1 => n21667, B2 => 
                           n21392, ZN => n6764);
   U18403 : OAI22_X1 port map( A1 => n21400, A2 => n14692, B1 => n21670, B2 => 
                           n21393, ZN => n6765);
   U18404 : OAI22_X1 port map( A1 => n21400, A2 => n14691, B1 => n21673, B2 => 
                           n21393, ZN => n6766);
   U18405 : OAI22_X1 port map( A1 => n21400, A2 => n14690, B1 => n21676, B2 => 
                           n21393, ZN => n6767);
   U18406 : OAI22_X1 port map( A1 => n21401, A2 => n14689, B1 => n21679, B2 => 
                           n21393, ZN => n6768);
   U18407 : OAI22_X1 port map( A1 => n21401, A2 => n14688, B1 => n21682, B2 => 
                           n21393, ZN => n6769);
   U18408 : OAI22_X1 port map( A1 => n21401, A2 => n14687, B1 => n21685, B2 => 
                           n21393, ZN => n6770);
   U18409 : OAI22_X1 port map( A1 => n21401, A2 => n14686, B1 => n21688, B2 => 
                           n21393, ZN => n6771);
   U18410 : OAI22_X1 port map( A1 => n21401, A2 => n14685, B1 => n21691, B2 => 
                           n21393, ZN => n6772);
   U18411 : OAI22_X1 port map( A1 => n21401, A2 => n14684, B1 => n21694, B2 => 
                           n21393, ZN => n6773);
   U18412 : OAI22_X1 port map( A1 => n21401, A2 => n14683, B1 => n21697, B2 => 
                           n21393, ZN => n6774);
   U18413 : OAI22_X1 port map( A1 => n21401, A2 => n14682, B1 => n21700, B2 => 
                           n21393, ZN => n6775);
   U18414 : OAI22_X1 port map( A1 => n21401, A2 => n14681, B1 => n21703, B2 => 
                           n21393, ZN => n6776);
   U18415 : OAI22_X1 port map( A1 => n21410, A2 => n14673, B1 => n21526, B2 => 
                           n21402, ZN => n6781);
   U18416 : OAI22_X1 port map( A1 => n21410, A2 => n14672, B1 => n21529, B2 => 
                           n21402, ZN => n6782);
   U18417 : OAI22_X1 port map( A1 => n21410, A2 => n14671, B1 => n21532, B2 => 
                           n21402, ZN => n6783);
   U18418 : OAI22_X1 port map( A1 => n21410, A2 => n14670, B1 => n21535, B2 => 
                           n21402, ZN => n6784);
   U18419 : OAI22_X1 port map( A1 => n21410, A2 => n14669, B1 => n21538, B2 => 
                           n21402, ZN => n6785);
   U18420 : OAI22_X1 port map( A1 => n21410, A2 => n14668, B1 => n21541, B2 => 
                           n21402, ZN => n6786);
   U18421 : OAI22_X1 port map( A1 => n21410, A2 => n14667, B1 => n21544, B2 => 
                           n21402, ZN => n6787);
   U18422 : OAI22_X1 port map( A1 => n21410, A2 => n14666, B1 => n21547, B2 => 
                           n21402, ZN => n6788);
   U18423 : OAI22_X1 port map( A1 => n21410, A2 => n14665, B1 => n21550, B2 => 
                           n21402, ZN => n6789);
   U18424 : OAI22_X1 port map( A1 => n21410, A2 => n14664, B1 => n21553, B2 => 
                           n21402, ZN => n6790);
   U18425 : OAI22_X1 port map( A1 => n21410, A2 => n14663, B1 => n21556, B2 => 
                           n21402, ZN => n6791);
   U18426 : OAI22_X1 port map( A1 => n21410, A2 => n14662, B1 => n21559, B2 => 
                           n21402, ZN => n6792);
   U18427 : OAI22_X1 port map( A1 => n21411, A2 => n14661, B1 => n21562, B2 => 
                           n21403, ZN => n6793);
   U18428 : OAI22_X1 port map( A1 => n21411, A2 => n14660, B1 => n21565, B2 => 
                           n21403, ZN => n6794);
   U18429 : OAI22_X1 port map( A1 => n21411, A2 => n14659, B1 => n21568, B2 => 
                           n21403, ZN => n6795);
   U18430 : OAI22_X1 port map( A1 => n21411, A2 => n14658, B1 => n21571, B2 => 
                           n21403, ZN => n6796);
   U18431 : OAI22_X1 port map( A1 => n21411, A2 => n14657, B1 => n21574, B2 => 
                           n21403, ZN => n6797);
   U18432 : OAI22_X1 port map( A1 => n21411, A2 => n14656, B1 => n21577, B2 => 
                           n21403, ZN => n6798);
   U18433 : OAI22_X1 port map( A1 => n21411, A2 => n14655, B1 => n21580, B2 => 
                           n21403, ZN => n6799);
   U18434 : OAI22_X1 port map( A1 => n21411, A2 => n14654, B1 => n21583, B2 => 
                           n21403, ZN => n6800);
   U18435 : OAI22_X1 port map( A1 => n21411, A2 => n14653, B1 => n21586, B2 => 
                           n21403, ZN => n6801);
   U18436 : OAI22_X1 port map( A1 => n21411, A2 => n14652, B1 => n21589, B2 => 
                           n21403, ZN => n6802);
   U18437 : OAI22_X1 port map( A1 => n21411, A2 => n14651, B1 => n21592, B2 => 
                           n21403, ZN => n6803);
   U18438 : OAI22_X1 port map( A1 => n21411, A2 => n14650, B1 => n21595, B2 => 
                           n21403, ZN => n6804);
   U18439 : OAI22_X1 port map( A1 => n21411, A2 => n14649, B1 => n21598, B2 => 
                           n21404, ZN => n6805);
   U18440 : OAI22_X1 port map( A1 => n21412, A2 => n14648, B1 => n21601, B2 => 
                           n21404, ZN => n6806);
   U18441 : OAI22_X1 port map( A1 => n21412, A2 => n14647, B1 => n21604, B2 => 
                           n21404, ZN => n6807);
   U18442 : OAI22_X1 port map( A1 => n21412, A2 => n14646, B1 => n21607, B2 => 
                           n21404, ZN => n6808);
   U18443 : OAI22_X1 port map( A1 => n21412, A2 => n14645, B1 => n21610, B2 => 
                           n21404, ZN => n6809);
   U18444 : OAI22_X1 port map( A1 => n21412, A2 => n14644, B1 => n21613, B2 => 
                           n21404, ZN => n6810);
   U18445 : OAI22_X1 port map( A1 => n21412, A2 => n14643, B1 => n21616, B2 => 
                           n21404, ZN => n6811);
   U18446 : OAI22_X1 port map( A1 => n21412, A2 => n14642, B1 => n21619, B2 => 
                           n21404, ZN => n6812);
   U18447 : OAI22_X1 port map( A1 => n21412, A2 => n14641, B1 => n21622, B2 => 
                           n21404, ZN => n6813);
   U18448 : OAI22_X1 port map( A1 => n21412, A2 => n14640, B1 => n21625, B2 => 
                           n21404, ZN => n6814);
   U18449 : OAI22_X1 port map( A1 => n21412, A2 => n14639, B1 => n21628, B2 => 
                           n21404, ZN => n6815);
   U18450 : OAI22_X1 port map( A1 => n21412, A2 => n14638, B1 => n21631, B2 => 
                           n21404, ZN => n6816);
   U18451 : OAI22_X1 port map( A1 => n21412, A2 => n14637, B1 => n21634, B2 => 
                           n21405, ZN => n6817);
   U18452 : OAI22_X1 port map( A1 => n21412, A2 => n14636, B1 => n21637, B2 => 
                           n21405, ZN => n6818);
   U18453 : OAI22_X1 port map( A1 => n21413, A2 => n14635, B1 => n21640, B2 => 
                           n21405, ZN => n6819);
   U18454 : OAI22_X1 port map( A1 => n21413, A2 => n14634, B1 => n21643, B2 => 
                           n21405, ZN => n6820);
   U18455 : OAI22_X1 port map( A1 => n21413, A2 => n14633, B1 => n21646, B2 => 
                           n21405, ZN => n6821);
   U18456 : OAI22_X1 port map( A1 => n21413, A2 => n14632, B1 => n21649, B2 => 
                           n21405, ZN => n6822);
   U18457 : OAI22_X1 port map( A1 => n21413, A2 => n14631, B1 => n21652, B2 => 
                           n21405, ZN => n6823);
   U18458 : OAI22_X1 port map( A1 => n21413, A2 => n14630, B1 => n21655, B2 => 
                           n21405, ZN => n6824);
   U18459 : OAI22_X1 port map( A1 => n21413, A2 => n14629, B1 => n21658, B2 => 
                           n21405, ZN => n6825);
   U18460 : OAI22_X1 port map( A1 => n21413, A2 => n14628, B1 => n21661, B2 => 
                           n21405, ZN => n6826);
   U18461 : OAI22_X1 port map( A1 => n21413, A2 => n14627, B1 => n21664, B2 => 
                           n21405, ZN => n6827);
   U18462 : OAI22_X1 port map( A1 => n21413, A2 => n14626, B1 => n21667, B2 => 
                           n21405, ZN => n6828);
   U18463 : OAI22_X1 port map( A1 => n21413, A2 => n14625, B1 => n21670, B2 => 
                           n21406, ZN => n6829);
   U18464 : OAI22_X1 port map( A1 => n21413, A2 => n14624, B1 => n21673, B2 => 
                           n21406, ZN => n6830);
   U18465 : OAI22_X1 port map( A1 => n21413, A2 => n14623, B1 => n21676, B2 => 
                           n21406, ZN => n6831);
   U18466 : OAI22_X1 port map( A1 => n21414, A2 => n14622, B1 => n21679, B2 => 
                           n21406, ZN => n6832);
   U18467 : OAI22_X1 port map( A1 => n21414, A2 => n14621, B1 => n21682, B2 => 
                           n21406, ZN => n6833);
   U18468 : OAI22_X1 port map( A1 => n21414, A2 => n14620, B1 => n21685, B2 => 
                           n21406, ZN => n6834);
   U18469 : OAI22_X1 port map( A1 => n21414, A2 => n14619, B1 => n21688, B2 => 
                           n21406, ZN => n6835);
   U18470 : OAI22_X1 port map( A1 => n21414, A2 => n14618, B1 => n21691, B2 => 
                           n21406, ZN => n6836);
   U18471 : OAI22_X1 port map( A1 => n21414, A2 => n14617, B1 => n21694, B2 => 
                           n21406, ZN => n6837);
   U18472 : OAI22_X1 port map( A1 => n21414, A2 => n14616, B1 => n21697, B2 => 
                           n21406, ZN => n6838);
   U18473 : OAI22_X1 port map( A1 => n21414, A2 => n14615, B1 => n21700, B2 => 
                           n21406, ZN => n6839);
   U18474 : OAI22_X1 port map( A1 => n21414, A2 => n14614, B1 => n21703, B2 => 
                           n21406, ZN => n6840);
   U18475 : OAI22_X1 port map( A1 => n21449, A2 => n14470, B1 => n21526, B2 => 
                           n21441, ZN => n6973);
   U18476 : OAI22_X1 port map( A1 => n21449, A2 => n14469, B1 => n21529, B2 => 
                           n21441, ZN => n6974);
   U18477 : OAI22_X1 port map( A1 => n21449, A2 => n14468, B1 => n21532, B2 => 
                           n21441, ZN => n6975);
   U18478 : OAI22_X1 port map( A1 => n21449, A2 => n14467, B1 => n21535, B2 => 
                           n21441, ZN => n6976);
   U18479 : OAI22_X1 port map( A1 => n21449, A2 => n14466, B1 => n21538, B2 => 
                           n21441, ZN => n6977);
   U18480 : OAI22_X1 port map( A1 => n21449, A2 => n14465, B1 => n21541, B2 => 
                           n21441, ZN => n6978);
   U18481 : OAI22_X1 port map( A1 => n21449, A2 => n14464, B1 => n21544, B2 => 
                           n21441, ZN => n6979);
   U18482 : OAI22_X1 port map( A1 => n21449, A2 => n14463, B1 => n21547, B2 => 
                           n21441, ZN => n6980);
   U18483 : OAI22_X1 port map( A1 => n21449, A2 => n14462, B1 => n21550, B2 => 
                           n21441, ZN => n6981);
   U18484 : OAI22_X1 port map( A1 => n21449, A2 => n14461, B1 => n21553, B2 => 
                           n21441, ZN => n6982);
   U18485 : OAI22_X1 port map( A1 => n21449, A2 => n14460, B1 => n21556, B2 => 
                           n21441, ZN => n6983);
   U18486 : OAI22_X1 port map( A1 => n21449, A2 => n14459, B1 => n21559, B2 => 
                           n21441, ZN => n6984);
   U18487 : OAI22_X1 port map( A1 => n21450, A2 => n14458, B1 => n21562, B2 => 
                           n21442, ZN => n6985);
   U18488 : OAI22_X1 port map( A1 => n21450, A2 => n14457, B1 => n21565, B2 => 
                           n21442, ZN => n6986);
   U18489 : OAI22_X1 port map( A1 => n21450, A2 => n14456, B1 => n21568, B2 => 
                           n21442, ZN => n6987);
   U18490 : OAI22_X1 port map( A1 => n21450, A2 => n14455, B1 => n21571, B2 => 
                           n21442, ZN => n6988);
   U18491 : OAI22_X1 port map( A1 => n21450, A2 => n14454, B1 => n21574, B2 => 
                           n21442, ZN => n6989);
   U18492 : OAI22_X1 port map( A1 => n21450, A2 => n14453, B1 => n21577, B2 => 
                           n21442, ZN => n6990);
   U18493 : OAI22_X1 port map( A1 => n21450, A2 => n14452, B1 => n21580, B2 => 
                           n21442, ZN => n6991);
   U18494 : OAI22_X1 port map( A1 => n21450, A2 => n14451, B1 => n21583, B2 => 
                           n21442, ZN => n6992);
   U18495 : OAI22_X1 port map( A1 => n21450, A2 => n14450, B1 => n21586, B2 => 
                           n21442, ZN => n6993);
   U18496 : OAI22_X1 port map( A1 => n21450, A2 => n14449, B1 => n21589, B2 => 
                           n21442, ZN => n6994);
   U18497 : OAI22_X1 port map( A1 => n21450, A2 => n14448, B1 => n21592, B2 => 
                           n21442, ZN => n6995);
   U18498 : OAI22_X1 port map( A1 => n21450, A2 => n14447, B1 => n21595, B2 => 
                           n21442, ZN => n6996);
   U18499 : OAI22_X1 port map( A1 => n21450, A2 => n14446, B1 => n21598, B2 => 
                           n21443, ZN => n6997);
   U18500 : OAI22_X1 port map( A1 => n21451, A2 => n14445, B1 => n21601, B2 => 
                           n21443, ZN => n6998);
   U18501 : OAI22_X1 port map( A1 => n21451, A2 => n14444, B1 => n21604, B2 => 
                           n21443, ZN => n6999);
   U18502 : OAI22_X1 port map( A1 => n21451, A2 => n14443, B1 => n21607, B2 => 
                           n21443, ZN => n7000);
   U18503 : OAI22_X1 port map( A1 => n21451, A2 => n14442, B1 => n21610, B2 => 
                           n21443, ZN => n7001);
   U18504 : OAI22_X1 port map( A1 => n21451, A2 => n14441, B1 => n21613, B2 => 
                           n21443, ZN => n7002);
   U18505 : OAI22_X1 port map( A1 => n21451, A2 => n14440, B1 => n21616, B2 => 
                           n21443, ZN => n7003);
   U18506 : OAI22_X1 port map( A1 => n21451, A2 => n14439, B1 => n21619, B2 => 
                           n21443, ZN => n7004);
   U18507 : OAI22_X1 port map( A1 => n21451, A2 => n14438, B1 => n21622, B2 => 
                           n21443, ZN => n7005);
   U18508 : OAI22_X1 port map( A1 => n21451, A2 => n14437, B1 => n21625, B2 => 
                           n21443, ZN => n7006);
   U18509 : OAI22_X1 port map( A1 => n21451, A2 => n14436, B1 => n21628, B2 => 
                           n21443, ZN => n7007);
   U18510 : OAI22_X1 port map( A1 => n21451, A2 => n14435, B1 => n21631, B2 => 
                           n21443, ZN => n7008);
   U18511 : OAI22_X1 port map( A1 => n21451, A2 => n14434, B1 => n21634, B2 => 
                           n21444, ZN => n7009);
   U18512 : OAI22_X1 port map( A1 => n21451, A2 => n14433, B1 => n21637, B2 => 
                           n21444, ZN => n7010);
   U18513 : OAI22_X1 port map( A1 => n21452, A2 => n14432, B1 => n21640, B2 => 
                           n21444, ZN => n7011);
   U18514 : OAI22_X1 port map( A1 => n21452, A2 => n14431, B1 => n21643, B2 => 
                           n21444, ZN => n7012);
   U18515 : OAI22_X1 port map( A1 => n21452, A2 => n14430, B1 => n21646, B2 => 
                           n21444, ZN => n7013);
   U18516 : OAI22_X1 port map( A1 => n21452, A2 => n14429, B1 => n21649, B2 => 
                           n21444, ZN => n7014);
   U18517 : OAI22_X1 port map( A1 => n21452, A2 => n14428, B1 => n21652, B2 => 
                           n21444, ZN => n7015);
   U18518 : OAI22_X1 port map( A1 => n21452, A2 => n14427, B1 => n21655, B2 => 
                           n21444, ZN => n7016);
   U18519 : OAI22_X1 port map( A1 => n21452, A2 => n14426, B1 => n21658, B2 => 
                           n21444, ZN => n7017);
   U18520 : OAI22_X1 port map( A1 => n21452, A2 => n14425, B1 => n21661, B2 => 
                           n21444, ZN => n7018);
   U18521 : OAI22_X1 port map( A1 => n21452, A2 => n14424, B1 => n21664, B2 => 
                           n21444, ZN => n7019);
   U18522 : OAI22_X1 port map( A1 => n21452, A2 => n14423, B1 => n21667, B2 => 
                           n21444, ZN => n7020);
   U18523 : OAI22_X1 port map( A1 => n21452, A2 => n14422, B1 => n21670, B2 => 
                           n21445, ZN => n7021);
   U18524 : OAI22_X1 port map( A1 => n21452, A2 => n14421, B1 => n21673, B2 => 
                           n21445, ZN => n7022);
   U18525 : OAI22_X1 port map( A1 => n21452, A2 => n14420, B1 => n21676, B2 => 
                           n21445, ZN => n7023);
   U18526 : OAI22_X1 port map( A1 => n21453, A2 => n14419, B1 => n21679, B2 => 
                           n21445, ZN => n7024);
   U18527 : OAI22_X1 port map( A1 => n21453, A2 => n14418, B1 => n21682, B2 => 
                           n21445, ZN => n7025);
   U18528 : OAI22_X1 port map( A1 => n21453, A2 => n14417, B1 => n21685, B2 => 
                           n21445, ZN => n7026);
   U18529 : OAI22_X1 port map( A1 => n21453, A2 => n14416, B1 => n21688, B2 => 
                           n21445, ZN => n7027);
   U18530 : OAI22_X1 port map( A1 => n21453, A2 => n14415, B1 => n21691, B2 => 
                           n21445, ZN => n7028);
   U18531 : OAI22_X1 port map( A1 => n21453, A2 => n14414, B1 => n21694, B2 => 
                           n21445, ZN => n7029);
   U18532 : OAI22_X1 port map( A1 => n21453, A2 => n14413, B1 => n21697, B2 => 
                           n21445, ZN => n7030);
   U18533 : OAI22_X1 port map( A1 => n21453, A2 => n14412, B1 => n21700, B2 => 
                           n21445, ZN => n7031);
   U18534 : OAI22_X1 port map( A1 => n21453, A2 => n14411, B1 => n21703, B2 => 
                           n21445, ZN => n7032);
   U18535 : OAI22_X1 port map( A1 => n21501, A2 => n14204, B1 => n21526, B2 => 
                           n21493, ZN => n7229);
   U18536 : OAI22_X1 port map( A1 => n21501, A2 => n14203, B1 => n21529, B2 => 
                           n21493, ZN => n7230);
   U18537 : OAI22_X1 port map( A1 => n21501, A2 => n14202, B1 => n21532, B2 => 
                           n21493, ZN => n7231);
   U18538 : OAI22_X1 port map( A1 => n21501, A2 => n14201, B1 => n21535, B2 => 
                           n21493, ZN => n7232);
   U18539 : OAI22_X1 port map( A1 => n21501, A2 => n14200, B1 => n21538, B2 => 
                           n21493, ZN => n7233);
   U18540 : OAI22_X1 port map( A1 => n21501, A2 => n14199, B1 => n21541, B2 => 
                           n21493, ZN => n7234);
   U18541 : OAI22_X1 port map( A1 => n21501, A2 => n14198, B1 => n21544, B2 => 
                           n21493, ZN => n7235);
   U18542 : OAI22_X1 port map( A1 => n21501, A2 => n14197, B1 => n21547, B2 => 
                           n21493, ZN => n7236);
   U18543 : OAI22_X1 port map( A1 => n21501, A2 => n14196, B1 => n21550, B2 => 
                           n21493, ZN => n7237);
   U18544 : OAI22_X1 port map( A1 => n21501, A2 => n14195, B1 => n21553, B2 => 
                           n21493, ZN => n7238);
   U18545 : OAI22_X1 port map( A1 => n21501, A2 => n14194, B1 => n21556, B2 => 
                           n21493, ZN => n7239);
   U18546 : OAI22_X1 port map( A1 => n21501, A2 => n14193, B1 => n21559, B2 => 
                           n21493, ZN => n7240);
   U18547 : OAI22_X1 port map( A1 => n21502, A2 => n14192, B1 => n21562, B2 => 
                           n21494, ZN => n7241);
   U18548 : OAI22_X1 port map( A1 => n21502, A2 => n14191, B1 => n21565, B2 => 
                           n21494, ZN => n7242);
   U18549 : OAI22_X1 port map( A1 => n21502, A2 => n14190, B1 => n21568, B2 => 
                           n21494, ZN => n7243);
   U18550 : OAI22_X1 port map( A1 => n21502, A2 => n14189, B1 => n21571, B2 => 
                           n21494, ZN => n7244);
   U18551 : OAI22_X1 port map( A1 => n21502, A2 => n14188, B1 => n21574, B2 => 
                           n21494, ZN => n7245);
   U18552 : OAI22_X1 port map( A1 => n21502, A2 => n14187, B1 => n21577, B2 => 
                           n21494, ZN => n7246);
   U18553 : OAI22_X1 port map( A1 => n21502, A2 => n14186, B1 => n21580, B2 => 
                           n21494, ZN => n7247);
   U18554 : OAI22_X1 port map( A1 => n21502, A2 => n14185, B1 => n21583, B2 => 
                           n21494, ZN => n7248);
   U18555 : OAI22_X1 port map( A1 => n21502, A2 => n14184, B1 => n21586, B2 => 
                           n21494, ZN => n7249);
   U18556 : OAI22_X1 port map( A1 => n21502, A2 => n14183, B1 => n21589, B2 => 
                           n21494, ZN => n7250);
   U18557 : OAI22_X1 port map( A1 => n21502, A2 => n14182, B1 => n21592, B2 => 
                           n21494, ZN => n7251);
   U18558 : OAI22_X1 port map( A1 => n21502, A2 => n14181, B1 => n21595, B2 => 
                           n21494, ZN => n7252);
   U18559 : OAI22_X1 port map( A1 => n21502, A2 => n14180, B1 => n21598, B2 => 
                           n21495, ZN => n7253);
   U18560 : OAI22_X1 port map( A1 => n21503, A2 => n14179, B1 => n21601, B2 => 
                           n21495, ZN => n7254);
   U18561 : OAI22_X1 port map( A1 => n21503, A2 => n14178, B1 => n21604, B2 => 
                           n21495, ZN => n7255);
   U18562 : OAI22_X1 port map( A1 => n21503, A2 => n14177, B1 => n21607, B2 => 
                           n21495, ZN => n7256);
   U18563 : OAI22_X1 port map( A1 => n21503, A2 => n14176, B1 => n21610, B2 => 
                           n21495, ZN => n7257);
   U18564 : OAI22_X1 port map( A1 => n21503, A2 => n14175, B1 => n21613, B2 => 
                           n21495, ZN => n7258);
   U18565 : OAI22_X1 port map( A1 => n21503, A2 => n14174, B1 => n21616, B2 => 
                           n21495, ZN => n7259);
   U18566 : OAI22_X1 port map( A1 => n21503, A2 => n14173, B1 => n21619, B2 => 
                           n21495, ZN => n7260);
   U18567 : OAI22_X1 port map( A1 => n21503, A2 => n14172, B1 => n21622, B2 => 
                           n21495, ZN => n7261);
   U18568 : OAI22_X1 port map( A1 => n21503, A2 => n14171, B1 => n21625, B2 => 
                           n21495, ZN => n7262);
   U18569 : OAI22_X1 port map( A1 => n21503, A2 => n14170, B1 => n21628, B2 => 
                           n21495, ZN => n7263);
   U18570 : OAI22_X1 port map( A1 => n21503, A2 => n14169, B1 => n21631, B2 => 
                           n21495, ZN => n7264);
   U18571 : OAI22_X1 port map( A1 => n21503, A2 => n14168, B1 => n21634, B2 => 
                           n21496, ZN => n7265);
   U18572 : OAI22_X1 port map( A1 => n21503, A2 => n14167, B1 => n21637, B2 => 
                           n21496, ZN => n7266);
   U18573 : OAI22_X1 port map( A1 => n21504, A2 => n14166, B1 => n21640, B2 => 
                           n21496, ZN => n7267);
   U18574 : OAI22_X1 port map( A1 => n21504, A2 => n14165, B1 => n21643, B2 => 
                           n21496, ZN => n7268);
   U18575 : OAI22_X1 port map( A1 => n21504, A2 => n14164, B1 => n21646, B2 => 
                           n21496, ZN => n7269);
   U18576 : OAI22_X1 port map( A1 => n21504, A2 => n14163, B1 => n21649, B2 => 
                           n21496, ZN => n7270);
   U18577 : OAI22_X1 port map( A1 => n21504, A2 => n14162, B1 => n21652, B2 => 
                           n21496, ZN => n7271);
   U18578 : OAI22_X1 port map( A1 => n21504, A2 => n14161, B1 => n21655, B2 => 
                           n21496, ZN => n7272);
   U18579 : OAI22_X1 port map( A1 => n21504, A2 => n14160, B1 => n21658, B2 => 
                           n21496, ZN => n7273);
   U18580 : OAI22_X1 port map( A1 => n21504, A2 => n14159, B1 => n21661, B2 => 
                           n21496, ZN => n7274);
   U18581 : OAI22_X1 port map( A1 => n21504, A2 => n14158, B1 => n21664, B2 => 
                           n21496, ZN => n7275);
   U18582 : OAI22_X1 port map( A1 => n21504, A2 => n14157, B1 => n21667, B2 => 
                           n21496, ZN => n7276);
   U18583 : OAI22_X1 port map( A1 => n21504, A2 => n14156, B1 => n21670, B2 => 
                           n21497, ZN => n7277);
   U18584 : OAI22_X1 port map( A1 => n21504, A2 => n14155, B1 => n21673, B2 => 
                           n21497, ZN => n7278);
   U18585 : OAI22_X1 port map( A1 => n21504, A2 => n14154, B1 => n21676, B2 => 
                           n21497, ZN => n7279);
   U18586 : OAI22_X1 port map( A1 => n21505, A2 => n14153, B1 => n21679, B2 => 
                           n21497, ZN => n7280);
   U18587 : OAI22_X1 port map( A1 => n21505, A2 => n14152, B1 => n21682, B2 => 
                           n21497, ZN => n7281);
   U18588 : OAI22_X1 port map( A1 => n21505, A2 => n14151, B1 => n21685, B2 => 
                           n21497, ZN => n7282);
   U18589 : OAI22_X1 port map( A1 => n21505, A2 => n14150, B1 => n21688, B2 => 
                           n21497, ZN => n7283);
   U18590 : OAI22_X1 port map( A1 => n21505, A2 => n14149, B1 => n21691, B2 => 
                           n21497, ZN => n7284);
   U18591 : OAI22_X1 port map( A1 => n21505, A2 => n14148, B1 => n21694, B2 => 
                           n21497, ZN => n7285);
   U18592 : OAI22_X1 port map( A1 => n21505, A2 => n14147, B1 => n21697, B2 => 
                           n21497, ZN => n7286);
   U18593 : OAI22_X1 port map( A1 => n21505, A2 => n14146, B1 => n21700, B2 => 
                           n21497, ZN => n7287);
   U18594 : OAI22_X1 port map( A1 => n21505, A2 => n14145, B1 => n21703, B2 => 
                           n21497, ZN => n7288);
   U18595 : OAI22_X1 port map( A1 => n21726, A2 => n14067, B1 => n21718, B2 => 
                           n21526, ZN => n7357);
   U18596 : OAI22_X1 port map( A1 => n21726, A2 => n14065, B1 => n21718, B2 => 
                           n21529, ZN => n7358);
   U18597 : OAI22_X1 port map( A1 => n21726, A2 => n14063, B1 => n21718, B2 => 
                           n21532, ZN => n7359);
   U18598 : OAI22_X1 port map( A1 => n21726, A2 => n14061, B1 => n21718, B2 => 
                           n21535, ZN => n7360);
   U18599 : OAI22_X1 port map( A1 => n21726, A2 => n14059, B1 => n21718, B2 => 
                           n21538, ZN => n7361);
   U18600 : OAI22_X1 port map( A1 => n21726, A2 => n14057, B1 => n21718, B2 => 
                           n21541, ZN => n7362);
   U18601 : OAI22_X1 port map( A1 => n21726, A2 => n14055, B1 => n21718, B2 => 
                           n21544, ZN => n7363);
   U18602 : OAI22_X1 port map( A1 => n21726, A2 => n14053, B1 => n21718, B2 => 
                           n21547, ZN => n7364);
   U18603 : OAI22_X1 port map( A1 => n21726, A2 => n14051, B1 => n21718, B2 => 
                           n21550, ZN => n7365);
   U18604 : OAI22_X1 port map( A1 => n21726, A2 => n14049, B1 => n21718, B2 => 
                           n21553, ZN => n7366);
   U18605 : OAI22_X1 port map( A1 => n21726, A2 => n14047, B1 => n21718, B2 => 
                           n21556, ZN => n7367);
   U18606 : OAI22_X1 port map( A1 => n21726, A2 => n14045, B1 => n21718, B2 => 
                           n21559, ZN => n7368);
   U18607 : INV_X1 port map( A => ADD_RD2(4), ZN => n18532);
   U18608 : INV_X1 port map( A => ADD_RD1(4), ZN => n17331);
   U18609 : INV_X1 port map( A => ADD_RD2(3), ZN => n18534);
   U18610 : INV_X1 port map( A => ADD_RD1(3), ZN => n17333);
   U18611 : INV_X1 port map( A => ADD_RD2(0), ZN => n18535);
   U18612 : INV_X1 port map( A => ADD_RD1(0), ZN => n17334);
   U18613 : INV_X1 port map( A => DATAIN(0), ZN => n14068);
   U18614 : INV_X1 port map( A => DATAIN(1), ZN => n14066);
   U18615 : INV_X1 port map( A => DATAIN(2), ZN => n14064);
   U18616 : INV_X1 port map( A => DATAIN(3), ZN => n14062);
   U18617 : INV_X1 port map( A => DATAIN(4), ZN => n14060);
   U18618 : INV_X1 port map( A => DATAIN(5), ZN => n14058);
   U18619 : INV_X1 port map( A => DATAIN(6), ZN => n14056);
   U18620 : INV_X1 port map( A => DATAIN(7), ZN => n14054);
   U18621 : INV_X1 port map( A => DATAIN(8), ZN => n14052);
   U18622 : INV_X1 port map( A => DATAIN(9), ZN => n14050);
   U18623 : INV_X1 port map( A => DATAIN(10), ZN => n14048);
   U18624 : INV_X1 port map( A => DATAIN(11), ZN => n14046);
   U18625 : INV_X1 port map( A => DATAIN(12), ZN => n14044);
   U18626 : INV_X1 port map( A => DATAIN(13), ZN => n14042);
   U18627 : INV_X1 port map( A => DATAIN(14), ZN => n14040);
   U18628 : INV_X1 port map( A => DATAIN(15), ZN => n14038);
   U18629 : INV_X1 port map( A => DATAIN(16), ZN => n14036);
   U18630 : INV_X1 port map( A => DATAIN(17), ZN => n14034);
   U18631 : INV_X1 port map( A => DATAIN(18), ZN => n14032);
   U18632 : INV_X1 port map( A => DATAIN(19), ZN => n14030);
   U18633 : INV_X1 port map( A => DATAIN(20), ZN => n14028);
   U18634 : INV_X1 port map( A => DATAIN(21), ZN => n14026);
   U18635 : INV_X1 port map( A => DATAIN(22), ZN => n14024);
   U18636 : INV_X1 port map( A => DATAIN(23), ZN => n14022);
   U18637 : INV_X1 port map( A => DATAIN(24), ZN => n14020);
   U18638 : INV_X1 port map( A => DATAIN(25), ZN => n14018);
   U18639 : INV_X1 port map( A => DATAIN(26), ZN => n14016);
   U18640 : INV_X1 port map( A => DATAIN(27), ZN => n14014);
   U18641 : INV_X1 port map( A => DATAIN(28), ZN => n14012);
   U18642 : INV_X1 port map( A => DATAIN(29), ZN => n14010);
   U18643 : INV_X1 port map( A => DATAIN(30), ZN => n14008);
   U18644 : INV_X1 port map( A => DATAIN(31), ZN => n14006);
   U18645 : INV_X1 port map( A => DATAIN(32), ZN => n14004);
   U18646 : INV_X1 port map( A => DATAIN(33), ZN => n14002);
   U18647 : INV_X1 port map( A => DATAIN(34), ZN => n14000);
   U18648 : INV_X1 port map( A => DATAIN(35), ZN => n13998);
   U18649 : INV_X1 port map( A => DATAIN(36), ZN => n13996);
   U18650 : INV_X1 port map( A => DATAIN(37), ZN => n13994);
   U18651 : INV_X1 port map( A => DATAIN(38), ZN => n13992);
   U18652 : INV_X1 port map( A => DATAIN(39), ZN => n13990);
   U18653 : INV_X1 port map( A => DATAIN(40), ZN => n13988);
   U18654 : INV_X1 port map( A => DATAIN(41), ZN => n13986);
   U18655 : INV_X1 port map( A => DATAIN(42), ZN => n13984);
   U18656 : INV_X1 port map( A => DATAIN(43), ZN => n13982);
   U18657 : INV_X1 port map( A => DATAIN(44), ZN => n13980);
   U18658 : INV_X1 port map( A => DATAIN(45), ZN => n13978);
   U18659 : INV_X1 port map( A => DATAIN(46), ZN => n13976);
   U18660 : INV_X1 port map( A => DATAIN(47), ZN => n13974);
   U18661 : INV_X1 port map( A => DATAIN(48), ZN => n13972);
   U18662 : INV_X1 port map( A => DATAIN(49), ZN => n13970);
   U18663 : INV_X1 port map( A => DATAIN(50), ZN => n13968);
   U18664 : INV_X1 port map( A => DATAIN(51), ZN => n13966);
   U18665 : INV_X1 port map( A => DATAIN(52), ZN => n13964);
   U18666 : INV_X1 port map( A => DATAIN(53), ZN => n13962);
   U18667 : INV_X1 port map( A => DATAIN(54), ZN => n13960);
   U18668 : INV_X1 port map( A => DATAIN(55), ZN => n13958);
   U18669 : INV_X1 port map( A => DATAIN(56), ZN => n13956);
   U18670 : INV_X1 port map( A => DATAIN(57), ZN => n13954);
   U18671 : INV_X1 port map( A => DATAIN(58), ZN => n13952);
   U18672 : INV_X1 port map( A => DATAIN(59), ZN => n13950);
   U18673 : INV_X1 port map( A => DATAIN(60), ZN => n13948);
   U18674 : INV_X1 port map( A => DATAIN(61), ZN => n13946);
   U18675 : INV_X1 port map( A => DATAIN(62), ZN => n13944);
   U18676 : INV_X1 port map( A => DATAIN(63), ZN => n13942);
   U18677 : INV_X1 port map( A => ADD_WR(3), ZN => n14473);
   U18678 : INV_X1 port map( A => ADD_WR(0), ZN => n14472);
   U18679 : INV_X1 port map( A => ADD_WR(1), ZN => n15738);
   U18680 : INV_X1 port map( A => ADD_RD2(1), ZN => n18538);
   U18681 : INV_X1 port map( A => ADD_RD1(1), ZN => n17337);
   U18682 : INV_X1 port map( A => ADD_RD2(2), ZN => n18539);
   U18683 : INV_X1 port map( A => ADD_RD1(2), ZN => n17338);
   U18684 : INV_X1 port map( A => ADD_WR(2), ZN => n15737);
   U18685 : INV_X1 port map( A => RESET, ZN => n14069);
   U18686 : CLKBUF_X1 port map( A => n17388, Z => n20723);
   U18687 : CLKBUF_X1 port map( A => n17387, Z => n20729);
   U18688 : CLKBUF_X1 port map( A => n17385, Z => n20735);
   U18689 : CLKBUF_X1 port map( A => n17384, Z => n20741);
   U18690 : CLKBUF_X1 port map( A => n17383, Z => n20747);
   U18691 : CLKBUF_X1 port map( A => n17382, Z => n20753);
   U18692 : CLKBUF_X1 port map( A => n17380, Z => n20759);
   U18693 : CLKBUF_X1 port map( A => n17379, Z => n20765);
   U18694 : CLKBUF_X1 port map( A => n17378, Z => n20771);
   U18695 : CLKBUF_X1 port map( A => n17377, Z => n20777);
   U18696 : CLKBUF_X1 port map( A => n17375, Z => n20783);
   U18697 : CLKBUF_X1 port map( A => n17374, Z => n20789);
   U18698 : CLKBUF_X1 port map( A => n17373, Z => n20795);
   U18699 : CLKBUF_X1 port map( A => n17371, Z => n20801);
   U18700 : CLKBUF_X1 port map( A => n17370, Z => n20807);
   U18701 : CLKBUF_X1 port map( A => n17365, Z => n20813);
   U18702 : CLKBUF_X1 port map( A => n17364, Z => n20819);
   U18703 : CLKBUF_X1 port map( A => n17363, Z => n20825);
   U18704 : CLKBUF_X1 port map( A => n17361, Z => n20831);
   U18705 : CLKBUF_X1 port map( A => n17360, Z => n20837);
   U18706 : CLKBUF_X1 port map( A => n17359, Z => n20843);
   U18707 : CLKBUF_X1 port map( A => n17358, Z => n20849);
   U18708 : CLKBUF_X1 port map( A => n17356, Z => n20855);
   U18709 : CLKBUF_X1 port map( A => n17355, Z => n20861);
   U18710 : CLKBUF_X1 port map( A => n17354, Z => n20867);
   U18711 : CLKBUF_X1 port map( A => n17353, Z => n20873);
   U18712 : CLKBUF_X1 port map( A => n17351, Z => n20879);
   U18713 : CLKBUF_X1 port map( A => n17350, Z => n20885);
   U18714 : CLKBUF_X1 port map( A => n17349, Z => n20891);
   U18715 : CLKBUF_X1 port map( A => n17348, Z => n20897);
   U18716 : CLKBUF_X1 port map( A => n17346, Z => n20903);
   U18717 : CLKBUF_X1 port map( A => n17345, Z => n20909);
   U18718 : CLKBUF_X1 port map( A => n16123, Z => n20915);
   U18719 : CLKBUF_X1 port map( A => n16122, Z => n20921);
   U18720 : CLKBUF_X1 port map( A => n16120, Z => n20927);
   U18721 : CLKBUF_X1 port map( A => n16119, Z => n20933);
   U18722 : CLKBUF_X1 port map( A => n16118, Z => n20939);
   U18723 : CLKBUF_X1 port map( A => n16117, Z => n20945);
   U18724 : CLKBUF_X1 port map( A => n16115, Z => n20951);
   U18725 : CLKBUF_X1 port map( A => n16114, Z => n20957);
   U18726 : CLKBUF_X1 port map( A => n16113, Z => n20963);
   U18727 : CLKBUF_X1 port map( A => n16112, Z => n20969);
   U18728 : CLKBUF_X1 port map( A => n16110, Z => n20975);
   U18729 : CLKBUF_X1 port map( A => n16109, Z => n20981);
   U18730 : CLKBUF_X1 port map( A => n20983, Z => n20994);
   U18731 : CLKBUF_X1 port map( A => n16107, Z => n21000);
   U18732 : CLKBUF_X1 port map( A => n16105, Z => n21006);
   U18733 : CLKBUF_X1 port map( A => n16104, Z => n21012);
   U18734 : CLKBUF_X1 port map( A => n16099, Z => n21018);
   U18735 : CLKBUF_X1 port map( A => n16098, Z => n21024);
   U18736 : CLKBUF_X1 port map( A => n16097, Z => n21030);
   U18737 : CLKBUF_X1 port map( A => n16095, Z => n21036);
   U18738 : CLKBUF_X1 port map( A => n16094, Z => n21042);
   U18739 : CLKBUF_X1 port map( A => n16093, Z => n21048);
   U18740 : CLKBUF_X1 port map( A => n16092, Z => n21054);
   U18741 : CLKBUF_X1 port map( A => n16090, Z => n21060);
   U18742 : CLKBUF_X1 port map( A => n16089, Z => n21066);
   U18743 : CLKBUF_X1 port map( A => n16088, Z => n21072);
   U18744 : CLKBUF_X1 port map( A => n16087, Z => n21078);
   U18745 : CLKBUF_X1 port map( A => n16084, Z => n21091);
   U18746 : CLKBUF_X1 port map( A => n16082, Z => n21097);
   U18747 : CLKBUF_X1 port map( A => n16081, Z => n21103);
   U18748 : CLKBUF_X1 port map( A => n16079, Z => n21109);
   U18749 : CLKBUF_X1 port map( A => n16078, Z => n21115);
   U18750 : CLKBUF_X1 port map( A => n16071, Z => n21121);
   U18751 : CLKBUF_X1 port map( A => n16005, Z => n21134);
   U18752 : CLKBUF_X1 port map( A => n15939, Z => n21147);
   U18753 : CLKBUF_X1 port map( A => n15873, Z => n21160);
   U18754 : CLKBUF_X1 port map( A => n15807, Z => n21173);
   U18755 : CLKBUF_X1 port map( A => n15741, Z => n21186);
   U18756 : CLKBUF_X1 port map( A => n15672, Z => n21199);
   U18757 : CLKBUF_X1 port map( A => n15605, Z => n21212);
   U18758 : CLKBUF_X1 port map( A => n15539, Z => n21225);
   U18759 : CLKBUF_X1 port map( A => n15472, Z => n21238);
   U18760 : CLKBUF_X1 port map( A => n15406, Z => n21251);
   U18761 : CLKBUF_X1 port map( A => n15340, Z => n21264);
   U18762 : CLKBUF_X1 port map( A => n15274, Z => n21277);
   U18763 : CLKBUF_X1 port map( A => n15208, Z => n21290);
   U18764 : CLKBUF_X1 port map( A => n15141, Z => n21303);
   U18765 : CLKBUF_X1 port map( A => n15074, Z => n21316);
   U18766 : CLKBUF_X1 port map( A => n15007, Z => n21329);
   U18767 : CLKBUF_X1 port map( A => n14941, Z => n21342);
   U18768 : CLKBUF_X1 port map( A => n14875, Z => n21355);
   U18769 : CLKBUF_X1 port map( A => n14809, Z => n21368);
   U18770 : CLKBUF_X1 port map( A => n14743, Z => n21381);
   U18771 : CLKBUF_X1 port map( A => n14677, Z => n21394);
   U18772 : CLKBUF_X1 port map( A => n14610, Z => n21407);
   U18773 : CLKBUF_X1 port map( A => n14543, Z => n21420);
   U18774 : CLKBUF_X1 port map( A => n14477, Z => n21433);
   U18775 : CLKBUF_X1 port map( A => n14407, Z => n21446);
   U18776 : CLKBUF_X1 port map( A => n14341, Z => n21459);
   U18777 : CLKBUF_X1 port map( A => n14274, Z => n21472);
   U18778 : CLKBUF_X1 port map( A => n14208, Z => n21485);
   U18779 : CLKBUF_X1 port map( A => n14141, Z => n21498);
   U18780 : CLKBUF_X1 port map( A => n14074, Z => n21511);
   U18781 : CLKBUF_X1 port map( A => n13941, Z => n21723);

end SYN_BEHAVIORAL;
