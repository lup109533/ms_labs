
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_BOOTHMUL_N32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_BOOTHMUL_N32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_1007 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1007;

architecture SYN_BEHAVIORAL of FA_1007 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net148762, net148733, net138080, n3, n4, n5 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n4);
   U2 : NAND2_X1 port map( A1 => n4, A2 => net138080, ZN => Co);
   U3 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : CLKBUF_X1 port map( A => A, Z => net148733);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U7 : CLKBUF_X1 port map( A => B, Z => net148762);
   U8 : NAND2_X1 port map( A1 => net148733, A2 => net148762, ZN => net138080);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_1006 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1006;

architecture SYN_BEHAVIORAL of FA_1006 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_1005 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1005;

architecture SYN_BEHAVIORAL of FA_1005 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_1004 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1004;

architecture SYN_BEHAVIORAL of FA_1004 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_1003 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1003;

architecture SYN_BEHAVIORAL of FA_1003 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_1002 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1002;

architecture SYN_BEHAVIORAL of FA_1002 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_1001 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1001;

architecture SYN_BEHAVIORAL of FA_1001 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_1000 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1000;

architecture SYN_BEHAVIORAL of FA_1000 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_999 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_999;

architecture SYN_BEHAVIORAL of FA_999 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_998 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_998;

architecture SYN_BEHAVIORAL of FA_998 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_997 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_997;

architecture SYN_BEHAVIORAL of FA_997 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_996 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_996;

architecture SYN_BEHAVIORAL of FA_996 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_995 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_995;

architecture SYN_BEHAVIORAL of FA_995 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_994 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_994;

architecture SYN_BEHAVIORAL of FA_994 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_993 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_993;

architecture SYN_BEHAVIORAL of FA_993 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_992 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_992;

architecture SYN_BEHAVIORAL of FA_992 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_991 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_991;

architecture SYN_BEHAVIORAL of FA_991 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_990 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_990;

architecture SYN_BEHAVIORAL of FA_990 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_989 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_989;

architecture SYN_BEHAVIORAL of FA_989 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_988 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_988;

architecture SYN_BEHAVIORAL of FA_988 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_987 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_987;

architecture SYN_BEHAVIORAL of FA_987 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_986 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_986;

architecture SYN_BEHAVIORAL of FA_986 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_985 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_985;

architecture SYN_BEHAVIORAL of FA_985 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_984 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_984;

architecture SYN_BEHAVIORAL of FA_984 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net137989, net137988, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net137989);
   U2 : NAND2_X1 port map( A1 => net137989, A2 => net137988, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n4);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137988);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_983 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_983;

architecture SYN_BEHAVIORAL of FA_983 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_982 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_982;

architecture SYN_BEHAVIORAL of FA_982 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_981 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_981;

architecture SYN_BEHAVIORAL of FA_981 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_980 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_980;

architecture SYN_BEHAVIORAL of FA_980 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_979 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_979;

architecture SYN_BEHAVIORAL of FA_979 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_978 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_978;

architecture SYN_BEHAVIORAL of FA_978 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_977 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_977;

architecture SYN_BEHAVIORAL of FA_977 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_976 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_976;

architecture SYN_BEHAVIORAL of FA_976 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_975 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_975;

architecture SYN_BEHAVIORAL of FA_975 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_974 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_974;

architecture SYN_BEHAVIORAL of FA_974 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_973 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_973;

architecture SYN_BEHAVIORAL of FA_973 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_972 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_972;

architecture SYN_BEHAVIORAL of FA_972 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_971 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_971;

architecture SYN_BEHAVIORAL of FA_971 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_970 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_970;

architecture SYN_BEHAVIORAL of FA_970 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_969 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_969;

architecture SYN_BEHAVIORAL of FA_969 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_968 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_968;

architecture SYN_BEHAVIORAL of FA_968 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_967 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_967;

architecture SYN_BEHAVIORAL of FA_967 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_966 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_966;

architecture SYN_BEHAVIORAL of FA_966 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_965 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_965;

architecture SYN_BEHAVIORAL of FA_965 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net137913, net137912, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net137913);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U4 : INV_X1 port map( A => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137912);
   U6 : NAND2_X1 port map( A1 => net137913, A2 => net137912, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_964 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_964;

architecture SYN_BEHAVIORAL of FA_964 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_963 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_963;

architecture SYN_BEHAVIORAL of FA_963 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_962 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_962;

architecture SYN_BEHAVIORAL of FA_962 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : INV_X1 port map( A => n3, ZN => n6);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_961 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_961;

architecture SYN_BEHAVIORAL of FA_961 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : INV_X1 port map( A => n3, ZN => n6);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_960 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_960;

architecture SYN_BEHAVIORAL of FA_960 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_959 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_959;

architecture SYN_BEHAVIORAL of FA_959 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : INV_X1 port map( A => n3, ZN => n6);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_958 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_958;

architecture SYN_BEHAVIORAL of FA_958 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_957 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_957;

architecture SYN_BEHAVIORAL of FA_957 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_956 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_956;

architecture SYN_BEHAVIORAL of FA_956 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_955 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_955;

architecture SYN_BEHAVIORAL of FA_955 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_954 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_954;

architecture SYN_BEHAVIORAL of FA_954 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_953 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_953;

architecture SYN_BEHAVIORAL of FA_953 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_952 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_952;

architecture SYN_BEHAVIORAL of FA_952 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : INV_X1 port map( A => n3, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_951 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_951;

architecture SYN_BEHAVIORAL of FA_951 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net137856, net137857, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net137857);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U4 : INV_X1 port map( A => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137856);
   U6 : NAND2_X1 port map( A1 => net137856, A2 => net137857, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_950 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_950;

architecture SYN_BEHAVIORAL of FA_950 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_949 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_949;

architecture SYN_BEHAVIORAL of FA_949 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_948 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_948;

architecture SYN_BEHAVIORAL of FA_948 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_947 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_947;

architecture SYN_BEHAVIORAL of FA_947 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_946 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_946;

architecture SYN_BEHAVIORAL of FA_946 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_945 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_945;

architecture SYN_BEHAVIORAL of FA_945 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_944 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_944;

architecture SYN_BEHAVIORAL of FA_944 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n5, B2 => n6, A => n4, ZN => Co);
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : CLKBUF_X1 port map( A => B, Z => n3);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_943 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_943;

architecture SYN_BEHAVIORAL of FA_943 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_942 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_942;

architecture SYN_BEHAVIORAL of FA_942 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_941 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_941;

architecture SYN_BEHAVIORAL of FA_941 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_940 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_940;

architecture SYN_BEHAVIORAL of FA_940 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_939 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_939;

architecture SYN_BEHAVIORAL of FA_939 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_938 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_938;

architecture SYN_BEHAVIORAL of FA_938 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_937 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_937;

architecture SYN_BEHAVIORAL of FA_937 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_936 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_936;

architecture SYN_BEHAVIORAL of FA_936 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_935 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_935;

architecture SYN_BEHAVIORAL of FA_935 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_934 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_934;

architecture SYN_BEHAVIORAL of FA_934 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_933 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_933;

architecture SYN_BEHAVIORAL of FA_933 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_932 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_932;

architecture SYN_BEHAVIORAL of FA_932 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_931 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_931;

architecture SYN_BEHAVIORAL of FA_931 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_930 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_930;

architecture SYN_BEHAVIORAL of FA_930 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_929 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_929;

architecture SYN_BEHAVIORAL of FA_929 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_928 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_928;

architecture SYN_BEHAVIORAL of FA_928 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_927 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_927;

architecture SYN_BEHAVIORAL of FA_927 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_926 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_926;

architecture SYN_BEHAVIORAL of FA_926 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_925 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_925;

architecture SYN_BEHAVIORAL of FA_925 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_924 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_924;

architecture SYN_BEHAVIORAL of FA_924 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_923 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_923;

architecture SYN_BEHAVIORAL of FA_923 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_922 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_922;

architecture SYN_BEHAVIORAL of FA_922 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_921 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_921;

architecture SYN_BEHAVIORAL of FA_921 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_920 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_920;

architecture SYN_BEHAVIORAL of FA_920 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net137734, net137732, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => net137734);
   U3 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U4 : CLKBUF_X1 port map( A => B, Z => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => net137732);
   U6 : NAND2_X1 port map( A1 => n5, A2 => net137732, ZN => Co);
   U7 : NAND2_X1 port map( A1 => net137734, A2 => Ci, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_919 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_919;

architecture SYN_BEHAVIORAL of FA_919 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_918 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_918;

architecture SYN_BEHAVIORAL of FA_918 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net137724, net137725, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net137725);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137724);
   U5 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U6 : NAND2_X1 port map( A1 => net137725, A2 => net137724, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_917 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_917;

architecture SYN_BEHAVIORAL of FA_917 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_916 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_916;

architecture SYN_BEHAVIORAL of FA_916 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_915 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_915;

architecture SYN_BEHAVIORAL of FA_915 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_914 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_914;

architecture SYN_BEHAVIORAL of FA_914 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_913 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_913;

architecture SYN_BEHAVIORAL of FA_913 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_912 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_912;

architecture SYN_BEHAVIORAL of FA_912 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : BUF_X1 port map( A => n8, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_911 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_911;

architecture SYN_BEHAVIORAL of FA_911 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_910 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_910;

architecture SYN_BEHAVIORAL of FA_910 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_909 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_909;

architecture SYN_BEHAVIORAL of FA_909 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_908 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_908;

architecture SYN_BEHAVIORAL of FA_908 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_907 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_907;

architecture SYN_BEHAVIORAL of FA_907 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_906 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_906;

architecture SYN_BEHAVIORAL of FA_906 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_905 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_905;

architecture SYN_BEHAVIORAL of FA_905 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_904 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_904;

architecture SYN_BEHAVIORAL of FA_904 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_903 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_903;

architecture SYN_BEHAVIORAL of FA_903 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_902 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_902;

architecture SYN_BEHAVIORAL of FA_902 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_901 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_901;

architecture SYN_BEHAVIORAL of FA_901 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net137656, net137657, net137658, n3, n4 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : INV_X1 port map( A => n4, ZN => net137658);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => net137656);
   U5 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => net137658, ZN => net137657);
   U7 : NAND2_X1 port map( A1 => net137656, A2 => net137657, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_900 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_900;

architecture SYN_BEHAVIORAL of FA_900 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_899 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_899;

architecture SYN_BEHAVIORAL of FA_899 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_898 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_898;

architecture SYN_BEHAVIORAL of FA_898 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_897 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_897;

architecture SYN_BEHAVIORAL of FA_897 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_896 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_896;

architecture SYN_BEHAVIORAL of FA_896 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_895 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_895;

architecture SYN_BEHAVIORAL of FA_895 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_894 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_894;

architecture SYN_BEHAVIORAL of FA_894 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_893 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_893;

architecture SYN_BEHAVIORAL of FA_893 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_892 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_892;

architecture SYN_BEHAVIORAL of FA_892 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_891 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_891;

architecture SYN_BEHAVIORAL of FA_891 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_890 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_890;

architecture SYN_BEHAVIORAL of FA_890 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_889 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_889;

architecture SYN_BEHAVIORAL of FA_889 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_888 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_888;

architecture SYN_BEHAVIORAL of FA_888 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_887 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_887;

architecture SYN_BEHAVIORAL of FA_887 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net137600, n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : NAND2_X1 port map( A1 => net137600, A2 => n5, ZN => Co);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137600);
   U5 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_886 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_886;

architecture SYN_BEHAVIORAL of FA_886 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net137596, net137597, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net137597);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U4 : INV_X1 port map( A => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137596);
   U6 : NAND2_X1 port map( A1 => net137596, A2 => net137597, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_885 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_885;

architecture SYN_BEHAVIORAL of FA_885 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_884 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_884;

architecture SYN_BEHAVIORAL of FA_884 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_883 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_883;

architecture SYN_BEHAVIORAL of FA_883 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_882 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_882;

architecture SYN_BEHAVIORAL of FA_882 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_881 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_881;

architecture SYN_BEHAVIORAL of FA_881 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_880 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_880;

architecture SYN_BEHAVIORAL of FA_880 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_879 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_879;

architecture SYN_BEHAVIORAL of FA_879 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_878 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_878;

architecture SYN_BEHAVIORAL of FA_878 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_877 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_877;

architecture SYN_BEHAVIORAL of FA_877 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_876 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_876;

architecture SYN_BEHAVIORAL of FA_876 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_875 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_875;

architecture SYN_BEHAVIORAL of FA_875 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_874 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_874;

architecture SYN_BEHAVIORAL of FA_874 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_873 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_873;

architecture SYN_BEHAVIORAL of FA_873 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_872 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_872;

architecture SYN_BEHAVIORAL of FA_872 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_871 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_871;

architecture SYN_BEHAVIORAL of FA_871 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_870 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_870;

architecture SYN_BEHAVIORAL of FA_870 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_869 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_869;

architecture SYN_BEHAVIORAL of FA_869 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_868 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_868;

architecture SYN_BEHAVIORAL of FA_868 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_867 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_867;

architecture SYN_BEHAVIORAL of FA_867 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_866 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_866;

architecture SYN_BEHAVIORAL of FA_866 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_865 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_865;

architecture SYN_BEHAVIORAL of FA_865 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_864 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_864;

architecture SYN_BEHAVIORAL of FA_864 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_863 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_863;

architecture SYN_BEHAVIORAL of FA_863 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_862 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_862;

architecture SYN_BEHAVIORAL of FA_862 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_861 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_861;

architecture SYN_BEHAVIORAL of FA_861 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_860 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_860;

architecture SYN_BEHAVIORAL of FA_860 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_859 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_859;

architecture SYN_BEHAVIORAL of FA_859 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_858 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_858;

architecture SYN_BEHAVIORAL of FA_858 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_857 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_857;

architecture SYN_BEHAVIORAL of FA_857 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_856 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_856;

architecture SYN_BEHAVIORAL of FA_856 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_855 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_855;

architecture SYN_BEHAVIORAL of FA_855 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_854 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_854;

architecture SYN_BEHAVIORAL of FA_854 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net137468, n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137468);
   U5 : NAND2_X1 port map( A1 => n5, A2 => net137468, ZN => Co);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_853 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_853;

architecture SYN_BEHAVIORAL of FA_853 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net137464, net137465, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => net137465);
   U5 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => net137464);
   U6 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U7 : NAND2_X1 port map( A1 => net137465, A2 => net137464, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_852 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_852;

architecture SYN_BEHAVIORAL of FA_852 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_851 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_851;

architecture SYN_BEHAVIORAL of FA_851 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_850 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_850;

architecture SYN_BEHAVIORAL of FA_850 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_849 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_849;

architecture SYN_BEHAVIORAL of FA_849 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_848 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_848;

architecture SYN_BEHAVIORAL of FA_848 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_847 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_847;

architecture SYN_BEHAVIORAL of FA_847 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_846 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_846;

architecture SYN_BEHAVIORAL of FA_846 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_845 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_845;

architecture SYN_BEHAVIORAL of FA_845 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_844 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_844;

architecture SYN_BEHAVIORAL of FA_844 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_843 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_843;

architecture SYN_BEHAVIORAL of FA_843 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_842 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_842;

architecture SYN_BEHAVIORAL of FA_842 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_841 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_841;

architecture SYN_BEHAVIORAL of FA_841 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_840 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_840;

architecture SYN_BEHAVIORAL of FA_840 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_839 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_839;

architecture SYN_BEHAVIORAL of FA_839 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_838 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_838;

architecture SYN_BEHAVIORAL of FA_838 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_837 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_837;

architecture SYN_BEHAVIORAL of FA_837 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net137401, net137400, net137399, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net137401);
   U2 : NAND2_X1 port map( A1 => net137401, A2 => net137400, ZN => Co);
   U3 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U4 : XNOR2_X1 port map( A => Ci, B => net137399, ZN => S);
   U5 : XNOR2_X1 port map( A => A, B => B, ZN => net137399);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137400);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_836 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_836;

architecture SYN_BEHAVIORAL of FA_836 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_835 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_835;

architecture SYN_BEHAVIORAL of FA_835 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U3 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_834 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_834;

architecture SYN_BEHAVIORAL of FA_834 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net137388, net137389, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net137389);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137388);
   U6 : NAND2_X1 port map( A1 => net137389, A2 => net137388, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_833 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_833;

architecture SYN_BEHAVIORAL of FA_833 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_832 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_832;

architecture SYN_BEHAVIORAL of FA_832 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_831 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_831;

architecture SYN_BEHAVIORAL of FA_831 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_830 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_830;

architecture SYN_BEHAVIORAL of FA_830 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_829 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_829;

architecture SYN_BEHAVIORAL of FA_829 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_828 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_828;

architecture SYN_BEHAVIORAL of FA_828 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_827 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_827;

architecture SYN_BEHAVIORAL of FA_827 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_826 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_826;

architecture SYN_BEHAVIORAL of FA_826 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_825 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_825;

architecture SYN_BEHAVIORAL of FA_825 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_824 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_824;

architecture SYN_BEHAVIORAL of FA_824 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_823 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_823;

architecture SYN_BEHAVIORAL of FA_823 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_822 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_822;

architecture SYN_BEHAVIORAL of FA_822 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net137340, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => net137340, A2 => n6, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137340);
   U6 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_821 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_821;

architecture SYN_BEHAVIORAL of FA_821 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net137336, net137337, n3, n4 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net137337);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137336);
   U6 : NAND2_X1 port map( A1 => net137336, A2 => net137337, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_820 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_820;

architecture SYN_BEHAVIORAL of FA_820 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_819 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_819;

architecture SYN_BEHAVIORAL of FA_819 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_818 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_818;

architecture SYN_BEHAVIORAL of FA_818 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_817 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_817;

architecture SYN_BEHAVIORAL of FA_817 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_816 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_816;

architecture SYN_BEHAVIORAL of FA_816 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : OAI21_X1 port map( B1 => n5, B2 => n4, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_815 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_815;

architecture SYN_BEHAVIORAL of FA_815 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_814 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_814;

architecture SYN_BEHAVIORAL of FA_814 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_813 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_813;

architecture SYN_BEHAVIORAL of FA_813 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_812 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_812;

architecture SYN_BEHAVIORAL of FA_812 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_811 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_811;

architecture SYN_BEHAVIORAL of FA_811 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_810 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_810;

architecture SYN_BEHAVIORAL of FA_810 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_809 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_809;

architecture SYN_BEHAVIORAL of FA_809 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_808 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_808;

architecture SYN_BEHAVIORAL of FA_808 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_807 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_807;

architecture SYN_BEHAVIORAL of FA_807 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_806 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_806;

architecture SYN_BEHAVIORAL of FA_806 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_805 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_805;

architecture SYN_BEHAVIORAL of FA_805 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_804 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_804;

architecture SYN_BEHAVIORAL of FA_804 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_803 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_803;

architecture SYN_BEHAVIORAL of FA_803 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_802 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_802;

architecture SYN_BEHAVIORAL of FA_802 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XOR2_X1 port map( A => Ci, B => n4, Z => S);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_801 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_801;

architecture SYN_BEHAVIORAL of FA_801 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_800 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_800;

architecture SYN_BEHAVIORAL of FA_800 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_799 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_799;

architecture SYN_BEHAVIORAL of FA_799 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_798 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_798;

architecture SYN_BEHAVIORAL of FA_798 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_797 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_797;

architecture SYN_BEHAVIORAL of FA_797 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_796 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_796;

architecture SYN_BEHAVIORAL of FA_796 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_795 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_795;

architecture SYN_BEHAVIORAL of FA_795 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_794 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_794;

architecture SYN_BEHAVIORAL of FA_794 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_793 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_793;

architecture SYN_BEHAVIORAL of FA_793 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_792 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_792;

architecture SYN_BEHAVIORAL of FA_792 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_791 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_791;

architecture SYN_BEHAVIORAL of FA_791 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_790 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_790;

architecture SYN_BEHAVIORAL of FA_790 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_789 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_789;

architecture SYN_BEHAVIORAL of FA_789 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net137210, net137208, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U2 : INV_X1 port map( A => n3, ZN => net137210);
   U3 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);
   U4 : CLKBUF_X1 port map( A => B, Z => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => net137208);
   U6 : NAND2_X1 port map( A1 => n5, A2 => net137208, ZN => Co);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => net137210, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_788 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_788;

architecture SYN_BEHAVIORAL of FA_788 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_787 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_787;

architecture SYN_BEHAVIORAL of FA_787 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net137200, net137201, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => net137201);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => net137200);
   U6 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U7 : NAND2_X1 port map( A1 => net137201, A2 => net137200, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_786 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_786;

architecture SYN_BEHAVIORAL of FA_786 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_785 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_785;

architecture SYN_BEHAVIORAL of FA_785 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_784 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_784;

architecture SYN_BEHAVIORAL of FA_784 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_783 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_783;

architecture SYN_BEHAVIORAL of FA_783 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_782 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_782;

architecture SYN_BEHAVIORAL of FA_782 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_781 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_781;

architecture SYN_BEHAVIORAL of FA_781 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_780 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_780;

architecture SYN_BEHAVIORAL of FA_780 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_779 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_779;

architecture SYN_BEHAVIORAL of FA_779 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_778 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_778;

architecture SYN_BEHAVIORAL of FA_778 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_777 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_777;

architecture SYN_BEHAVIORAL of FA_777 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_776 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_776;

architecture SYN_BEHAVIORAL of FA_776 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_775 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_775;

architecture SYN_BEHAVIORAL of FA_775 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_774 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_774;

architecture SYN_BEHAVIORAL of FA_774 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_773 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_773;

architecture SYN_BEHAVIORAL of FA_773 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_772 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_772;

architecture SYN_BEHAVIORAL of FA_772 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_771 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_771;

architecture SYN_BEHAVIORAL of FA_771 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_770 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_770;

architecture SYN_BEHAVIORAL of FA_770 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net137133, net137132, net137131, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net137133);
   U2 : NAND2_X1 port map( A1 => net137133, A2 => net137132, ZN => Co);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U4 : XNOR2_X1 port map( A => Ci, B => net137131, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => net137131);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net137132);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_769 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_769;

architecture SYN_BEHAVIORAL of FA_769 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_768 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_768;

architecture SYN_BEHAVIORAL of FA_768 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_767 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_767;

architecture SYN_BEHAVIORAL of FA_767 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U6 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_766 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_766;

architecture SYN_BEHAVIORAL of FA_766 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U4 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U6 : CLKBUF_X1 port map( A => B, Z => n7);
   U7 : NAND2_X1 port map( A1 => A, A2 => n7, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_765 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_765;

architecture SYN_BEHAVIORAL of FA_765 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_764 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_764;

architecture SYN_BEHAVIORAL of FA_764 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_763 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_763;

architecture SYN_BEHAVIORAL of FA_763 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U3 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_762 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_762;

architecture SYN_BEHAVIORAL of FA_762 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n7);
   U5 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U6 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n5);
   U7 : XNOR2_X1 port map( A => A, B => B, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_761 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_761;

architecture SYN_BEHAVIORAL of FA_761 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n6, A2 => Ci, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_760 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_760;

architecture SYN_BEHAVIORAL of FA_760 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net137092, net137093, n3, n4 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net137093);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net137092);
   U6 : NAND2_X1 port map( A1 => net137093, A2 => net137092, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_759 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_759;

architecture SYN_BEHAVIORAL of FA_759 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_758 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_758;

architecture SYN_BEHAVIORAL of FA_758 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_757 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_757;

architecture SYN_BEHAVIORAL of FA_757 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net137080, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => net137080, A2 => n6, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137080);
   U6 : XNOR2_X1 port map( A => Ci, B => n5, ZN => S);
   U7 : XNOR2_X1 port map( A => A, B => B, ZN => n5);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_756 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_756;

architecture SYN_BEHAVIORAL of FA_756 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net137076, net137077, n3, n4 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net137077);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net137076);
   U6 : NAND2_X1 port map( A1 => net137076, A2 => net137077, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_755 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_755;

architecture SYN_BEHAVIORAL of FA_755 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_754 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_754;

architecture SYN_BEHAVIORAL of FA_754 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_753 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_753;

architecture SYN_BEHAVIORAL of FA_753 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_752 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_752;

architecture SYN_BEHAVIORAL of FA_752 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U3 : OAI21_X1 port map( B1 => n6, B2 => n5, A => n4, ZN => Co);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U5 : INV_X1 port map( A => Ci, ZN => n6);
   U6 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_751 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_751;

architecture SYN_BEHAVIORAL of FA_751 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_750 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_750;

architecture SYN_BEHAVIORAL of FA_750 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => n8, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_749 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_749;

architecture SYN_BEHAVIORAL of FA_749 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_748 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_748;

architecture SYN_BEHAVIORAL of FA_748 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_747 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_747;

architecture SYN_BEHAVIORAL of FA_747 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_746 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_746;

architecture SYN_BEHAVIORAL of FA_746 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_745 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_745;

architecture SYN_BEHAVIORAL of FA_745 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_744 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_744;

architecture SYN_BEHAVIORAL of FA_744 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_743 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_743;

architecture SYN_BEHAVIORAL of FA_743 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_742 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_742;

architecture SYN_BEHAVIORAL of FA_742 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_741 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_741;

architecture SYN_BEHAVIORAL of FA_741 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_740 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_740;

architecture SYN_BEHAVIORAL of FA_740 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_739 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_739;

architecture SYN_BEHAVIORAL of FA_739 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_738 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_738;

architecture SYN_BEHAVIORAL of FA_738 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => n8, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_737 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_737;

architecture SYN_BEHAVIORAL of FA_737 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_736 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_736;

architecture SYN_BEHAVIORAL of FA_736 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_735 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_735;

architecture SYN_BEHAVIORAL of FA_735 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_734 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_734;

architecture SYN_BEHAVIORAL of FA_734 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_733 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_733;

architecture SYN_BEHAVIORAL of FA_733 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_732 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_732;

architecture SYN_BEHAVIORAL of FA_732 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_731 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_731;

architecture SYN_BEHAVIORAL of FA_731 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_730 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_730;

architecture SYN_BEHAVIORAL of FA_730 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_729 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_729;

architecture SYN_BEHAVIORAL of FA_729 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_728 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_728;

architecture SYN_BEHAVIORAL of FA_728 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_727 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_727;

architecture SYN_BEHAVIORAL of FA_727 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_726 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_726;

architecture SYN_BEHAVIORAL of FA_726 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_725 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_725;

architecture SYN_BEHAVIORAL of FA_725 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_724 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_724;

architecture SYN_BEHAVIORAL of FA_724 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_723 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_723;

architecture SYN_BEHAVIORAL of FA_723 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136945, net136944, net148804, net136943, n3 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => net136943, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => net136943);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => net148804, ZN => net136945);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136944);
   U6 : XNOR2_X1 port map( A => B, B => n3, ZN => net148804);
   U7 : NAND2_X1 port map( A1 => net136945, A2 => net136944, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_722 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_722;

architecture SYN_BEHAVIORAL of FA_722 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U7 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_721 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_721;

architecture SYN_BEHAVIORAL of FA_721 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n7);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U7 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_720 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_720;

architecture SYN_BEHAVIORAL of FA_720 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U3 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U5 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U7 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_719 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_719;

architecture SYN_BEHAVIORAL of FA_719 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_718 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_718;

architecture SYN_BEHAVIORAL of FA_718 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_717 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_717;

architecture SYN_BEHAVIORAL of FA_717 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136920, net136921, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net136921);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136920);
   U6 : NAND2_X1 port map( A1 => net136921, A2 => net136920, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_716 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_716;

architecture SYN_BEHAVIORAL of FA_716 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_715 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_715;

architecture SYN_BEHAVIORAL of FA_715 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_714 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_714;

architecture SYN_BEHAVIORAL of FA_714 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_713 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_713;

architecture SYN_BEHAVIORAL of FA_713 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_712 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_712;

architecture SYN_BEHAVIORAL of FA_712 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_711 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_711;

architecture SYN_BEHAVIORAL of FA_711 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_710 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_710;

architecture SYN_BEHAVIORAL of FA_710 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_709 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_709;

architecture SYN_BEHAVIORAL of FA_709 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_708 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_708;

architecture SYN_BEHAVIORAL of FA_708 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_707 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_707;

architecture SYN_BEHAVIORAL of FA_707 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_706 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_706;

architecture SYN_BEHAVIORAL of FA_706 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_705 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_705;

architecture SYN_BEHAVIORAL of FA_705 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_704 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_704;

architecture SYN_BEHAVIORAL of FA_704 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_703 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_703;

architecture SYN_BEHAVIORAL of FA_703 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_702 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_702;

architecture SYN_BEHAVIORAL of FA_702 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_701 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_701;

architecture SYN_BEHAVIORAL of FA_701 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_700 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_700;

architecture SYN_BEHAVIORAL of FA_700 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_699 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_699;

architecture SYN_BEHAVIORAL of FA_699 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_698 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_698;

architecture SYN_BEHAVIORAL of FA_698 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_697 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_697;

architecture SYN_BEHAVIORAL of FA_697 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_696 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_696;

architecture SYN_BEHAVIORAL of FA_696 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136837, net136836, net136835, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net136837);
   U2 : NAND2_X1 port map( A1 => net136836, A2 => net136837, ZN => Co);
   U3 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U4 : XNOR2_X1 port map( A => Ci, B => net136835, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => net136835);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net136836);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_695 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_695;

architecture SYN_BEHAVIORAL of FA_695 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U3 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U4 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U5 : NAND2_X1 port map( A1 => A, A2 => n7, ZN => n4);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U7 : CLKBUF_X1 port map( A => B, Z => n7);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_694 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_694;

architecture SYN_BEHAVIORAL of FA_694 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136828, net136829, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net136829);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136828);
   U6 : NAND2_X1 port map( A1 => net136829, A2 => net136828, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_693 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_693;

architecture SYN_BEHAVIORAL of FA_693 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_692 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_692;

architecture SYN_BEHAVIORAL of FA_692 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136820, net136821, net152734, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136820);
   U4 : XOR2_X1 port map( A => A, B => B, Z => net152734);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => net152734, ZN => net136821);
   U6 : NAND2_X1 port map( A1 => net136821, A2 => net136820, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_691 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_691;

architecture SYN_BEHAVIORAL of FA_691 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_690 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_690;

architecture SYN_BEHAVIORAL of FA_690 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_689 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_689;

architecture SYN_BEHAVIORAL of FA_689 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_688 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_688;

architecture SYN_BEHAVIORAL of FA_688 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_687 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_687;

architecture SYN_BEHAVIORAL of FA_687 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_686 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_686;

architecture SYN_BEHAVIORAL of FA_686 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_685 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_685;

architecture SYN_BEHAVIORAL of FA_685 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_684 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_684;

architecture SYN_BEHAVIORAL of FA_684 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_683 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_683;

architecture SYN_BEHAVIORAL of FA_683 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_682 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_682;

architecture SYN_BEHAVIORAL of FA_682 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_681 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_681;

architecture SYN_BEHAVIORAL of FA_681 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_680 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_680;

architecture SYN_BEHAVIORAL of FA_680 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_679 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_679;

architecture SYN_BEHAVIORAL of FA_679 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_678 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_678;

architecture SYN_BEHAVIORAL of FA_678 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_677 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_677;

architecture SYN_BEHAVIORAL of FA_677 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_676 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_676;

architecture SYN_BEHAVIORAL of FA_676 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_675 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_675;

architecture SYN_BEHAVIORAL of FA_675 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_674 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_674;

architecture SYN_BEHAVIORAL of FA_674 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_673 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_673;

architecture SYN_BEHAVIORAL of FA_673 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_672 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_672;

architecture SYN_BEHAVIORAL of FA_672 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_671 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_671;

architecture SYN_BEHAVIORAL of FA_671 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_670 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_670;

architecture SYN_BEHAVIORAL of FA_670 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_669 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_669;

architecture SYN_BEHAVIORAL of FA_669 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_668 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_668;

architecture SYN_BEHAVIORAL of FA_668 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_667 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_667;

architecture SYN_BEHAVIORAL of FA_667 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_666 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_666;

architecture SYN_BEHAVIORAL of FA_666 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_665 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_665;

architecture SYN_BEHAVIORAL of FA_665 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_664 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_664;

architecture SYN_BEHAVIORAL of FA_664 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_663 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_663;

architecture SYN_BEHAVIORAL of FA_663 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_662 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_662;

architecture SYN_BEHAVIORAL of FA_662 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_661 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_661;

architecture SYN_BEHAVIORAL of FA_661 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_660 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_660;

architecture SYN_BEHAVIORAL of FA_660 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_659 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_659;

architecture SYN_BEHAVIORAL of FA_659 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136687, net136688, net136689, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net136689);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => net136687);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136688);
   U5 : NAND2_X1 port map( A1 => net136689, A2 => net136688, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => net136687, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_658 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_658;

architecture SYN_BEHAVIORAL of FA_658 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136684, net136685, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net136685);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136684);
   U6 : NAND2_X1 port map( A1 => net136685, A2 => net136684, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_657 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_657;

architecture SYN_BEHAVIORAL of FA_657 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_656 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_656;

architecture SYN_BEHAVIORAL of FA_656 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_655 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_655;

architecture SYN_BEHAVIORAL of FA_655 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_654 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_654;

architecture SYN_BEHAVIORAL of FA_654 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_653 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_653;

architecture SYN_BEHAVIORAL of FA_653 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136664, n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : NAND2_X1 port map( A1 => n5, A2 => net136664, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136664);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U6 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_652 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_652;

architecture SYN_BEHAVIORAL of FA_652 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136660, net136661, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net136661);
   U5 : XNOR2_X1 port map( A => n5, B => B, ZN => n4);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net136660);
   U7 : NAND2_X1 port map( A1 => net136661, A2 => net136660, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_651 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_651;

architecture SYN_BEHAVIORAL of FA_651 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_650 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_650;

architecture SYN_BEHAVIORAL of FA_650 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_649 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_649;

architecture SYN_BEHAVIORAL of FA_649 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_648 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_648;

architecture SYN_BEHAVIORAL of FA_648 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_647 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_647;

architecture SYN_BEHAVIORAL of FA_647 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_646 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_646;

architecture SYN_BEHAVIORAL of FA_646 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_645 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_645;

architecture SYN_BEHAVIORAL of FA_645 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_644 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_644;

architecture SYN_BEHAVIORAL of FA_644 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_643 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_643;

architecture SYN_BEHAVIORAL of FA_643 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_642 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_642;

architecture SYN_BEHAVIORAL of FA_642 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U4 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => Ci, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_641 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_641;

architecture SYN_BEHAVIORAL of FA_641 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_640 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_640;

architecture SYN_BEHAVIORAL of FA_640 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_639 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_639;

architecture SYN_BEHAVIORAL of FA_639 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_638 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_638;

architecture SYN_BEHAVIORAL of FA_638 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_637 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_637;

architecture SYN_BEHAVIORAL of FA_637 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_636 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_636;

architecture SYN_BEHAVIORAL of FA_636 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_635 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_635;

architecture SYN_BEHAVIORAL of FA_635 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_634 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_634;

architecture SYN_BEHAVIORAL of FA_634 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_633 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_633;

architecture SYN_BEHAVIORAL of FA_633 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_632 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_632;

architecture SYN_BEHAVIORAL of FA_632 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_631 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_631;

architecture SYN_BEHAVIORAL of FA_631 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_630 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_630;

architecture SYN_BEHAVIORAL of FA_630 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136572, net136573, net149086, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U3 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => net136572);
   U4 : XOR2_X1 port map( A => B, B => A, Z => net149086);
   U5 : CLKBUF_X1 port map( A => B, Z => n4);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => net149086, ZN => net136573);
   U7 : NAND2_X1 port map( A1 => net136573, A2 => net136572, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_629 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_629;

architecture SYN_BEHAVIORAL of FA_629 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_628 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_628;

architecture SYN_BEHAVIORAL of FA_628 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136564, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : NAND2_X1 port map( A1 => net136564, A2 => n5, ZN => Co);
   U3 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n5);
   U4 : NAND2_X1 port map( A1 => A, A2 => n6, ZN => net136564);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_627 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_627;

architecture SYN_BEHAVIORAL of FA_627 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136560, net136561, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U3 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => net136561);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136560);
   U6 : NAND2_X1 port map( A1 => net136560, A2 => net136561, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_626 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_626;

architecture SYN_BEHAVIORAL of FA_626 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_625 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_625;

architecture SYN_BEHAVIORAL of FA_625 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_624 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_624;

architecture SYN_BEHAVIORAL of FA_624 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_623 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_623;

architecture SYN_BEHAVIORAL of FA_623 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_622 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_622;

architecture SYN_BEHAVIORAL of FA_622 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_621 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_621;

architecture SYN_BEHAVIORAL of FA_621 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n5, A2 => Ci, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => n8, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_620 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_620;

architecture SYN_BEHAVIORAL of FA_620 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_619 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_619;

architecture SYN_BEHAVIORAL of FA_619 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_618 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_618;

architecture SYN_BEHAVIORAL of FA_618 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_617 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_617;

architecture SYN_BEHAVIORAL of FA_617 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_616 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_616;

architecture SYN_BEHAVIORAL of FA_616 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_615 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_615;

architecture SYN_BEHAVIORAL of FA_615 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_614 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_614;

architecture SYN_BEHAVIORAL of FA_614 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_613 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_613;

architecture SYN_BEHAVIORAL of FA_613 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_612 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_612;

architecture SYN_BEHAVIORAL of FA_612 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_611 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_611;

architecture SYN_BEHAVIORAL of FA_611 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_610 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_610;

architecture SYN_BEHAVIORAL of FA_610 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_609 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_609;

architecture SYN_BEHAVIORAL of FA_609 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_608 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_608;

architecture SYN_BEHAVIORAL of FA_608 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_607 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_607;

architecture SYN_BEHAVIORAL of FA_607 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_606 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_606;

architecture SYN_BEHAVIORAL of FA_606 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_605 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_605;

architecture SYN_BEHAVIORAL of FA_605 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_604 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_604;

architecture SYN_BEHAVIORAL of FA_604 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_603 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_603;

architecture SYN_BEHAVIORAL of FA_603 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_602 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_602;

architecture SYN_BEHAVIORAL of FA_602 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_601 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_601;

architecture SYN_BEHAVIORAL of FA_601 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_600 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_600;

architecture SYN_BEHAVIORAL of FA_600 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_599 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_599;

architecture SYN_BEHAVIORAL of FA_599 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_598 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_598;

architecture SYN_BEHAVIORAL of FA_598 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_597 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_597;

architecture SYN_BEHAVIORAL of FA_597 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_596 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_596;

architecture SYN_BEHAVIORAL of FA_596 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_595 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_595;

architecture SYN_BEHAVIORAL of FA_595 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_594 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_594;

architecture SYN_BEHAVIORAL of FA_594 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136427, net136428, net136429, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net136429);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => net136427);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136428);
   U5 : NAND2_X1 port map( A1 => net136429, A2 => net136428, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => net136427, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_593 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_593;

architecture SYN_BEHAVIORAL of FA_593 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136424, net136425, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net136425);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136424);
   U6 : NAND2_X1 port map( A1 => net136425, A2 => net136424, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_592 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_592;

architecture SYN_BEHAVIORAL of FA_592 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_591 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_591;

architecture SYN_BEHAVIORAL of FA_591 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_590 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_590;

architecture SYN_BEHAVIORAL of FA_590 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_589 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_589;

architecture SYN_BEHAVIORAL of FA_589 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_588 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_588;

architecture SYN_BEHAVIORAL of FA_588 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136404, net136405, net148805, n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => net148805, ZN => net136405);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136404);
   U6 : XNOR2_X1 port map( A => B, B => n4, ZN => net148805);
   U7 : NAND2_X1 port map( A1 => net136404, A2 => net136405, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_587 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_587;

architecture SYN_BEHAVIORAL of FA_587 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_586 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_586;

architecture SYN_BEHAVIORAL of FA_586 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_585 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_585;

architecture SYN_BEHAVIORAL of FA_585 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_584 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_584;

architecture SYN_BEHAVIORAL of FA_584 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_583 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_583;

architecture SYN_BEHAVIORAL of FA_583 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_582 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_582;

architecture SYN_BEHAVIORAL of FA_582 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_581 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_581;

architecture SYN_BEHAVIORAL of FA_581 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_580 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_580;

architecture SYN_BEHAVIORAL of FA_580 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_579 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_579;

architecture SYN_BEHAVIORAL of FA_579 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_578 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_578;

architecture SYN_BEHAVIORAL of FA_578 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : INV_X1 port map( A => A, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_577 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_577;

architecture SYN_BEHAVIORAL of FA_577 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_576 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_576;

architecture SYN_BEHAVIORAL of FA_576 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_575 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_575;

architecture SYN_BEHAVIORAL of FA_575 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_574 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_574;

architecture SYN_BEHAVIORAL of FA_574 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_573 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_573;

architecture SYN_BEHAVIORAL of FA_573 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_572 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_572;

architecture SYN_BEHAVIORAL of FA_572 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_571 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_571;

architecture SYN_BEHAVIORAL of FA_571 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_570 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_570;

architecture SYN_BEHAVIORAL of FA_570 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_569 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_569;

architecture SYN_BEHAVIORAL of FA_569 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : CLKBUF_X1 port map( A => B, Z => n5);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => n5, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_568 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_568;

architecture SYN_BEHAVIORAL of FA_568 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_567 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_567;

architecture SYN_BEHAVIORAL of FA_567 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_566 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_566;

architecture SYN_BEHAVIORAL of FA_566 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136317, net136316, net136315, n3, n4 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net136317);
   U3 : NAND2_X1 port map( A1 => net136316, A2 => net136317, ZN => Co);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => net136315, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => net136315);
   U7 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => net136316);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_565 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_565;

architecture SYN_BEHAVIORAL of FA_565 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136312, net136313, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => net136313);
   U5 : XOR2_X1 port map( A => A, B => B, Z => n5);
   U6 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => net136312);
   U7 : NAND2_X1 port map( A1 => net136312, A2 => net136313, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_564 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_564;

architecture SYN_BEHAVIORAL of FA_564 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_563 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_563;

architecture SYN_BEHAVIORAL of FA_563 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136304, net136305, net149729, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net136304);
   U4 : XOR2_X1 port map( A => A, B => B, Z => net149729);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => net149729, ZN => net136305);
   U6 : NAND2_X1 port map( A1 => net136304, A2 => net136305, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_562 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_562;

architecture SYN_BEHAVIORAL of FA_562 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_561 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_561;

architecture SYN_BEHAVIORAL of FA_561 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_560 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_560;

architecture SYN_BEHAVIORAL of FA_560 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_559 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_559;

architecture SYN_BEHAVIORAL of FA_559 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_558 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_558;

architecture SYN_BEHAVIORAL of FA_558 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_557 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_557;

architecture SYN_BEHAVIORAL of FA_557 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_556 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_556;

architecture SYN_BEHAVIORAL of FA_556 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_555 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_555;

architecture SYN_BEHAVIORAL of FA_555 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_554 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_554;

architecture SYN_BEHAVIORAL of FA_554 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_553 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_553;

architecture SYN_BEHAVIORAL of FA_553 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_552 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_552;

architecture SYN_BEHAVIORAL of FA_552 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_551 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_551;

architecture SYN_BEHAVIORAL of FA_551 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_550 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_550;

architecture SYN_BEHAVIORAL of FA_550 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_549 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_549;

architecture SYN_BEHAVIORAL of FA_549 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_548 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_548;

architecture SYN_BEHAVIORAL of FA_548 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_547 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_547;

architecture SYN_BEHAVIORAL of FA_547 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_546 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_546;

architecture SYN_BEHAVIORAL of FA_546 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_545 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_545;

architecture SYN_BEHAVIORAL of FA_545 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_544 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_544;

architecture SYN_BEHAVIORAL of FA_544 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_543 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_543;

architecture SYN_BEHAVIORAL of FA_543 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_542 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_542;

architecture SYN_BEHAVIORAL of FA_542 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_541 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_541;

architecture SYN_BEHAVIORAL of FA_541 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_540 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_540;

architecture SYN_BEHAVIORAL of FA_540 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_539 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_539;

architecture SYN_BEHAVIORAL of FA_539 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_538 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_538;

architecture SYN_BEHAVIORAL of FA_538 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_537 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_537;

architecture SYN_BEHAVIORAL of FA_537 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_536 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_536;

architecture SYN_BEHAVIORAL of FA_536 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_535 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_535;

architecture SYN_BEHAVIORAL of FA_535 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_534 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_534;

architecture SYN_BEHAVIORAL of FA_534 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_533 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_533;

architecture SYN_BEHAVIORAL of FA_533 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_532 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_532;

architecture SYN_BEHAVIORAL of FA_532 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_531 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_531;

architecture SYN_BEHAVIORAL of FA_531 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_530 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_530;

architecture SYN_BEHAVIORAL of FA_530 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_529 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_529;

architecture SYN_BEHAVIORAL of FA_529 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136167, net136168, net136169, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net136169);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => net136167);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net136168);
   U5 : NAND2_X1 port map( A1 => net136169, A2 => net136168, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => net136167, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_528 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_528;

architecture SYN_BEHAVIORAL of FA_528 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136164, net136165, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net136165);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net136164);
   U6 : NAND2_X1 port map( A1 => net136165, A2 => net136164, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_527 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_527;

architecture SYN_BEHAVIORAL of FA_527 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_526 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_526;

architecture SYN_BEHAVIORAL of FA_526 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_525 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_525;

architecture SYN_BEHAVIORAL of FA_525 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_524 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_524;

architecture SYN_BEHAVIORAL of FA_524 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136149, net136148, net136147, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => net136149, A2 => net136148, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net136149);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net136148);
   U5 : XNOR2_X1 port map( A => Ci, B => net136147, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => net136147);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_523 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_523;

architecture SYN_BEHAVIORAL of FA_523 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_522 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_522;

architecture SYN_BEHAVIORAL of FA_522 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_521 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_521;

architecture SYN_BEHAVIORAL of FA_521 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_520 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_520;

architecture SYN_BEHAVIORAL of FA_520 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => n6, ZN => n4);
   U3 : CLKBUF_X1 port map( A => B, Z => n6);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U5 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_519 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_519;

architecture SYN_BEHAVIORAL of FA_519 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : XNOR2_X1 port map( A => n7, B => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_518 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_518;

architecture SYN_BEHAVIORAL of FA_518 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U7 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_517 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_517;

architecture SYN_BEHAVIORAL of FA_517 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U5 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_516 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_516;

architecture SYN_BEHAVIORAL of FA_516 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_515 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_515;

architecture SYN_BEHAVIORAL of FA_515 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U5 : NAND2_X1 port map( A1 => n7, A2 => Ci, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U7 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_514 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_514;

architecture SYN_BEHAVIORAL of FA_514 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_513 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_513;

architecture SYN_BEHAVIORAL of FA_513 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U7 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_512 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_512;

architecture SYN_BEHAVIORAL of FA_512 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => n6, ZN => n4);
   U3 : CLKBUF_X1 port map( A => B, Z => n6);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U5 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_511 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_511;

architecture SYN_BEHAVIORAL of FA_511 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n5);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n6, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_510 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_510;

architecture SYN_BEHAVIORAL of FA_510 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_509 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_509;

architecture SYN_BEHAVIORAL of FA_509 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136088, net136089, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => net136089);
   U5 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U6 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => net136088);
   U7 : NAND2_X1 port map( A1 => net136088, A2 => net136089, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_508 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_508;

architecture SYN_BEHAVIORAL of FA_508 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_507 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_507;

architecture SYN_BEHAVIORAL of FA_507 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_506 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_506;

architecture SYN_BEHAVIORAL of FA_506 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_505 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_505;

architecture SYN_BEHAVIORAL of FA_505 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_504 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_504;

architecture SYN_BEHAVIORAL of FA_504 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_503 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_503;

architecture SYN_BEHAVIORAL of FA_503 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_502 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_502;

architecture SYN_BEHAVIORAL of FA_502 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_501 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_501;

architecture SYN_BEHAVIORAL of FA_501 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136057, net136056, net136055, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net136057);
   U2 : NAND2_X1 port map( A1 => net136056, A2 => net136057, ZN => Co);
   U3 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U4 : XNOR2_X1 port map( A => Ci, B => net136055, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => net136055);
   U6 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => net136056);
   U7 : CLKBUF_X1 port map( A => B, Z => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_500 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_500;

architecture SYN_BEHAVIORAL of FA_500 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net136052, net136053, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net136053);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net136052);
   U5 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U6 : NAND2_X1 port map( A1 => net136052, A2 => net136053, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_499 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_499;

architecture SYN_BEHAVIORAL of FA_499 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net136048, net136049, net149575, n3, n4 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U4 : XOR2_X1 port map( A => A, B => B, Z => net149575);
   U5 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => net136048);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => net149575, ZN => net136049);
   U7 : NAND2_X1 port map( A1 => net136048, A2 => net136049, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_498 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_498;

architecture SYN_BEHAVIORAL of FA_498 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_497 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_497;

architecture SYN_BEHAVIORAL of FA_497 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n7, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_496 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_496;

architecture SYN_BEHAVIORAL of FA_496 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_495 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_495;

architecture SYN_BEHAVIORAL of FA_495 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_494 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_494;

architecture SYN_BEHAVIORAL of FA_494 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_493 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_493;

architecture SYN_BEHAVIORAL of FA_493 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_492 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_492;

architecture SYN_BEHAVIORAL of FA_492 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_491 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_491;

architecture SYN_BEHAVIORAL of FA_491 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_490 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_490;

architecture SYN_BEHAVIORAL of FA_490 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_489 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_489;

architecture SYN_BEHAVIORAL of FA_489 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_488 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_488;

architecture SYN_BEHAVIORAL of FA_488 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_487 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_487;

architecture SYN_BEHAVIORAL of FA_487 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_486 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_486;

architecture SYN_BEHAVIORAL of FA_486 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_485 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_485;

architecture SYN_BEHAVIORAL of FA_485 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_484 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_484;

architecture SYN_BEHAVIORAL of FA_484 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_483 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_483;

architecture SYN_BEHAVIORAL of FA_483 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_482 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_482;

architecture SYN_BEHAVIORAL of FA_482 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_481 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_481;

architecture SYN_BEHAVIORAL of FA_481 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_480 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_480;

architecture SYN_BEHAVIORAL of FA_480 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_479 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_479;

architecture SYN_BEHAVIORAL of FA_479 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_478 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_478;

architecture SYN_BEHAVIORAL of FA_478 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_477 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_477;

architecture SYN_BEHAVIORAL of FA_477 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_476 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_476;

architecture SYN_BEHAVIORAL of FA_476 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_475 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_475;

architecture SYN_BEHAVIORAL of FA_475 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_474 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_474;

architecture SYN_BEHAVIORAL of FA_474 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_473 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_473;

architecture SYN_BEHAVIORAL of FA_473 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_472 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_472;

architecture SYN_BEHAVIORAL of FA_472 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_471 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_471;

architecture SYN_BEHAVIORAL of FA_471 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_470 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_470;

architecture SYN_BEHAVIORAL of FA_470 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_469 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_469;

architecture SYN_BEHAVIORAL of FA_469 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_468 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_468;

architecture SYN_BEHAVIORAL of FA_468 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_467 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_467;

architecture SYN_BEHAVIORAL of FA_467 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_466 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_466;

architecture SYN_BEHAVIORAL of FA_466 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_465 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_465;

architecture SYN_BEHAVIORAL of FA_465 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_464 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_464;

architecture SYN_BEHAVIORAL of FA_464 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net135907, net135908, net135909, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net135909);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => net135907);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net135908);
   U5 : NAND2_X1 port map( A1 => net135909, A2 => net135908, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => net135907, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_463 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_463;

architecture SYN_BEHAVIORAL of FA_463 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135904, net135905, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net135905);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net135904);
   U6 : NAND2_X1 port map( A1 => net135904, A2 => net135905, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_462 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_462;

architecture SYN_BEHAVIORAL of FA_462 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_461 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_461;

architecture SYN_BEHAVIORAL of FA_461 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_460 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_460;

architecture SYN_BEHAVIORAL of FA_460 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_459 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_459;

architecture SYN_BEHAVIORAL of FA_459 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_458 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_458;

architecture SYN_BEHAVIORAL of FA_458 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_457 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_457;

architecture SYN_BEHAVIORAL of FA_457 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_456 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_456;

architecture SYN_BEHAVIORAL of FA_456 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_455 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_455;

architecture SYN_BEHAVIORAL of FA_455 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_454 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_454;

architecture SYN_BEHAVIORAL of FA_454 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_453 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_453;

architecture SYN_BEHAVIORAL of FA_453 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_452 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_452;

architecture SYN_BEHAVIORAL of FA_452 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_451 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_451;

architecture SYN_BEHAVIORAL of FA_451 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_450 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_450;

architecture SYN_BEHAVIORAL of FA_450 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_449 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_449;

architecture SYN_BEHAVIORAL of FA_449 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_448 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_448;

architecture SYN_BEHAVIORAL of FA_448 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_447 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_447;

architecture SYN_BEHAVIORAL of FA_447 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_446 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_446;

architecture SYN_BEHAVIORAL of FA_446 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_445 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_445;

architecture SYN_BEHAVIORAL of FA_445 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135833, net135832, net135831, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => net135833, A2 => net135832, ZN => Co);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net135832);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net135833);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => net135831);
   U6 : XNOR2_X1 port map( A => Ci, B => net135831, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_444 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_444;

architecture SYN_BEHAVIORAL of FA_444 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => n7, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_443 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_443;

architecture SYN_BEHAVIORAL of FA_443 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n5);
   U6 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_442 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_442;

architecture SYN_BEHAVIORAL of FA_442 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n8);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : NAND2_X1 port map( A1 => A, A2 => n7, ZN => n5);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n8, ZN => n6);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U8 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_441 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_441;

architecture SYN_BEHAVIORAL of FA_441 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U5 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n5);
   U7 : XNOR2_X1 port map( A => n4, B => Ci, ZN => S);
   U8 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_440 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_440;

architecture SYN_BEHAVIORAL of FA_440 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U5 : XNOR2_X1 port map( A => B, B => n8, ZN => n7);
   U6 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n5);
   U7 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U8 : XNOR2_X1 port map( A => B, B => A, ZN => n4);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_439 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_439;

architecture SYN_BEHAVIORAL of FA_439 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U3 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n7, ZN => n6);
   U5 : XOR2_X1 port map( A => B, B => A, Z => n7);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U7 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_438 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_438;

architecture SYN_BEHAVIORAL of FA_438 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net135804, net135805, n3, n4, n5 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => net135805);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => net135804);
   U6 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U7 : NAND2_X1 port map( A1 => net135805, A2 => net135804, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_437 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_437;

architecture SYN_BEHAVIORAL of FA_437 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_436 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_436;

architecture SYN_BEHAVIORAL of FA_436 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135796, net135797, net148884, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U3 : XOR2_X1 port map( A => B, B => A, Z => net148884);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net135796);
   U5 : NAND2_X1 port map( A1 => net148884, A2 => Ci, ZN => net135797);
   U6 : NAND2_X1 port map( A1 => net135797, A2 => net135796, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_435 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_435;

architecture SYN_BEHAVIORAL of FA_435 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135792, net135793, net149073, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => net149073);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n5);
   U5 : XNOR2_X1 port map( A => n5, B => Ci, ZN => S);
   U6 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => net135792);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => net149073, ZN => net135793);
   U8 : NAND2_X1 port map( A1 => net135792, A2 => net135793, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_434 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_434;

architecture SYN_BEHAVIORAL of FA_434 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_433 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_433;

architecture SYN_BEHAVIORAL of FA_433 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_432 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_432;

architecture SYN_BEHAVIORAL of FA_432 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_431 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_431;

architecture SYN_BEHAVIORAL of FA_431 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_430 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_430;

architecture SYN_BEHAVIORAL of FA_430 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_429 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_429;

architecture SYN_BEHAVIORAL of FA_429 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_428 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_428;

architecture SYN_BEHAVIORAL of FA_428 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_427 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_427;

architecture SYN_BEHAVIORAL of FA_427 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_426 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_426;

architecture SYN_BEHAVIORAL of FA_426 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_425 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_425;

architecture SYN_BEHAVIORAL of FA_425 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_424 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_424;

architecture SYN_BEHAVIORAL of FA_424 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_423 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_423;

architecture SYN_BEHAVIORAL of FA_423 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_422 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_422;

architecture SYN_BEHAVIORAL of FA_422 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_421 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_421;

architecture SYN_BEHAVIORAL of FA_421 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_420 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_420;

architecture SYN_BEHAVIORAL of FA_420 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_419 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_419;

architecture SYN_BEHAVIORAL of FA_419 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_418 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_418;

architecture SYN_BEHAVIORAL of FA_418 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_417 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_417;

architecture SYN_BEHAVIORAL of FA_417 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_416 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_416;

architecture SYN_BEHAVIORAL of FA_416 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_415 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_415;

architecture SYN_BEHAVIORAL of FA_415 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_414 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_414;

architecture SYN_BEHAVIORAL of FA_414 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_413 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_413;

architecture SYN_BEHAVIORAL of FA_413 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_412 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_412;

architecture SYN_BEHAVIORAL of FA_412 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_411 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_411;

architecture SYN_BEHAVIORAL of FA_411 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_410 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_410;

architecture SYN_BEHAVIORAL of FA_410 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_409 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_409;

architecture SYN_BEHAVIORAL of FA_409 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_408 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_408;

architecture SYN_BEHAVIORAL of FA_408 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_407 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_407;

architecture SYN_BEHAVIORAL of FA_407 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_406 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_406;

architecture SYN_BEHAVIORAL of FA_406 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_405 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_405;

architecture SYN_BEHAVIORAL of FA_405 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_404 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_404;

architecture SYN_BEHAVIORAL of FA_404 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_403 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_403;

architecture SYN_BEHAVIORAL of FA_403 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_402 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_402;

architecture SYN_BEHAVIORAL of FA_402 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_401 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_401;

architecture SYN_BEHAVIORAL of FA_401 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_400 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_400;

architecture SYN_BEHAVIORAL of FA_400 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_399 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_399;

architecture SYN_BEHAVIORAL of FA_399 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net135647, net135648, net135649, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net135649);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => net135647);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net135648);
   U5 : NAND2_X1 port map( A1 => net135649, A2 => net135648, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => net135647, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_398 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_398;

architecture SYN_BEHAVIORAL of FA_398 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_397 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_397;

architecture SYN_BEHAVIORAL of FA_397 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => n7, B => B, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_396 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_396;

architecture SYN_BEHAVIORAL of FA_396 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_395 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_395;

architecture SYN_BEHAVIORAL of FA_395 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135632, net135633, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => net135633);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net135632);
   U7 : NAND2_X1 port map( A1 => net135633, A2 => net135632, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_394 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_394;

architecture SYN_BEHAVIORAL of FA_394 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_393 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_393;

architecture SYN_BEHAVIORAL of FA_393 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_392 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_392;

architecture SYN_BEHAVIORAL of FA_392 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_391 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_391;

architecture SYN_BEHAVIORAL of FA_391 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_390 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_390;

architecture SYN_BEHAVIORAL of FA_390 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_389 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_389;

architecture SYN_BEHAVIORAL of FA_389 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_388 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_388;

architecture SYN_BEHAVIORAL of FA_388 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_387 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_387;

architecture SYN_BEHAVIORAL of FA_387 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_386 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_386;

architecture SYN_BEHAVIORAL of FA_386 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_385 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_385;

architecture SYN_BEHAVIORAL of FA_385 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_384 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_384;

architecture SYN_BEHAVIORAL of FA_384 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_383 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_383;

architecture SYN_BEHAVIORAL of FA_383 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_382 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_382;

architecture SYN_BEHAVIORAL of FA_382 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_381 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_381;

architecture SYN_BEHAVIORAL of FA_381 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_380 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_380;

architecture SYN_BEHAVIORAL of FA_380 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_379 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_379;

architecture SYN_BEHAVIORAL of FA_379 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_378 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_378;

architecture SYN_BEHAVIORAL of FA_378 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_377 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_377;

architecture SYN_BEHAVIORAL of FA_377 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_376 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_376;

architecture SYN_BEHAVIORAL of FA_376 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_375 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_375;

architecture SYN_BEHAVIORAL of FA_375 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_374 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_374;

architecture SYN_BEHAVIORAL of FA_374 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135548, net135549, net148779, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => net148779);
   U6 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => net135548);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => net148779, ZN => net135549);
   U8 : NAND2_X1 port map( A1 => net135549, A2 => net135548, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_373 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_373;

architecture SYN_BEHAVIORAL of FA_373 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_372 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_372;

architecture SYN_BEHAVIORAL of FA_372 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net135541, net135540, net135539, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => net135541);
   U2 : NAND2_X1 port map( A1 => net135541, A2 => net135540, ZN => Co);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U4 : XNOR2_X1 port map( A => Ci, B => net135539, ZN => S);
   U5 : CLKBUF_X1 port map( A => B, Z => n4);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => net135539);
   U7 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => net135540);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_371 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_371;

architecture SYN_BEHAVIORAL of FA_371 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135536, net135537, net149082, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => net149082, ZN => net135537);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net135536);
   U5 : XOR2_X1 port map( A => B, B => A, Z => net149082);
   U6 : NAND2_X1 port map( A1 => net135537, A2 => net135536, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_370 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_370;

architecture SYN_BEHAVIORAL of FA_370 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_369 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_369;

architecture SYN_BEHAVIORAL of FA_369 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n7, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_368 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_368;

architecture SYN_BEHAVIORAL of FA_368 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_367 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_367;

architecture SYN_BEHAVIORAL of FA_367 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_366 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_366;

architecture SYN_BEHAVIORAL of FA_366 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_365 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_365;

architecture SYN_BEHAVIORAL of FA_365 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_364 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_364;

architecture SYN_BEHAVIORAL of FA_364 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_363 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_363;

architecture SYN_BEHAVIORAL of FA_363 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_362 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_362;

architecture SYN_BEHAVIORAL of FA_362 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_361 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_361;

architecture SYN_BEHAVIORAL of FA_361 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_360 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_360;

architecture SYN_BEHAVIORAL of FA_360 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_359 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_359;

architecture SYN_BEHAVIORAL of FA_359 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_358 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_358;

architecture SYN_BEHAVIORAL of FA_358 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_357 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_357;

architecture SYN_BEHAVIORAL of FA_357 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_356 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_356;

architecture SYN_BEHAVIORAL of FA_356 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_355 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_355;

architecture SYN_BEHAVIORAL of FA_355 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_354 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_354;

architecture SYN_BEHAVIORAL of FA_354 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_353 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_353;

architecture SYN_BEHAVIORAL of FA_353 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_352 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_352;

architecture SYN_BEHAVIORAL of FA_352 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_351 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_351;

architecture SYN_BEHAVIORAL of FA_351 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_350 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_350;

architecture SYN_BEHAVIORAL of FA_350 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_349 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_349;

architecture SYN_BEHAVIORAL of FA_349 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_348 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_348;

architecture SYN_BEHAVIORAL of FA_348 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_347 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_347;

architecture SYN_BEHAVIORAL of FA_347 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_346 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_346;

architecture SYN_BEHAVIORAL of FA_346 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_345 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_345;

architecture SYN_BEHAVIORAL of FA_345 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_344 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_344;

architecture SYN_BEHAVIORAL of FA_344 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_343 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_343;

architecture SYN_BEHAVIORAL of FA_343 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_342 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_342;

architecture SYN_BEHAVIORAL of FA_342 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_341 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_341;

architecture SYN_BEHAVIORAL of FA_341 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_340 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_340;

architecture SYN_BEHAVIORAL of FA_340 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_339 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_339;

architecture SYN_BEHAVIORAL of FA_339 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_338 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_338;

architecture SYN_BEHAVIORAL of FA_338 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_337 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_337;

architecture SYN_BEHAVIORAL of FA_337 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_336 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_336;

architecture SYN_BEHAVIORAL of FA_336 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_335 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_335;

architecture SYN_BEHAVIORAL of FA_335 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_334 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_334;

architecture SYN_BEHAVIORAL of FA_334 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_333 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_333;

architecture SYN_BEHAVIORAL of FA_333 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_332 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_332;

architecture SYN_BEHAVIORAL of FA_332 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_331 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_331;

architecture SYN_BEHAVIORAL of FA_331 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135376, net135377, net148753, n3 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net135376);
   U4 : XOR2_X1 port map( A => A, B => B, Z => net148753);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => net148753, ZN => net135377);
   U6 : NAND2_X1 port map( A1 => net135377, A2 => net135376, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_330 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_330;

architecture SYN_BEHAVIORAL of FA_330 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_329 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_329;

architecture SYN_BEHAVIORAL of FA_329 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_328 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_328;

architecture SYN_BEHAVIORAL of FA_328 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_327 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_327;

architecture SYN_BEHAVIORAL of FA_327 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_326 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_326;

architecture SYN_BEHAVIORAL of FA_326 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_325 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_325;

architecture SYN_BEHAVIORAL of FA_325 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_324 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_324;

architecture SYN_BEHAVIORAL of FA_324 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_323 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_323;

architecture SYN_BEHAVIORAL of FA_323 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_322 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_322;

architecture SYN_BEHAVIORAL of FA_322 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_321 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_321;

architecture SYN_BEHAVIORAL of FA_321 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_320 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_320;

architecture SYN_BEHAVIORAL of FA_320 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_319 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_319;

architecture SYN_BEHAVIORAL of FA_319 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_318 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_318;

architecture SYN_BEHAVIORAL of FA_318 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_317 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_317;

architecture SYN_BEHAVIORAL of FA_317 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_316 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_316;

architecture SYN_BEHAVIORAL of FA_316 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_315 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_315;

architecture SYN_BEHAVIORAL of FA_315 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_314 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_314;

architecture SYN_BEHAVIORAL of FA_314 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n5);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_313 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_313;

architecture SYN_BEHAVIORAL of FA_313 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_312 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_312;

architecture SYN_BEHAVIORAL of FA_312 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_311 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_311;

architecture SYN_BEHAVIORAL of FA_311 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_310 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_310;

architecture SYN_BEHAVIORAL of FA_310 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135293, net135292, net135291, n3 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => net135293, A2 => net135292, ZN => Co);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net135292);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net135293);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => net135291);
   U6 : XNOR2_X1 port map( A => Ci, B => net135291, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_309 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_309;

architecture SYN_BEHAVIORAL of FA_309 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n6);
   U4 : NAND2_X1 port map( A1 => A, A2 => n7, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n7);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_308 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_308;

architecture SYN_BEHAVIORAL of FA_308 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n6);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U6 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_307 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_307;

architecture SYN_BEHAVIORAL of FA_307 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net135281, net135280, net135279, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net135281);
   U2 : NAND2_X1 port map( A1 => net135281, A2 => net135280, ZN => Co);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U4 : XNOR2_X1 port map( A => Ci, B => net135279, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => A, ZN => net135279);
   U6 : CLKBUF_X1 port map( A => B, Z => n4);
   U7 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => net135280);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_306 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_306;

architecture SYN_BEHAVIORAL of FA_306 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135276, net135277, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : INV_X1 port map( A => n3, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net135277);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : NAND2_X1 port map( A1 => A, A2 => n5, ZN => net135276);
   U7 : NAND2_X1 port map( A1 => net135276, A2 => net135277, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_305 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_305;

architecture SYN_BEHAVIORAL of FA_305 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n7);
   U5 : INV_X1 port map( A => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_304 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_304;

architecture SYN_BEHAVIORAL of FA_304 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_303 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_303;

architecture SYN_BEHAVIORAL of FA_303 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_302 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_302;

architecture SYN_BEHAVIORAL of FA_302 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_301 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_301;

architecture SYN_BEHAVIORAL of FA_301 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_300 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_300;

architecture SYN_BEHAVIORAL of FA_300 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_299 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_299;

architecture SYN_BEHAVIORAL of FA_299 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_298 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_298;

architecture SYN_BEHAVIORAL of FA_298 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_297 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_297;

architecture SYN_BEHAVIORAL of FA_297 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_296 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_296;

architecture SYN_BEHAVIORAL of FA_296 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_295 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_295;

architecture SYN_BEHAVIORAL of FA_295 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_294 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_294;

architecture SYN_BEHAVIORAL of FA_294 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_293 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_293;

architecture SYN_BEHAVIORAL of FA_293 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_292 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_292;

architecture SYN_BEHAVIORAL of FA_292 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_291 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_291;

architecture SYN_BEHAVIORAL of FA_291 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_290 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_290;

architecture SYN_BEHAVIORAL of FA_290 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_289 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_289;

architecture SYN_BEHAVIORAL of FA_289 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_288 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_288;

architecture SYN_BEHAVIORAL of FA_288 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_287 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_287;

architecture SYN_BEHAVIORAL of FA_287 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_286 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_286;

architecture SYN_BEHAVIORAL of FA_286 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_285 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_285;

architecture SYN_BEHAVIORAL of FA_285 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_284 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_284;

architecture SYN_BEHAVIORAL of FA_284 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_283 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_283;

architecture SYN_BEHAVIORAL of FA_283 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_282 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_282;

architecture SYN_BEHAVIORAL of FA_282 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_281 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_281;

architecture SYN_BEHAVIORAL of FA_281 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_280 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_280;

architecture SYN_BEHAVIORAL of FA_280 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_279 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_279;

architecture SYN_BEHAVIORAL of FA_279 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_278 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_278;

architecture SYN_BEHAVIORAL of FA_278 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_277 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_277;

architecture SYN_BEHAVIORAL of FA_277 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_276 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_276;

architecture SYN_BEHAVIORAL of FA_276 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_275 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_275;

architecture SYN_BEHAVIORAL of FA_275 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_274 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_274;

architecture SYN_BEHAVIORAL of FA_274 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_273 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_273;

architecture SYN_BEHAVIORAL of FA_273 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_272 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_272;

architecture SYN_BEHAVIORAL of FA_272 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_271 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_271;

architecture SYN_BEHAVIORAL of FA_271 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_270 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_270;

architecture SYN_BEHAVIORAL of FA_270 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_269 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_269;

architecture SYN_BEHAVIORAL of FA_269 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_268 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_268;

architecture SYN_BEHAVIORAL of FA_268 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_267 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_267;

architecture SYN_BEHAVIORAL of FA_267 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135120, net135121, net147396, n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => net147396);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net135120);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => net147396, ZN => net135121);
   U7 : NAND2_X1 port map( A1 => net135121, A2 => net135120, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_266 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_266;

architecture SYN_BEHAVIORAL of FA_266 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_265 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_265;

architecture SYN_BEHAVIORAL of FA_265 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => n4, A2 => Ci, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_264 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_264;

architecture SYN_BEHAVIORAL of FA_264 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_263 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_263;

architecture SYN_BEHAVIORAL of FA_263 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_262 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_262;

architecture SYN_BEHAVIORAL of FA_262 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_261 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_261;

architecture SYN_BEHAVIORAL of FA_261 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_260 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_260;

architecture SYN_BEHAVIORAL of FA_260 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_259 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_259;

architecture SYN_BEHAVIORAL of FA_259 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_258 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_258;

architecture SYN_BEHAVIORAL of FA_258 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_257 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_257;

architecture SYN_BEHAVIORAL of FA_257 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_256 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_256;

architecture SYN_BEHAVIORAL of FA_256 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_255 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_255;

architecture SYN_BEHAVIORAL of FA_255 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_254 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_254;

architecture SYN_BEHAVIORAL of FA_254 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_253 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_253;

architecture SYN_BEHAVIORAL of FA_253 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_252 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_252;

architecture SYN_BEHAVIORAL of FA_252 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_251 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_251;

architecture SYN_BEHAVIORAL of FA_251 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_250 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_250;

architecture SYN_BEHAVIORAL of FA_250 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_249 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_249;

architecture SYN_BEHAVIORAL of FA_249 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_248 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_248;

architecture SYN_BEHAVIORAL of FA_248 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_247 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_247;

architecture SYN_BEHAVIORAL of FA_247 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_246 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_246;

architecture SYN_BEHAVIORAL of FA_246 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_245 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_245;

architecture SYN_BEHAVIORAL of FA_245 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_244 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_244;

architecture SYN_BEHAVIORAL of FA_244 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_243 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_243;

architecture SYN_BEHAVIORAL of FA_243 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135024, net135025, net148778, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : CLKBUF_X1 port map( A => B, Z => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U5 : XNOR2_X1 port map( A => B, B => n5, ZN => net148778);
   U6 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => net135024);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => net148778, ZN => net135025);
   U8 : NAND2_X1 port map( A1 => net135024, A2 => net135025, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_242 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_242;

architecture SYN_BEHAVIORAL of FA_242 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net135020, net135021, net148887, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XOR2_X1 port map( A => B, B => A, Z => net148887);
   U5 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => net135020);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => net148887, ZN => net135021);
   U7 : NAND2_X1 port map( A1 => net135020, A2 => net135021, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_241 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_241;

architecture SYN_BEHAVIORAL of FA_241 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : CLKBUF_X1 port map( A => n9, Z => n4);
   U3 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n9);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n8);
   U6 : INV_X1 port map( A => n4, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => n7);
   U8 : NAND2_X1 port map( A1 => n8, A2 => n7, ZN => Co);
   U9 : XNOR2_X1 port map( A => n9, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_240 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_240;

architecture SYN_BEHAVIORAL of FA_240 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_239 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_239;

architecture SYN_BEHAVIORAL of FA_239 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_238 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_238;

architecture SYN_BEHAVIORAL of FA_238 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_237 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_237;

architecture SYN_BEHAVIORAL of FA_237 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_236 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_236;

architecture SYN_BEHAVIORAL of FA_236 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_235 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_235;

architecture SYN_BEHAVIORAL of FA_235 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_234 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_234;

architecture SYN_BEHAVIORAL of FA_234 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_233 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_233;

architecture SYN_BEHAVIORAL of FA_233 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_232 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_232;

architecture SYN_BEHAVIORAL of FA_232 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_231 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_231;

architecture SYN_BEHAVIORAL of FA_231 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => n6, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_230 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_230;

architecture SYN_BEHAVIORAL of FA_230 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_229 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_229;

architecture SYN_BEHAVIORAL of FA_229 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_228 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_228;

architecture SYN_BEHAVIORAL of FA_228 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_227 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_227;

architecture SYN_BEHAVIORAL of FA_227 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_226 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_226;

architecture SYN_BEHAVIORAL of FA_226 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_225 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_225;

architecture SYN_BEHAVIORAL of FA_225 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_224 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_224;

architecture SYN_BEHAVIORAL of FA_224 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n7, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_223 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_223;

architecture SYN_BEHAVIORAL of FA_223 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_222 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_222;

architecture SYN_BEHAVIORAL of FA_222 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_221 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_221;

architecture SYN_BEHAVIORAL of FA_221 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_220 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_220;

architecture SYN_BEHAVIORAL of FA_220 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_219 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_219;

architecture SYN_BEHAVIORAL of FA_219 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n7, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_218 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_218;

architecture SYN_BEHAVIORAL of FA_218 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_217 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_217;

architecture SYN_BEHAVIORAL of FA_217 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_216 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_216;

architecture SYN_BEHAVIORAL of FA_216 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_215 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_215;

architecture SYN_BEHAVIORAL of FA_215 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_214 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_214;

architecture SYN_BEHAVIORAL of FA_214 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_213 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_213;

architecture SYN_BEHAVIORAL of FA_213 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_212 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_212;

architecture SYN_BEHAVIORAL of FA_212 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_211 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_211;

architecture SYN_BEHAVIORAL of FA_211 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_210 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_210;

architecture SYN_BEHAVIORAL of FA_210 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_209 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_209;

architecture SYN_BEHAVIORAL of FA_209 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_208 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_208;

architecture SYN_BEHAVIORAL of FA_208 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_207 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_207;

architecture SYN_BEHAVIORAL of FA_207 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_206 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_206;

architecture SYN_BEHAVIORAL of FA_206 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_205 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_205;

architecture SYN_BEHAVIORAL of FA_205 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_204 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_204;

architecture SYN_BEHAVIORAL of FA_204 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_203 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_203;

architecture SYN_BEHAVIORAL of FA_203 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net134863, net134864, net134865, n3 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => net134865);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net134864);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => net134863);
   U5 : NAND2_X1 port map( A1 => net134865, A2 => net134864, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => net134863, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_202 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_202;

architecture SYN_BEHAVIORAL of FA_202 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_201 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_201;

architecture SYN_BEHAVIORAL of FA_201 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_200 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_200;

architecture SYN_BEHAVIORAL of FA_200 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_199 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_199;

architecture SYN_BEHAVIORAL of FA_199 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => n3, B => B, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_198 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_198;

architecture SYN_BEHAVIORAL of FA_198 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_197 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_197;

architecture SYN_BEHAVIORAL of FA_197 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_196 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_196;

architecture SYN_BEHAVIORAL of FA_196 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_195 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_195;

architecture SYN_BEHAVIORAL of FA_195 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_194 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_194;

architecture SYN_BEHAVIORAL of FA_194 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_193 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_193;

architecture SYN_BEHAVIORAL of FA_193 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_192 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_192;

architecture SYN_BEHAVIORAL of FA_192 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_191 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_191;

architecture SYN_BEHAVIORAL of FA_191 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_190 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_190;

architecture SYN_BEHAVIORAL of FA_190 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => n7, B => B, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_189 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_189;

architecture SYN_BEHAVIORAL of FA_189 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_188 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_188;

architecture SYN_BEHAVIORAL of FA_188 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n7);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n4);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U5 : XNOR2_X1 port map( A => B, B => n7, ZN => n6);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_187 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_187;

architecture SYN_BEHAVIORAL of FA_187 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_186 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_186;

architecture SYN_BEHAVIORAL of FA_186 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_185 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_185;

architecture SYN_BEHAVIORAL of FA_185 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_184 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_184;

architecture SYN_BEHAVIORAL of FA_184 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_183 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_183;

architecture SYN_BEHAVIORAL of FA_183 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_182 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_182;

architecture SYN_BEHAVIORAL of FA_182 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n8);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U3 : NAND2_X1 port map( A1 => n7, A2 => A, ZN => n4);
   U4 : CLKBUF_X1 port map( A => B, Z => n7);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n6, ZN => n5);
   U6 : XNOR2_X1 port map( A => B, B => n8, ZN => n6);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U8 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_181 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_181;

architecture SYN_BEHAVIORAL of FA_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net134776, net134777, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => net134777);
   U4 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n5);
   U6 : NAND2_X1 port map( A1 => A, A2 => n5, ZN => net134776);
   U7 : NAND2_X1 port map( A1 => net134777, A2 => net134776, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_180 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_180;

architecture SYN_BEHAVIORAL of FA_180 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : CLKBUF_X1 port map( A => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_179 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_179;

architecture SYN_BEHAVIORAL of FA_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net134768, net134769, net148793, n3, n4 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => n4, ZN => net148793);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => net134768);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => net148793, ZN => net134769);
   U7 : NAND2_X1 port map( A1 => net134769, A2 => net134768, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_178 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_178;

architecture SYN_BEHAVIORAL of FA_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net134764, net134765, net148581, n3, n4 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XOR2_X1 port map( A => B, B => A, Z => net148581);
   U5 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => net134764);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => net148581, ZN => net134765);
   U7 : NAND2_X1 port map( A1 => net134765, A2 => net134764, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_177 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_177;

architecture SYN_BEHAVIORAL of FA_177 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n7);
   U5 : INV_X1 port map( A => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_176 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_176;

architecture SYN_BEHAVIORAL of FA_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_175 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_175;

architecture SYN_BEHAVIORAL of FA_175 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_174 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_174;

architecture SYN_BEHAVIORAL of FA_174 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_173 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_173;

architecture SYN_BEHAVIORAL of FA_173 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_172 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_172;

architecture SYN_BEHAVIORAL of FA_172 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_171 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_171;

architecture SYN_BEHAVIORAL of FA_171 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_170 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_170;

architecture SYN_BEHAVIORAL of FA_170 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_169 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_169;

architecture SYN_BEHAVIORAL of FA_169 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_168 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_168;

architecture SYN_BEHAVIORAL of FA_168 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_167 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_167;

architecture SYN_BEHAVIORAL of FA_167 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_166 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_166;

architecture SYN_BEHAVIORAL of FA_166 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_165 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_165;

architecture SYN_BEHAVIORAL of FA_165 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_164 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_164;

architecture SYN_BEHAVIORAL of FA_164 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_163 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_163;

architecture SYN_BEHAVIORAL of FA_163 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_162 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_162;

architecture SYN_BEHAVIORAL of FA_162 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_161 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_161;

architecture SYN_BEHAVIORAL of FA_161 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_160 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_160;

architecture SYN_BEHAVIORAL of FA_160 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_159 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_159;

architecture SYN_BEHAVIORAL of FA_159 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_158 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_158;

architecture SYN_BEHAVIORAL of FA_158 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_157 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_157;

architecture SYN_BEHAVIORAL of FA_157 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_156 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_156;

architecture SYN_BEHAVIORAL of FA_156 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_155 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_155;

architecture SYN_BEHAVIORAL of FA_155 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_154 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_154;

architecture SYN_BEHAVIORAL of FA_154 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_153 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_153;

architecture SYN_BEHAVIORAL of FA_153 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_152 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_152;

architecture SYN_BEHAVIORAL of FA_152 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_151 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_151;

architecture SYN_BEHAVIORAL of FA_151 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_150 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_150;

architecture SYN_BEHAVIORAL of FA_150 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_149 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_149;

architecture SYN_BEHAVIORAL of FA_149 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_148 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_148;

architecture SYN_BEHAVIORAL of FA_148 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_147 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_147;

architecture SYN_BEHAVIORAL of FA_147 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_146 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_146;

architecture SYN_BEHAVIORAL of FA_146 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : INV_X1 port map( A => n3, ZN => n4);
   U3 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n5, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_145 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_145;

architecture SYN_BEHAVIORAL of FA_145 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_144 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_144;

architecture SYN_BEHAVIORAL of FA_144 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_143 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_143;

architecture SYN_BEHAVIORAL of FA_143 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : CLKBUF_X1 port map( A => n8, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => n3, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_142 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_142;

architecture SYN_BEHAVIORAL of FA_142 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_141 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_141;

architecture SYN_BEHAVIORAL of FA_141 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_140 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_140;

architecture SYN_BEHAVIORAL of FA_140 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_139 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_139;

architecture SYN_BEHAVIORAL of FA_139 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XOR2_X1 port map( A => A, B => B, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_138 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_138;

architecture SYN_BEHAVIORAL of FA_138 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n7, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_137 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_137;

architecture SYN_BEHAVIORAL of FA_137 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n7, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_136 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_136;

architecture SYN_BEHAVIORAL of FA_136 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U2 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_135 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_135;

architecture SYN_BEHAVIORAL of FA_135 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n7, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_134 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_134;

architecture SYN_BEHAVIORAL of FA_134 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_133 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_133;

architecture SYN_BEHAVIORAL of FA_133 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => Ci, Z => n3);
   U2 : INV_X1 port map( A => A, ZN => n4);
   U3 : XNOR2_X1 port map( A => n4, B => B, ZN => n5);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => n3, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_132 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_132;

architecture SYN_BEHAVIORAL of FA_132 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_131 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_131;

architecture SYN_BEHAVIORAL of FA_131 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_130 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_130;

architecture SYN_BEHAVIORAL of FA_130 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_129 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_129;

architecture SYN_BEHAVIORAL of FA_129 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_128 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_128;

architecture SYN_BEHAVIORAL of FA_128 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_127 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_127;

architecture SYN_BEHAVIORAL of FA_127 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_126 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_126;

architecture SYN_BEHAVIORAL of FA_126 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_125 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_125;

architecture SYN_BEHAVIORAL of FA_125 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n6);
   U3 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n5);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_124 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_124;

architecture SYN_BEHAVIORAL of FA_124 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U3 : XNOR2_X1 port map( A => n4, B => B, ZN => n3);
   U4 : INV_X1 port map( A => n3, ZN => n5);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n8);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n7);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => Co);
   U8 : XNOR2_X1 port map( A => n6, B => n5, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_123 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_123;

architecture SYN_BEHAVIORAL of FA_123 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_122 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_122;

architecture SYN_BEHAVIORAL of FA_122 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => B, Z => n3);
   U2 : CLKBUF_X1 port map( A => n3, Z => n4);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U4 : XNOR2_X1 port map( A => n3, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_121 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_121;

architecture SYN_BEHAVIORAL of FA_121 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : INV_X1 port map( A => n3, ZN => n7);
   U3 : XNOR2_X1 port map( A => B, B => n4, ZN => n3);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n7, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_120 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_120;

architecture SYN_BEHAVIORAL of FA_120 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => n3, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_119 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_119;

architecture SYN_BEHAVIORAL of FA_119 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X32
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => B, B => n3, ZN => n4);
   U2 : INV_X32 port map( A => A, ZN => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_118 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_118;

architecture SYN_BEHAVIORAL of FA_118 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_117 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_117;

architecture SYN_BEHAVIORAL of FA_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net134520, net134521, net147405, n3, n4 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U3 : XNOR2_X1 port map( A => Ci, B => n4, ZN => S);
   U4 : XOR2_X1 port map( A => B, B => A, Z => net147405);
   U5 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => net134520);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => net147405, ZN => net134521);
   U7 : NAND2_X1 port map( A1 => net134521, A2 => net134520, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_116 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_116;

architecture SYN_BEHAVIORAL of FA_116 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => B, Z => n3);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U4 : NAND2_X1 port map( A1 => n3, A2 => A, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_115 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_115;

architecture SYN_BEHAVIORAL of FA_115 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net134513, net134512, net134511, n3, n4, n5 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : NAND2_X1 port map( A1 => net134513, A2 => net134512, ZN => Co);
   U4 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => net134512);
   U5 : CLKBUF_X1 port map( A => B, Z => n4);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => net134513);
   U7 : XNOR2_X1 port map( A => B, B => A, ZN => net134511);
   U8 : XNOR2_X1 port map( A => Ci, B => net134511, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_114 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_114;

architecture SYN_BEHAVIORAL of FA_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal net134509, net134508, net134507, n3, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => net134509);
   U2 : NAND2_X1 port map( A1 => net134509, A2 => net134508, ZN => Co);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U4 : XNOR2_X1 port map( A => Ci, B => net134507, ZN => S);
   U5 : CLKBUF_X1 port map( A => B, Z => n4);
   U6 : XNOR2_X1 port map( A => B, B => A, ZN => net134507);
   U7 : NAND2_X1 port map( A1 => A, A2 => n4, ZN => net134508);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_113 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_113;

architecture SYN_BEHAVIORAL of FA_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net134504, net134506, net149730, net149817, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : CLKBUF_X1 port map( A => Ci, Z => net149817);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U4 : CLKBUF_X1 port map( A => n3, Z => net149730);
   U5 : CLKBUF_X1 port map( A => B, Z => n4);
   U6 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => net134504);
   U7 : INV_X1 port map( A => net149730, ZN => net134506);
   U8 : NAND2_X1 port map( A1 => net149817, A2 => net134506, ZN => n5);
   U9 : NAND2_X1 port map( A1 => net134504, A2 => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_112 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_112;

architecture SYN_BEHAVIORAL of FA_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => n4, B => n5, Z => S);
   U2 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n3, ZN => Co);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n4);
   U4 : INV_X1 port map( A => Ci, ZN => n5);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n3);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_111 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_111;

architecture SYN_BEHAVIORAL of FA_111 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_110 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_110;

architecture SYN_BEHAVIORAL of FA_110 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_109 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_109;

architecture SYN_BEHAVIORAL of FA_109 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_108 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_108;

architecture SYN_BEHAVIORAL of FA_108 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_107 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_107;

architecture SYN_BEHAVIORAL of FA_107 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_106 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_106;

architecture SYN_BEHAVIORAL of FA_106 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_105 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_105;

architecture SYN_BEHAVIORAL of FA_105 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_104 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_104;

architecture SYN_BEHAVIORAL of FA_104 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_103 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_103;

architecture SYN_BEHAVIORAL of FA_103 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_102 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_102;

architecture SYN_BEHAVIORAL of FA_102 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_101 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_101;

architecture SYN_BEHAVIORAL of FA_101 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_100 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_100;

architecture SYN_BEHAVIORAL of FA_100 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_99 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_99;

architecture SYN_BEHAVIORAL of FA_99 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => n3, A2 => Ci, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_98 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_98;

architecture SYN_BEHAVIORAL of FA_98 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_97 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_97;

architecture SYN_BEHAVIORAL of FA_97 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_96 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_96;

architecture SYN_BEHAVIORAL of FA_96 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n4);
   U2 : INV_X1 port map( A => n3, ZN => n7);
   U3 : XNOR2_X1 port map( A => n4, B => B, ZN => n3);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => Ci, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => n4);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => n4);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => n4);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);
   U3 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U5 : INV_X1 port map( A => n7, ZN => n4);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => n5);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U8 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => Ci, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);
   U2 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U4 : INV_X1 port map( A => n6, ZN => n3);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U6 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => n5);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U8 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U2 : XNOR2_X1 port map( A => B, B => A, ZN => n7);
   U3 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n6);
   U4 : INV_X1 port map( A => n7, ZN => n4);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n5);
   U6 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => Co);
   U7 : XNOR2_X1 port map( A => n3, B => n7, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => n5);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U8 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);
   U4 : XNOR2_X1 port map( A => A, B => B, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => n5);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U8 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => Ci, Z => n4);
   U2 : CLKBUF_X1 port map( A => n8, Z => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n7, A2 => n6, ZN => Co);
   U8 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => A, B => B, ZN => n6);
   U2 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n5);
   U3 : INV_X1 port map( A => n6, ZN => n3);
   U4 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n4);
   U5 : NAND2_X1 port map( A1 => n5, A2 => n4, ZN => Co);
   U6 : XNOR2_X1 port map( A => Ci, B => n6, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : XOR2_X1 port map( A => n6, B => n3, Z => S);
   U3 : CLKBUF_X1 port map( A => n4, Z => n3);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => Ci, Z => n6);
   U6 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n8);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n7);
   U8 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => n5);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U8 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => n4, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U4 : NAND2_X1 port map( A1 => B, A2 => A, ZN => n7);
   U5 : INV_X1 port map( A => n8, ZN => n5);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => A, B => B, Z => n3);
   U2 : INV_X1 port map( A => n3, ZN => n4);
   U3 : CLKBUF_X1 port map( A => Ci, Z => n5);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U7 : XNOR2_X1 port map( A => n5, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : CLKBUF_X1 port map( A => n8, Z => n3);
   U2 : CLKBUF_X1 port map( A => Ci, Z => n4);
   U3 : XNOR2_X1 port map( A => n4, B => n3, ZN => S);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => A, A2 => B, ZN => n7);
   U6 : INV_X1 port map( A => n8, ZN => n5);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U8 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net134264, n3, n4, n5, n6 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => Ci, Z => n5);
   U2 : XOR2_X1 port map( A => B, B => A, Z => n3);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n4);
   U4 : NAND2_X1 port map( A1 => A, A2 => B, ZN => net134264);
   U5 : NAND2_X1 port map( A1 => Ci, A2 => n3, ZN => n6);
   U6 : NAND2_X1 port map( A1 => n6, A2 => net134264, ZN => Co);
   U7 : XNOR2_X1 port map( A => n5, B => n4, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8, n9 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n5);
   U2 : INV_X1 port map( A => n4, ZN => n9);
   U3 : CLKBUF_X1 port map( A => Ci, Z => n3);
   U4 : XNOR2_X1 port map( A => B, B => n5, ZN => n4);
   U5 : CLKBUF_X1 port map( A => B, Z => n6);
   U6 : NAND2_X1 port map( A1 => A, A2 => n6, ZN => n8);
   U7 : NAND2_X1 port map( A1 => Ci, A2 => n4, ZN => n7);
   U8 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => Co);
   U9 : XNOR2_X1 port map( A => n3, B => n9, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => Ci, Z => n3);
   U2 : BUF_X1 port map( A => B, Z => n4);
   U3 : XOR2_X1 port map( A => B, B => A, Z => n5);
   U4 : XNOR2_X1 port map( A => n4, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => n3, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n3, n4, n5, n6, n7, n8 : std_logic;

begin
   
   U1 : INV_X1 port map( A => A, ZN => n3);
   U2 : XNOR2_X1 port map( A => B, B => n3, ZN => n5);
   U3 : CLKBUF_X1 port map( A => B, Z => n4);
   U4 : XNOR2_X1 port map( A => B, B => A, ZN => n8);
   U5 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => n7);
   U6 : NAND2_X1 port map( A1 => Ci, A2 => n5, ZN => n6);
   U7 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => Co);
   U8 : XNOR2_X1 port map( A => Ci, B => n8, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net134248, net134250, net148436, net148468, n3, n4, n5 : std_logic;

begin
   
   U1 : XNOR2_X1 port map( A => Ci, B => n3, ZN => S);
   U2 : CLKBUF_X1 port map( A => Ci, Z => net148436);
   U3 : XNOR2_X1 port map( A => B, B => A, ZN => n3);
   U4 : CLKBUF_X1 port map( A => n3, Z => net148468);
   U5 : CLKBUF_X1 port map( A => B, Z => n4);
   U6 : NAND2_X1 port map( A1 => n4, A2 => A, ZN => net134248);
   U7 : INV_X1 port map( A => net148468, ZN => net134250);
   U8 : NAND2_X1 port map( A1 => net148436, A2 => net134250, ZN => n5);
   U9 : NAND2_X1 port map( A1 => net134248, A2 => n5, ZN => Co);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_14 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_14;

architecture SYN_STRUCTURAL of RCA_generic_N64_14 is

   component FA_881
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_882
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_883
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_884
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_885
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_886
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_887
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_888
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_889
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_890
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_891
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_892
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_893
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_894
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_895
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_896
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_897
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_898
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_899
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_900
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_901
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_902
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_903
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_904
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_905
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_906
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_907
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_908
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_909
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_910
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_911
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_912
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_913
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_914
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_915
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_916
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_917
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_918
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_919
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_920
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_921
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_922
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_923
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_924
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_925
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_926
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_927
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_928
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_929
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_930
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_931
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_932
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_933
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_934
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_935
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_936
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_937
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_938
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_939
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_940
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_941
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_942
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_943
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_944
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_944 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_943 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_942 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_941 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_940 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_939 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_938 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_937 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_936 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_935 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_934 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_933 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_932 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_931 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_930 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_929 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_928 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_927 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_926 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_925 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_924 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_923 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_922 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_921 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_920 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_919 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_918 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_917 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_916 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_915 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_914 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_913 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_912 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_911 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_910 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_909 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_908 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_907 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_906 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_905 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_904 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_903 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_902 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_901 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_900 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_899 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_898 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_897 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_896 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_895 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_894 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_893 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_892 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_891 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_890 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_889 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_888 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_887 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_886 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_885 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_884 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_883 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_882 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_881 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_13 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_13;

architecture SYN_STRUCTURAL of RCA_generic_N64_13 is

   component FA_817
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_818
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_819
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_820
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_821
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_822
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_823
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_824
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_825
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_826
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_827
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_828
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_829
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_830
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_831
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_832
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_833
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_834
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_835
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_836
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_837
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_838
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_839
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_840
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_841
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_842
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_843
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_844
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_845
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_846
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_847
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_848
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_849
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_850
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_851
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_852
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_853
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_854
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_855
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_856
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_857
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_858
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_859
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_860
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_861
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_862
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_863
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_864
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_865
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_866
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_867
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_868
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_869
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_870
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_871
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_872
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_873
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_874
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_875
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_876
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_877
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_878
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_879
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_880
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_880 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_879 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_878 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_877 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_876 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_875 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_874 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_873 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_872 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_871 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_870 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_869 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_868 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_867 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_866 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_865 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_864 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_863 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_862 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_861 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_860 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_859 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_858 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_857 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_856 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_855 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_854 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_853 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_852 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_851 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_850 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_849 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_848 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_847 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_846 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_845 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_844 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_843 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_842 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_841 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_840 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_839 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_838 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_837 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_836 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_835 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_834 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_833 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_832 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_831 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_830 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_829 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_828 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_827 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_826 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_825 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_824 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_823 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_822 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_821 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_820 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_819 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_818 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_817 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_12 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_12;

architecture SYN_STRUCTURAL of RCA_generic_N64_12 is

   component FA_753
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_754
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_755
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_756
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_757
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_758
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_759
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_760
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_761
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_762
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_763
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_764
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_765
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_766
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_767
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_768
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_769
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_770
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_771
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_772
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_773
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_774
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_775
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_776
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_777
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_778
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_779
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_780
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_781
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_782
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_783
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_784
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_785
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_786
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_787
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_788
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_789
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_790
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_791
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_792
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_793
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_794
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_795
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_796
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_797
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_798
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_799
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_800
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_801
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_802
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_803
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_804
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_805
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_806
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_807
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_808
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_809
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_810
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_811
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_812
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_813
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_814
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_815
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_816
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_816 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_815 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_814 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_813 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_812 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_811 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_810 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_809 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_808 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_807 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_806 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_805 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_804 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_803 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_802 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_801 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_800 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_799 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_798 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_797 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_796 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_795 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_794 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_793 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_792 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_791 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_790 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_789 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_788 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_787 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_786 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_785 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_784 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_783 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_782 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_781 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_780 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_779 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_778 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_777 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_776 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_775 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_774 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_773 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_772 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_771 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_770 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_769 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_768 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_767 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_766 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_765 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_764 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_763 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_762 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_761 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_760 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_759 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_758 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_757 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_756 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_755 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_754 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_753 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_11 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_11;

architecture SYN_STRUCTURAL of RCA_generic_N64_11 is

   component FA_689
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_690
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_691
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_692
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_693
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_694
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_695
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_696
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_697
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_698
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_699
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_700
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_701
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_702
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_703
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_704
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_705
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_706
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_707
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_708
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_709
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_710
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_711
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_712
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_713
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_714
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_715
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_716
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_717
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_718
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_719
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_720
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_721
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_722
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_723
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_724
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_725
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_726
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_727
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_728
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_729
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_730
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_731
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_732
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_733
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_734
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_735
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_736
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_737
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_738
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_739
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_740
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_741
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_742
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_743
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_744
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_745
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_746
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_747
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_748
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_749
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_750
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_751
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_752
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_752 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_751 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_750 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_749 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_748 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_747 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_746 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_745 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_744 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_743 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_742 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_741 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_740 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_739 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_738 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_737 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_736 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_735 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_734 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_733 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_732 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_731 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_730 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_729 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_728 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_727 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_726 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_725 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_724 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_723 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_722 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_721 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_720 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_719 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_718 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_717 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_716 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_715 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_714 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_713 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_712 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_711 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_710 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_709 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_708 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_707 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_706 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_705 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_704 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_703 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_702 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_701 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_700 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_699 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_698 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_697 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_696 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_695 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_694 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_693 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_692 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_691 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_690 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_689 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_10 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_10;

architecture SYN_STRUCTURAL of RCA_generic_N64_10 is

   component FA_625
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_626
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_627
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_628
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_629
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_630
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_631
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_632
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_633
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_634
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_635
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_636
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_637
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_638
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_639
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_640
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_641
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_642
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_643
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_644
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_645
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_646
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_647
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_648
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_649
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_650
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_651
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_652
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_653
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_654
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_655
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_656
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_657
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_658
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_659
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_660
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_661
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_662
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_663
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_664
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_665
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_666
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_667
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_668
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_669
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_670
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_671
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_672
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_673
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_674
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_675
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_676
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_677
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_678
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_679
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_680
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_681
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_682
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_683
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_684
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_685
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_686
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_687
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_688
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_688 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_687 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_686 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_685 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_684 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_683 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_682 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_681 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_680 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_679 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_678 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_677 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_676 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_675 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_674 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_673 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_672 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_671 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_670 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_669 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_668 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_667 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_666 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_665 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_664 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_663 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_662 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_661 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_660 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_659 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_658 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_657 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_656 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_655 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_654 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_653 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_652 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_651 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_650 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_649 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_648 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_647 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_646 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_645 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_644 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_643 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_642 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_641 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_640 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_639 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_638 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_637 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_636 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_635 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_634 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_633 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_632 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_631 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_630 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_629 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_628 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_627 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_626 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_625 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_9 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_9;

architecture SYN_STRUCTURAL of RCA_generic_N64_9 is

   component FA_561
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_562
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_563
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_564
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_565
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_566
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_567
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_568
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_569
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_570
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_571
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_572
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_573
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_574
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_575
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_576
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_577
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_578
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_579
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_580
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_581
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_582
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_583
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_584
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_585
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_586
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_587
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_588
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_589
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_590
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_591
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_592
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_593
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_594
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_595
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_596
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_597
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_598
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_599
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_600
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_601
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_602
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_603
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_604
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_605
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_606
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_607
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_608
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_609
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_610
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_611
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_612
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_613
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_614
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_615
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_616
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_617
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_618
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_619
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_620
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_621
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_622
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_623
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_624
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_624 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_623 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_622 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_621 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_620 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_619 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_618 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_617 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_616 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_615 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_614 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_613 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_612 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_611 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_610 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_609 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_608 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_607 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_606 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_605 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_604 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_603 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_602 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_601 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_600 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_599 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_598 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_597 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_596 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_595 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_594 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_593 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_592 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_591 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_590 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_589 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_588 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_587 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_586 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_585 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_584 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_583 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_582 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_581 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_580 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_579 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_578 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_577 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_576 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_575 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_574 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_573 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_572 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_571 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_570 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_569 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_568 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_567 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_566 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_565 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_564 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_563 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_562 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_561 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_8 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_8;

architecture SYN_STRUCTURAL of RCA_generic_N64_8 is

   component FA_497
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_498
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_499
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_500
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_501
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_502
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_503
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_504
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_505
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_506
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_507
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_508
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_509
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_510
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_511
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_512
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_513
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_514
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_515
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_516
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_517
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_518
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_519
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_520
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_521
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_522
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_523
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_524
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_525
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_526
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_527
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_528
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_529
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_530
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_531
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_532
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_533
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_534
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_535
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_536
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_537
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_538
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_539
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_540
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_541
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_542
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_543
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_544
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_545
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_546
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_547
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_548
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_549
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_550
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_551
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_552
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_553
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_554
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_555
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_556
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_557
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_558
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_559
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_560
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_560 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_559 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_558 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_557 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_556 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_555 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_554 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_553 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_552 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_551 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_550 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_549 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_548 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_547 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_546 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_545 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_544 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_543 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_542 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_541 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_540 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_539 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_538 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_537 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_536 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_535 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_534 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_533 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_532 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_531 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_530 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_529 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_528 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_527 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_526 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_525 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_524 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_523 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_522 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_521 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_520 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_519 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_518 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_517 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_516 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_515 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_514 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_513 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_512 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_511 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_510 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_509 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_508 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_507 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_506 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_505 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_504 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_503 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_502 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_501 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_500 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_499 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_498 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_497 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_7 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_7;

architecture SYN_STRUCTURAL of RCA_generic_N64_7 is

   component FA_433
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_434
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_435
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_436
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_437
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_438
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_439
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_440
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_441
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_442
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_443
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_444
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_445
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_446
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_447
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_448
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_449
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_450
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_451
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_452
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_453
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_454
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_455
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_456
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_457
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_458
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_459
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_460
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_461
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_462
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_463
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_464
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_465
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_466
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_467
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_468
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_469
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_470
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_471
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_472
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_473
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_474
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_475
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_476
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_477
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_478
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_479
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_480
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_481
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_482
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_483
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_484
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_485
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_486
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_487
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_488
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_489
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_490
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_491
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_492
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_493
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_494
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_495
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_496
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_496 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_495 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_494 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_493 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_492 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_491 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_490 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_489 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_488 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_487 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_486 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_485 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_484 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_483 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_482 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_481 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_480 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_479 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_478 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_477 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_476 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_475 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_474 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_473 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_472 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_471 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_470 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_469 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_468 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_467 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_466 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_465 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_464 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_463 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_462 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_461 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_460 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_459 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_458 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_457 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_456 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_455 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_454 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_453 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_452 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_451 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_450 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_449 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_448 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_447 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_446 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_445 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_444 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_443 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_442 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_441 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_440 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_439 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_438 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_437 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_436 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_435 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_434 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_433 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_6 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_6;

architecture SYN_STRUCTURAL of RCA_generic_N64_6 is

   component FA_369
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_370
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_371
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_372
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_373
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_374
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_375
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_376
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_377
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_378
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_379
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_380
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_381
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_382
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_383
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_384
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_385
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_386
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_387
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_388
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_389
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_390
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_391
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_392
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_393
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_394
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_395
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_396
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_397
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_398
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_399
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_400
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_401
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_402
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_403
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_404
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_405
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_406
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_407
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_408
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_409
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_410
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_411
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_412
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_413
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_414
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_415
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_416
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_417
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_418
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_419
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_420
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_421
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_422
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_423
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_424
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_425
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_426
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_427
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_428
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_429
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_430
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_431
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_432
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_432 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_431 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_430 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_429 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_428 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_427 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_426 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_425 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_424 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_423 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_422 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_421 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_420 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_419 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_418 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_417 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_416 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_415 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_414 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_413 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_412 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_411 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_410 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_409 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_408 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_407 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_406 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_405 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_404 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_403 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_402 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_401 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_400 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_399 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_398 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_397 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_396 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_395 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_394 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_393 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_392 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_391 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_390 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_389 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_388 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_387 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_386 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_385 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_384 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_383 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_382 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_381 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_380 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_379 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_378 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_377 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_376 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_375 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_374 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_373 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_372 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_371 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_370 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_369 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_5 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_5;

architecture SYN_STRUCTURAL of RCA_generic_N64_5 is

   component FA_305
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_306
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_307
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_308
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_309
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_310
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_311
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_312
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_313
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_314
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_315
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_316
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_317
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_318
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_319
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_320
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_321
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_322
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_323
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_324
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_325
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_326
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_327
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_328
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_329
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_330
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_331
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_332
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_333
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_334
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_335
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_336
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_337
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_338
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_339
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_340
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_341
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_342
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_343
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_344
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_345
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_346
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_347
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_348
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_349
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_350
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_351
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_352
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_353
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_354
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_355
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_356
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_357
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_358
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_359
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_360
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_361
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_362
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_363
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_364
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_365
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_366
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_367
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_368
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_368 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_367 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_366 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_365 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_364 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_363 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_362 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_361 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_360 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_359 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_358 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_357 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_356 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_355 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_354 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_353 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_352 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_351 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_350 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_349 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_348 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_347 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_346 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_345 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_344 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_343 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_342 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_341 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_340 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_339 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_338 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_337 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_336 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_335 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_334 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_333 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_332 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_331 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_330 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_329 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_328 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_327 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_326 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_325 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_324 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_323 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_322 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_321 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_320 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_319 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_318 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_317 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_316 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_315 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_314 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_313 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_312 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_311 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_310 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_309 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_308 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_307 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_306 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_305 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_4 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_4;

architecture SYN_STRUCTURAL of RCA_generic_N64_4 is

   component FA_241
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_242
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_243
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_244
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_245
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_246
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_247
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_248
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_249
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_250
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_251
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_252
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_253
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_254
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_255
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_256
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_257
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_258
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_259
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_260
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_261
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_262
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_263
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_264
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_265
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_266
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_267
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_268
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_269
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_270
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_271
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_272
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_273
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_274
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_275
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_276
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_277
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_278
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_279
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_280
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_281
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_282
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_283
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_284
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_285
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_286
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_287
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_288
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_289
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_290
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_291
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_292
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_293
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_294
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_295
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_296
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_297
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_298
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_299
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_300
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_301
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_302
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_303
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_304
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_304 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_303 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_302 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_301 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_300 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_299 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_298 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_297 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_296 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_295 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_294 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_293 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_292 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_291 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_290 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_289 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_288 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_287 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_286 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_285 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_284 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_283 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_282 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_281 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_280 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_279 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_278 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_277 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_276 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_275 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_274 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_273 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_272 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_271 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_270 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_269 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_268 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_267 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_266 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_265 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_264 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_263 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_262 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_261 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_260 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_259 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_258 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_257 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_256 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_255 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_254 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_253 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_252 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_251 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_250 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_249 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_248 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_247 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_246 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_245 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_244 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_243 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_242 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_241 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_3 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_3;

architecture SYN_STRUCTURAL of RCA_generic_N64_3 is

   component FA_177
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_178
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_179
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_180
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_181
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_182
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_183
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_184
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_185
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_186
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_187
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_188
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_189
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_190
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_191
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_192
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_193
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_194
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_195
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_196
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_197
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_198
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_199
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_200
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_201
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_202
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_203
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_204
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_205
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_206
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_207
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_208
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_209
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_210
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_211
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_212
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_213
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_214
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_215
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_216
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_217
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_218
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_219
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_220
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_221
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_222
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_223
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_224
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_225
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_226
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_227
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_228
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_229
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_230
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_231
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_232
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_233
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_234
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_235
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_236
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_237
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_238
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_239
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_240
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_240 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_239 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_238 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_237 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_236 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_235 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_234 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_233 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_232 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_231 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_230 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_229 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_228 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_227 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_226 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_225 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_224 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_223 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_222 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_221 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_220 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_219 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_218 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_217 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_216 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_215 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_214 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_213 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_212 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_211 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_210 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_209 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_208 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_207 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_206 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_205 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_204 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_203 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_202 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_201 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_200 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_199 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_198 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_197 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_196 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_195 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_194 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_193 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_192 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_191 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_190 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_189 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_188 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_187 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_186 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_185 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_184 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_183 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_182 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_181 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_180 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_179 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_178 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_177 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_2 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_2;

architecture SYN_STRUCTURAL of RCA_generic_N64_2 is

   component FA_113
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_114
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_115
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_116
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_117
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_118
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_119
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_120
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_121
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_122
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_123
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_124
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_125
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_126
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_127
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_128
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_129
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_130
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_131
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_132
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_133
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_134
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_135
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_136
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_137
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_138
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_139
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_140
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_141
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_142
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_143
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_144
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_145
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_146
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_147
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_148
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_149
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_150
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_151
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_152
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_153
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_154
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_155
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_156
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_157
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_158
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_159
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_160
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_161
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_162
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_163
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_164
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_165
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_166
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_167
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_168
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_169
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_170
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_171
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_172
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_173
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_174
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_175
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_176
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_176 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_175 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_174 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_173 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_172 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_171 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_170 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_169 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_168 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_167 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_166 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_165 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_164 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_163 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_162 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_161 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_160 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_159 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_158 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_157 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_156 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_155 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_154 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_153 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_152 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_151 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_150 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_149 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_148 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_147 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_146 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_145 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_144 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_143 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_142 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_141 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_140 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_139 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_138 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_137 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_136 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_135 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_134 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_133 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_132 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_131 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_130 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_129 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_128 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_127 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_126 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_125 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_124 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_123 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_122 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_121 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_120 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_119 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_118 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_117 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_116 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_115 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_114 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_113 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_1 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_1;

architecture SYN_STRUCTURAL of RCA_generic_N64_1 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_96
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_97
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_98
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_99
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_100
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_101
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_102
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_103
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_104
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_105
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_106
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_107
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_108
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_109
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_110
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_111
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_112
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_112 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_111 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1),
                           Co => CTMP_2_port);
   FAI_3 : FA_110 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2),
                           Co => CTMP_3_port);
   FAI_4 : FA_109 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3),
                           Co => CTMP_4_port);
   FAI_5 : FA_108 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4),
                           Co => CTMP_5_port);
   FAI_6 : FA_107 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5),
                           Co => CTMP_6_port);
   FAI_7 : FA_106 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6),
                           Co => CTMP_7_port);
   FAI_8 : FA_105 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7),
                           Co => CTMP_8_port);
   FAI_9 : FA_104 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8),
                           Co => CTMP_9_port);
   FAI_10 : FA_103 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_102 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_101 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_100 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_99 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_98 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_97 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_96 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_95 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_94 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_93 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_92 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_91 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_90 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_89 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_88 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_87 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_86 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_85 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_84 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_83 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_82 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_81 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_80 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_79 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_78 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_77 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_76 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_75 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_74 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_73 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_72 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_71 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_70 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_69 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_68 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_67 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_66 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_65 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_64 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_63 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_62 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_61 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_60 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_59 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_58 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_57 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_56 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_55 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_54 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_53 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_52 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_51 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_50 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_49 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_15 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_15;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_15 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net141885, net141886, net141888, net142145, net146767, net146765, 
      net146761, net146759, net146781, net146779, net146777, net146775, 
      net146793, net146791, net146789, net146787, net146785, net146805, 
      net146803, net146801, net146799, net146797, net146817, net146815, 
      net146813, net146811, net146809, net148625, net142137, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
      n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
      n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
      n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, 
      n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, 
      n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, 
      n406, n407, n408 : std_logic;

begin
   
   U1 : AND2_X2 port map( A1 => n153, A2 => n149, ZN => n139);
   U2 : INV_X1 port map( A => E(1), ZN => n140);
   U3 : BUF_X1 port map( A => net141885, Z => net146781);
   U4 : OR2_X1 port map( A1 => net142145, A2 => n140, ZN => n160);
   U5 : BUF_X4 port map( A => n145, Z => net146767);
   U6 : NOR2_X1 port map( A1 => n151, A2 => SEL(2), ZN => n153);
   U7 : AND2_X1 port map( A1 => SEL(1), A2 => n152, ZN => n141);
   U8 : BUF_X2 port map( A => net141886, Z => net146787);
   U9 : NOR2_X1 port map( A1 => n143, A2 => n144, ZN => n142);
   U10 : AND2_X1 port map( A1 => net141886, A2 => D(1), ZN => n143);
   U11 : AND2_X1 port map( A1 => B(1), A2 => n139, ZN => n144);
   U12 : CLKBUF_X1 port map( A => n139, Z => net146797);
   U13 : AND2_X1 port map( A1 => n152, A2 => SEL(1), ZN => n145);
   U14 : AND2_X1 port map( A1 => n148, A2 => n149, ZN => n146);
   U15 : AND2_X2 port map( A1 => n154, A2 => SEL(1), ZN => net141886);
   U16 : INV_X1 port map( A => n151, ZN => n147);
   U17 : NOR2_X1 port map( A1 => n147, A2 => SEL(1), ZN => n150);
   U18 : INV_X1 port map( A => SEL(1), ZN => n149);
   U19 : INV_X1 port map( A => SEL(0), ZN => n151);
   U20 : NOR2_X1 port map( A1 => n151, A2 => SEL(2), ZN => n154);
   U21 : NOR2_X1 port map( A1 => n155, A2 => SEL(2), ZN => n148);
   U22 : NOR2_X1 port map( A1 => SEL(2), A2 => n155, ZN => n152);
   U23 : NAND2_X1 port map( A1 => SEL(2), A2 => E(0), ZN => net142137);
   U24 : OAI21_X1 port map( B1 => SEL(2), B2 => n150, A => net148625, ZN => 
                           net142145);
   U25 : BUF_X1 port map( A => SEL(0), Z => n155);
   U26 : NAND2_X1 port map( A1 => n148, A2 => n149, ZN => net148625);
   U27 : NAND4_X1 port map( A1 => n158, A2 => net142137, A3 => n156, A4 => n157
                           , ZN => Y(0));
   U28 : NAND2_X1 port map( A1 => D(0), A2 => net141886, ZN => n157);
   U29 : NAND2_X1 port map( A1 => B(0), A2 => n139, ZN => n156);
   U30 : AOI22_X1 port map( A1 => C(0), A2 => n141, B1 => n146, B2 => A(0), ZN 
                           => n158);
   U31 : NAND3_X1 port map( A1 => n160, A2 => n159, A3 => n142, ZN => Y(1));
   U32 : BUF_X4 port map( A => net141888, Z => net146809);
   U33 : CLKBUF_X1 port map( A => net141888, Z => net146815);
   U34 : BUF_X4 port map( A => net141885, Z => net146779);
   U35 : CLKBUF_X1 port map( A => net141886, Z => net146791);
   U36 : CLKBUF_X1 port map( A => net141886, Z => net146789);
   U37 : CLKBUF_X1 port map( A => net141886, Z => net146785);
   U38 : CLKBUF_X1 port map( A => net141888, Z => net146811);
   U39 : CLKBUF_X1 port map( A => net141888, Z => net146813);
   U40 : CLKBUF_X1 port map( A => n139, Z => net146803);
   U41 : CLKBUF_X1 port map( A => n139, Z => net146801);
   U42 : CLKBUF_X1 port map( A => n139, Z => net146799);
   U43 : CLKBUF_X1 port map( A => n145, Z => net146759);
   U44 : CLKBUF_X1 port map( A => n145, Z => net146761);
   U45 : CLKBUF_X1 port map( A => n145, Z => net146765);
   U46 : CLKBUF_X1 port map( A => net141885, Z => net146775);
   U47 : CLKBUF_X1 port map( A => net141885, Z => net146777);
   U48 : CLKBUF_X1 port map( A => net141888, Z => net146817);
   U49 : CLKBUF_X1 port map( A => n139, Z => net146805);
   U50 : CLKBUF_X1 port map( A => net141886, Z => net146793);
   U51 : INV_X1 port map( A => net142145, ZN => net141888);
   U52 : INV_X1 port map( A => net148625, ZN => net141885);
   U53 : AOI22_X1 port map( A1 => C(1), A2 => n145, B1 => A(1), B2 => net141885
                           , ZN => n159);
   U54 : NAND2_X1 port map( A1 => E(2), A2 => net141888, ZN => n164);
   U55 : NAND2_X1 port map( A1 => B(2), A2 => net146805, ZN => n163);
   U56 : NAND2_X1 port map( A1 => D(2), A2 => net146787, ZN => n162);
   U57 : AOI22_X1 port map( A1 => C(2), A2 => net146759, B1 => A(2), B2 => 
                           net146775, ZN => n161);
   U58 : NAND4_X1 port map( A1 => n164, A2 => n163, A3 => n162, A4 => n161, ZN 
                           => Y(2));
   U59 : NAND2_X1 port map( A1 => E(3), A2 => net146815, ZN => n168);
   U60 : NAND2_X1 port map( A1 => B(3), A2 => net146797, ZN => n167);
   U61 : NAND2_X1 port map( A1 => D(3), A2 => net146785, ZN => n166);
   U62 : AOI22_X1 port map( A1 => C(3), A2 => net146759, B1 => A(3), B2 => 
                           net146781, ZN => n165);
   U63 : NAND4_X1 port map( A1 => n168, A2 => n167, A3 => n166, A4 => n165, ZN 
                           => Y(3));
   U64 : NAND2_X1 port map( A1 => E(4), A2 => net146811, ZN => n172);
   U65 : NAND2_X1 port map( A1 => B(4), A2 => net146799, ZN => n171);
   U66 : NAND2_X1 port map( A1 => D(4), A2 => net146793, ZN => n170);
   U67 : AOI22_X1 port map( A1 => C(4), A2 => net146761, B1 => A(4), B2 => 
                           net146781, ZN => n169);
   U68 : NAND4_X1 port map( A1 => n172, A2 => n171, A3 => n170, A4 => n169, ZN 
                           => Y(4));
   U69 : NAND2_X1 port map( A1 => E(5), A2 => net146813, ZN => n176);
   U70 : NAND2_X1 port map( A1 => B(5), A2 => net146801, ZN => n175);
   U71 : NAND2_X1 port map( A1 => D(5), A2 => net146791, ZN => n174);
   U72 : AOI22_X1 port map( A1 => C(5), A2 => net146761, B1 => A(5), B2 => 
                           net146781, ZN => n173);
   U73 : NAND4_X1 port map( A1 => n176, A2 => n175, A3 => n174, A4 => n173, ZN 
                           => Y(5));
   U74 : NAND2_X1 port map( A1 => E(6), A2 => net146817, ZN => n180);
   U75 : NAND2_X1 port map( A1 => B(6), A2 => net146803, ZN => n179);
   U76 : NAND2_X1 port map( A1 => D(6), A2 => net146789, ZN => n178);
   U77 : AOI22_X1 port map( A1 => C(6), A2 => net146765, B1 => A(6), B2 => 
                           net146777, ZN => n177);
   U78 : NAND4_X1 port map( A1 => n180, A2 => n179, A3 => n178, A4 => n177, ZN 
                           => Y(6));
   U79 : NAND2_X1 port map( A1 => E(7), A2 => net146809, ZN => n184);
   U80 : NAND2_X1 port map( A1 => B(7), A2 => net146803, ZN => n183);
   U81 : NAND2_X1 port map( A1 => D(7), A2 => net146787, ZN => n182);
   U82 : AOI22_X1 port map( A1 => C(7), A2 => net146767, B1 => A(7), B2 => 
                           net146779, ZN => n181);
   U83 : NAND4_X1 port map( A1 => n184, A2 => n183, A3 => n182, A4 => n181, ZN 
                           => Y(7));
   U84 : NAND2_X1 port map( A1 => E(8), A2 => net146809, ZN => n188);
   U85 : NAND2_X1 port map( A1 => B(8), A2 => net146803, ZN => n187);
   U86 : NAND2_X1 port map( A1 => D(8), A2 => net146785, ZN => n186);
   U87 : AOI22_X1 port map( A1 => C(8), A2 => net146767, B1 => A(8), B2 => 
                           net146779, ZN => n185);
   U88 : NAND4_X1 port map( A1 => n188, A2 => n187, A3 => n186, A4 => n185, ZN 
                           => Y(8));
   U89 : NAND2_X1 port map( A1 => E(9), A2 => net146809, ZN => n192);
   U90 : NAND2_X1 port map( A1 => B(9), A2 => net146803, ZN => n191);
   U91 : NAND2_X1 port map( A1 => D(9), A2 => net146793, ZN => n190);
   U92 : AOI22_X1 port map( A1 => C(9), A2 => net146767, B1 => A(9), B2 => 
                           net146779, ZN => n189);
   U93 : NAND4_X1 port map( A1 => n192, A2 => n191, A3 => n190, A4 => n189, ZN 
                           => Y(9));
   U94 : NAND2_X1 port map( A1 => E(10), A2 => net146809, ZN => n196);
   U95 : NAND2_X1 port map( A1 => B(10), A2 => net146803, ZN => n195);
   U96 : NAND2_X1 port map( A1 => D(10), A2 => net146791, ZN => n194);
   U97 : AOI22_X1 port map( A1 => C(10), A2 => net146767, B1 => A(10), B2 => 
                           net146779, ZN => n193);
   U98 : NAND4_X1 port map( A1 => n196, A2 => n195, A3 => n194, A4 => n193, ZN 
                           => Y(10));
   U99 : NAND2_X1 port map( A1 => E(11), A2 => net146809, ZN => n200);
   U100 : NAND2_X1 port map( A1 => B(11), A2 => net146803, ZN => n199);
   U101 : NAND2_X1 port map( A1 => D(11), A2 => net146789, ZN => n198);
   U102 : AOI22_X1 port map( A1 => C(11), A2 => net146767, B1 => A(11), B2 => 
                           net146779, ZN => n197);
   U103 : NAND4_X1 port map( A1 => n200, A2 => n199, A3 => n198, A4 => n197, ZN
                           => Y(11));
   U104 : NAND2_X1 port map( A1 => E(12), A2 => net146809, ZN => n204);
   U105 : NAND2_X1 port map( A1 => B(12), A2 => net146797, ZN => n203);
   U106 : NAND2_X1 port map( A1 => D(12), A2 => net146787, ZN => n202);
   U107 : AOI22_X1 port map( A1 => C(12), A2 => net146767, B1 => A(12), B2 => 
                           net146779, ZN => n201);
   U108 : NAND4_X1 port map( A1 => n204, A2 => n203, A3 => n202, A4 => n201, ZN
                           => Y(12));
   U109 : NAND2_X1 port map( A1 => E(13), A2 => net146809, ZN => n208);
   U110 : NAND2_X1 port map( A1 => B(13), A2 => net146797, ZN => n207);
   U111 : NAND2_X1 port map( A1 => D(13), A2 => net146785, ZN => n206);
   U112 : AOI22_X1 port map( A1 => C(13), A2 => net146767, B1 => A(13), B2 => 
                           net146779, ZN => n205);
   U113 : NAND4_X1 port map( A1 => n208, A2 => n207, A3 => n206, A4 => n205, ZN
                           => Y(13));
   U114 : NAND2_X1 port map( A1 => E(14), A2 => net146809, ZN => n212);
   U115 : NAND2_X1 port map( A1 => B(14), A2 => net146797, ZN => n211);
   U116 : NAND2_X1 port map( A1 => D(14), A2 => net146793, ZN => n210);
   U117 : AOI22_X1 port map( A1 => C(14), A2 => net146767, B1 => A(14), B2 => 
                           net146779, ZN => n209);
   U118 : NAND4_X1 port map( A1 => n212, A2 => n211, A3 => n210, A4 => n209, ZN
                           => Y(14));
   U119 : NAND2_X1 port map( A1 => E(15), A2 => net146809, ZN => n216);
   U120 : NAND2_X1 port map( A1 => B(15), A2 => net146797, ZN => n215);
   U121 : NAND2_X1 port map( A1 => D(15), A2 => net146791, ZN => n214);
   U122 : AOI22_X1 port map( A1 => C(15), A2 => net146767, B1 => A(15), B2 => 
                           net146779, ZN => n213);
   U123 : NAND4_X1 port map( A1 => n216, A2 => n215, A3 => n214, A4 => n213, ZN
                           => Y(15));
   U124 : NAND2_X1 port map( A1 => E(16), A2 => net146809, ZN => n220);
   U125 : NAND2_X1 port map( A1 => B(16), A2 => net146797, ZN => n219);
   U126 : NAND2_X1 port map( A1 => D(16), A2 => net146789, ZN => n218);
   U127 : AOI22_X1 port map( A1 => C(16), A2 => net146767, B1 => A(16), B2 => 
                           net146779, ZN => n217);
   U128 : NAND4_X1 port map( A1 => n220, A2 => n219, A3 => n218, A4 => n217, ZN
                           => Y(16));
   U129 : NAND2_X1 port map( A1 => E(17), A2 => net146809, ZN => n224);
   U130 : NAND2_X1 port map( A1 => B(17), A2 => net146797, ZN => n223);
   U131 : NAND2_X1 port map( A1 => D(17), A2 => net146787, ZN => n222);
   U132 : AOI22_X1 port map( A1 => C(17), A2 => net146767, B1 => A(17), B2 => 
                           net146779, ZN => n221);
   U133 : NAND4_X1 port map( A1 => n224, A2 => n223, A3 => n222, A4 => n221, ZN
                           => Y(17));
   U134 : NAND2_X1 port map( A1 => E(18), A2 => net146817, ZN => n228);
   U135 : NAND2_X1 port map( A1 => B(18), A2 => net146797, ZN => n227);
   U136 : NAND2_X1 port map( A1 => D(18), A2 => net146785, ZN => n226);
   U137 : AOI22_X1 port map( A1 => C(18), A2 => net146767, B1 => A(18), B2 => 
                           net146779, ZN => n225);
   U138 : NAND4_X1 port map( A1 => n228, A2 => n227, A3 => n226, A4 => n225, ZN
                           => Y(18));
   U139 : NAND2_X1 port map( A1 => E(19), A2 => net146809, ZN => n232);
   U140 : NAND2_X1 port map( A1 => B(19), A2 => net146797, ZN => n231);
   U141 : NAND2_X1 port map( A1 => D(19), A2 => net146793, ZN => n230);
   U142 : AOI22_X1 port map( A1 => C(19), A2 => net146767, B1 => A(19), B2 => 
                           net146779, ZN => n229);
   U143 : NAND4_X1 port map( A1 => n232, A2 => n231, A3 => n230, A4 => n229, ZN
                           => Y(19));
   U144 : NAND2_X1 port map( A1 => E(20), A2 => net146817, ZN => n236);
   U145 : NAND2_X1 port map( A1 => B(20), A2 => net146797, ZN => n235);
   U146 : NAND2_X1 port map( A1 => D(20), A2 => net146791, ZN => n234);
   U147 : AOI22_X1 port map( A1 => C(20), A2 => net146767, B1 => A(20), B2 => 
                           net146779, ZN => n233);
   U148 : NAND4_X1 port map( A1 => n236, A2 => n235, A3 => n234, A4 => n233, ZN
                           => Y(20));
   U149 : NAND2_X1 port map( A1 => E(21), A2 => net146809, ZN => n240);
   U150 : NAND2_X1 port map( A1 => B(21), A2 => net146797, ZN => n239);
   U151 : NAND2_X1 port map( A1 => D(21), A2 => net146789, ZN => n238);
   U152 : AOI22_X1 port map( A1 => C(21), A2 => net146767, B1 => A(21), B2 => 
                           net146779, ZN => n237);
   U153 : NAND4_X1 port map( A1 => n240, A2 => n239, A3 => n238, A4 => n237, ZN
                           => Y(21));
   U154 : NAND2_X1 port map( A1 => E(22), A2 => net146817, ZN => n244);
   U155 : NAND2_X1 port map( A1 => B(22), A2 => net146797, ZN => n243);
   U156 : NAND2_X1 port map( A1 => D(22), A2 => net146787, ZN => n242);
   U157 : AOI22_X1 port map( A1 => C(22), A2 => net146767, B1 => A(22), B2 => 
                           net146779, ZN => n241);
   U158 : NAND4_X1 port map( A1 => n244, A2 => n243, A3 => n242, A4 => n241, ZN
                           => Y(22));
   U159 : NAND2_X1 port map( A1 => E(23), A2 => net146809, ZN => n248);
   U160 : NAND2_X1 port map( A1 => B(23), A2 => net146797, ZN => n247);
   U161 : NAND2_X1 port map( A1 => D(23), A2 => net146785, ZN => n246);
   U162 : AOI22_X1 port map( A1 => C(23), A2 => net146767, B1 => A(23), B2 => 
                           net146779, ZN => n245);
   U163 : NAND4_X1 port map( A1 => n248, A2 => n247, A3 => n246, A4 => n245, ZN
                           => Y(23));
   U164 : NAND2_X1 port map( A1 => E(24), A2 => net146817, ZN => n252);
   U165 : NAND2_X1 port map( A1 => B(24), A2 => net146799, ZN => n251);
   U166 : NAND2_X1 port map( A1 => D(24), A2 => net146793, ZN => n250);
   U167 : AOI22_X1 port map( A1 => C(24), A2 => net146767, B1 => A(24), B2 => 
                           net146779, ZN => n249);
   U168 : NAND4_X1 port map( A1 => n252, A2 => n251, A3 => n250, A4 => n249, ZN
                           => Y(24));
   U169 : NAND2_X1 port map( A1 => E(25), A2 => net146809, ZN => n256);
   U170 : NAND2_X1 port map( A1 => B(25), A2 => net146799, ZN => n255);
   U171 : NAND2_X1 port map( A1 => D(25), A2 => net146791, ZN => n254);
   U172 : AOI22_X1 port map( A1 => C(25), A2 => net146767, B1 => A(25), B2 => 
                           net146779, ZN => n253);
   U173 : NAND4_X1 port map( A1 => n256, A2 => n255, A3 => n254, A4 => n253, ZN
                           => Y(25));
   U174 : NAND2_X1 port map( A1 => E(26), A2 => net146817, ZN => n260);
   U175 : NAND2_X1 port map( A1 => B(26), A2 => net146799, ZN => n259);
   U176 : NAND2_X1 port map( A1 => D(26), A2 => net146789, ZN => n258);
   U177 : AOI22_X1 port map( A1 => C(26), A2 => net146767, B1 => A(26), B2 => 
                           net146779, ZN => n257);
   U178 : NAND4_X1 port map( A1 => n260, A2 => n259, A3 => n258, A4 => n257, ZN
                           => Y(26));
   U179 : NAND2_X1 port map( A1 => E(27), A2 => net146809, ZN => n264);
   U180 : NAND2_X1 port map( A1 => B(27), A2 => net146799, ZN => n263);
   U181 : NAND2_X1 port map( A1 => D(27), A2 => net146787, ZN => n262);
   U182 : AOI22_X1 port map( A1 => C(27), A2 => net146767, B1 => A(27), B2 => 
                           net146779, ZN => n261);
   U183 : NAND4_X1 port map( A1 => n264, A2 => n263, A3 => n262, A4 => n261, ZN
                           => Y(27));
   U184 : NAND2_X1 port map( A1 => E(28), A2 => net146817, ZN => n268);
   U185 : NAND2_X1 port map( A1 => B(28), A2 => net146799, ZN => n267);
   U186 : NAND2_X1 port map( A1 => D(28), A2 => net146785, ZN => n266);
   U187 : AOI22_X1 port map( A1 => C(28), A2 => net146767, B1 => A(28), B2 => 
                           net146779, ZN => n265);
   U188 : NAND4_X1 port map( A1 => n268, A2 => n267, A3 => n266, A4 => n265, ZN
                           => Y(28));
   U189 : NAND2_X1 port map( A1 => E(29), A2 => net146809, ZN => n272);
   U190 : NAND2_X1 port map( A1 => B(29), A2 => net146799, ZN => n271);
   U191 : NAND2_X1 port map( A1 => D(29), A2 => net146793, ZN => n270);
   U192 : AOI22_X1 port map( A1 => C(29), A2 => net146767, B1 => A(29), B2 => 
                           net146779, ZN => n269);
   U193 : NAND4_X1 port map( A1 => n272, A2 => n271, A3 => n270, A4 => n269, ZN
                           => Y(29));
   U194 : NAND2_X1 port map( A1 => E(30), A2 => net146817, ZN => n276);
   U195 : NAND2_X1 port map( A1 => B(30), A2 => net146799, ZN => n275);
   U196 : NAND2_X1 port map( A1 => D(30), A2 => net146791, ZN => n274);
   U197 : AOI22_X1 port map( A1 => C(30), A2 => net146767, B1 => A(30), B2 => 
                           net146777, ZN => n273);
   U198 : NAND4_X1 port map( A1 => n276, A2 => n275, A3 => n274, A4 => n273, ZN
                           => Y(30));
   U199 : NAND2_X1 port map( A1 => E(31), A2 => net146809, ZN => n280);
   U200 : NAND2_X1 port map( A1 => B(31), A2 => net146799, ZN => n279);
   U201 : NAND2_X1 port map( A1 => D(31), A2 => net146789, ZN => n278);
   U202 : AOI22_X1 port map( A1 => C(31), A2 => net146765, B1 => A(31), B2 => 
                           net146779, ZN => n277);
   U203 : NAND4_X1 port map( A1 => n280, A2 => n279, A3 => n278, A4 => n277, ZN
                           => Y(31));
   U204 : NAND2_X1 port map( A1 => E(32), A2 => net146817, ZN => n284);
   U205 : NAND2_X1 port map( A1 => B(32), A2 => net146799, ZN => n283);
   U206 : NAND2_X1 port map( A1 => D(32), A2 => net146787, ZN => n282);
   U207 : AOI22_X1 port map( A1 => C(32), A2 => net146767, B1 => A(32), B2 => 
                           net146779, ZN => n281);
   U208 : NAND4_X1 port map( A1 => n284, A2 => n283, A3 => n282, A4 => n281, ZN
                           => Y(32));
   U209 : NAND2_X1 port map( A1 => E(33), A2 => net146817, ZN => n288);
   U210 : NAND2_X1 port map( A1 => B(33), A2 => net146799, ZN => n287);
   U211 : NAND2_X1 port map( A1 => D(33), A2 => net146785, ZN => n286);
   U212 : AOI22_X1 port map( A1 => C(33), A2 => net146767, B1 => A(33), B2 => 
                           net146779, ZN => n285);
   U213 : NAND4_X1 port map( A1 => n288, A2 => n287, A3 => n286, A4 => n285, ZN
                           => Y(33));
   U214 : NAND2_X1 port map( A1 => E(34), A2 => net146817, ZN => n292);
   U215 : NAND2_X1 port map( A1 => B(34), A2 => net146799, ZN => n291);
   U216 : NAND2_X1 port map( A1 => D(34), A2 => net146793, ZN => n290);
   U217 : AOI22_X1 port map( A1 => C(34), A2 => net146765, B1 => A(34), B2 => 
                           net146777, ZN => n289);
   U218 : NAND4_X1 port map( A1 => n292, A2 => n291, A3 => n290, A4 => n289, ZN
                           => Y(34));
   U219 : NAND2_X1 port map( A1 => E(35), A2 => net146809, ZN => n296);
   U220 : NAND2_X1 port map( A1 => B(35), A2 => net146799, ZN => n295);
   U221 : NAND2_X1 port map( A1 => D(35), A2 => net146791, ZN => n294);
   U222 : AOI22_X1 port map( A1 => C(35), A2 => net146767, B1 => A(35), B2 => 
                           net146779, ZN => n293);
   U223 : NAND4_X1 port map( A1 => n296, A2 => n295, A3 => n294, A4 => n293, ZN
                           => Y(35));
   U224 : NAND2_X1 port map( A1 => E(36), A2 => net146813, ZN => n300);
   U225 : NAND2_X1 port map( A1 => B(36), A2 => net146801, ZN => n299);
   U226 : NAND2_X1 port map( A1 => D(36), A2 => net146789, ZN => n298);
   U227 : AOI22_X1 port map( A1 => C(36), A2 => net146765, B1 => A(36), B2 => 
                           net146779, ZN => n297);
   U228 : NAND4_X1 port map( A1 => n300, A2 => n299, A3 => n298, A4 => n297, ZN
                           => Y(36));
   U229 : NAND2_X1 port map( A1 => E(37), A2 => net146809, ZN => n304);
   U230 : NAND2_X1 port map( A1 => B(37), A2 => net146801, ZN => n303);
   U231 : NAND2_X1 port map( A1 => D(37), A2 => net146787, ZN => n302);
   U232 : AOI22_X1 port map( A1 => C(37), A2 => net146767, B1 => A(37), B2 => 
                           net146779, ZN => n301);
   U233 : NAND4_X1 port map( A1 => n304, A2 => n303, A3 => n302, A4 => n301, ZN
                           => Y(37));
   U234 : NAND2_X1 port map( A1 => E(38), A2 => net146817, ZN => n308);
   U235 : NAND2_X1 port map( A1 => B(38), A2 => net146801, ZN => n307);
   U236 : NAND2_X1 port map( A1 => D(38), A2 => net146785, ZN => n306);
   U237 : AOI22_X1 port map( A1 => C(38), A2 => net146767, B1 => A(38), B2 => 
                           net146777, ZN => n305);
   U238 : NAND4_X1 port map( A1 => n308, A2 => n307, A3 => n306, A4 => n305, ZN
                           => Y(38));
   U239 : NAND2_X1 port map( A1 => E(39), A2 => net146813, ZN => n312);
   U240 : NAND2_X1 port map( A1 => B(39), A2 => net146801, ZN => n311);
   U241 : NAND2_X1 port map( A1 => D(39), A2 => net146793, ZN => n310);
   U242 : AOI22_X1 port map( A1 => C(39), A2 => net146765, B1 => A(39), B2 => 
                           net146779, ZN => n309);
   U243 : NAND4_X1 port map( A1 => n312, A2 => n311, A3 => n310, A4 => n309, ZN
                           => Y(39));
   U244 : NAND2_X1 port map( A1 => E(40), A2 => net146809, ZN => n316);
   U245 : NAND2_X1 port map( A1 => B(40), A2 => net146801, ZN => n315);
   U246 : NAND2_X1 port map( A1 => D(40), A2 => net146791, ZN => n314);
   U247 : AOI22_X1 port map( A1 => C(40), A2 => net146767, B1 => A(40), B2 => 
                           net146779, ZN => n313);
   U248 : NAND4_X1 port map( A1 => n316, A2 => n315, A3 => n314, A4 => n313, ZN
                           => Y(40));
   U249 : NAND2_X1 port map( A1 => E(41), A2 => net146817, ZN => n320);
   U250 : NAND2_X1 port map( A1 => B(41), A2 => net146801, ZN => n319);
   U251 : NAND2_X1 port map( A1 => D(41), A2 => net146789, ZN => n318);
   U252 : AOI22_X1 port map( A1 => C(41), A2 => net146765, B1 => A(41), B2 => 
                           net146777, ZN => n317);
   U253 : NAND4_X1 port map( A1 => n320, A2 => n319, A3 => n318, A4 => n317, ZN
                           => Y(41));
   U254 : NAND2_X1 port map( A1 => E(42), A2 => net146813, ZN => n324);
   U255 : NAND2_X1 port map( A1 => B(42), A2 => net146801, ZN => n323);
   U256 : NAND2_X1 port map( A1 => D(42), A2 => net146787, ZN => n322);
   U257 : AOI22_X1 port map( A1 => C(42), A2 => net146767, B1 => A(42), B2 => 
                           net146779, ZN => n321);
   U258 : NAND4_X1 port map( A1 => n324, A2 => n323, A3 => n322, A4 => n321, ZN
                           => Y(42));
   U259 : NAND2_X1 port map( A1 => E(43), A2 => net146809, ZN => n328);
   U260 : NAND2_X1 port map( A1 => B(43), A2 => net146801, ZN => n327);
   U261 : NAND2_X1 port map( A1 => D(43), A2 => net146785, ZN => n326);
   U262 : AOI22_X1 port map( A1 => C(43), A2 => net146765, B1 => A(43), B2 => 
                           net146779, ZN => n325);
   U263 : NAND4_X1 port map( A1 => n328, A2 => n327, A3 => n326, A4 => n325, ZN
                           => Y(43));
   U264 : NAND2_X1 port map( A1 => E(44), A2 => net146813, ZN => n332);
   U265 : NAND2_X1 port map( A1 => B(44), A2 => net146801, ZN => n331);
   U266 : NAND2_X1 port map( A1 => D(44), A2 => net146793, ZN => n330);
   U267 : AOI22_X1 port map( A1 => C(44), A2 => net146767, B1 => A(44), B2 => 
                           net146779, ZN => n329);
   U268 : NAND4_X1 port map( A1 => n332, A2 => n331, A3 => n330, A4 => n329, ZN
                           => Y(44));
   U269 : NAND2_X1 port map( A1 => E(45), A2 => net146817, ZN => n336);
   U270 : NAND2_X1 port map( A1 => B(45), A2 => net146801, ZN => n335);
   U271 : NAND2_X1 port map( A1 => D(45), A2 => net146791, ZN => n334);
   U272 : AOI22_X1 port map( A1 => C(45), A2 => net146767, B1 => A(45), B2 => 
                           net146777, ZN => n333);
   U273 : NAND4_X1 port map( A1 => n336, A2 => n335, A3 => n334, A4 => n333, ZN
                           => Y(45));
   U274 : NAND2_X1 port map( A1 => E(46), A2 => net146809, ZN => n340);
   U275 : NAND2_X1 port map( A1 => B(46), A2 => net146801, ZN => n339);
   U276 : NAND2_X1 port map( A1 => D(46), A2 => net146789, ZN => n338);
   U277 : AOI22_X1 port map( A1 => C(46), A2 => net146765, B1 => A(46), B2 => 
                           net146779, ZN => n337);
   U278 : NAND4_X1 port map( A1 => n340, A2 => n339, A3 => n338, A4 => n337, ZN
                           => Y(46));
   U279 : NAND2_X1 port map( A1 => E(47), A2 => net146813, ZN => n344);
   U280 : NAND2_X1 port map( A1 => B(47), A2 => net146801, ZN => n343);
   U281 : NAND2_X1 port map( A1 => D(47), A2 => net146787, ZN => n342);
   U282 : AOI22_X1 port map( A1 => C(47), A2 => net146767, B1 => A(47), B2 => 
                           net146779, ZN => n341);
   U283 : NAND4_X1 port map( A1 => n344, A2 => n343, A3 => n342, A4 => n341, ZN
                           => Y(47));
   U284 : NAND2_X1 port map( A1 => E(48), A2 => net146817, ZN => n348);
   U285 : NAND2_X1 port map( A1 => B(48), A2 => net146803, ZN => n347);
   U286 : NAND2_X1 port map( A1 => D(48), A2 => net146785, ZN => n346);
   U287 : AOI22_X1 port map( A1 => C(48), A2 => net146765, B1 => A(48), B2 => 
                           net146779, ZN => n345);
   U288 : NAND4_X1 port map( A1 => n348, A2 => n347, A3 => n346, A4 => n345, ZN
                           => Y(48));
   U289 : NAND2_X1 port map( A1 => E(49), A2 => net146809, ZN => n352);
   U290 : NAND2_X1 port map( A1 => B(49), A2 => net146803, ZN => n351);
   U291 : NAND2_X1 port map( A1 => D(49), A2 => net146793, ZN => n350);
   U292 : AOI22_X1 port map( A1 => C(49), A2 => net146765, B1 => A(49), B2 => 
                           net146781, ZN => n349);
   U293 : NAND4_X1 port map( A1 => n352, A2 => n351, A3 => n350, A4 => n349, ZN
                           => Y(49));
   U294 : NAND2_X1 port map( A1 => E(50), A2 => net146811, ZN => n356);
   U295 : NAND2_X1 port map( A1 => B(50), A2 => net146803, ZN => n355);
   U296 : NAND2_X1 port map( A1 => D(50), A2 => net146791, ZN => n354);
   U297 : AOI22_X1 port map( A1 => C(50), A2 => net146765, B1 => A(50), B2 => 
                           net146777, ZN => n353);
   U298 : NAND4_X1 port map( A1 => n356, A2 => n355, A3 => n354, A4 => n353, ZN
                           => Y(50));
   U299 : NAND2_X1 port map( A1 => E(51), A2 => net146813, ZN => n360);
   U300 : NAND2_X1 port map( A1 => B(51), A2 => net146803, ZN => n359);
   U301 : NAND2_X1 port map( A1 => D(51), A2 => net146789, ZN => n358);
   U302 : AOI22_X1 port map( A1 => C(51), A2 => net146767, B1 => A(51), B2 => 
                           net146779, ZN => n357);
   U303 : NAND4_X1 port map( A1 => n360, A2 => n359, A3 => n358, A4 => n357, ZN
                           => Y(51));
   U304 : NAND2_X1 port map( A1 => E(52), A2 => net146817, ZN => n364);
   U305 : NAND2_X1 port map( A1 => B(52), A2 => net146803, ZN => n363);
   U306 : NAND2_X1 port map( A1 => D(52), A2 => net146787, ZN => n362);
   U307 : AOI22_X1 port map( A1 => C(52), A2 => net146765, B1 => A(52), B2 => 
                           net146779, ZN => n361);
   U308 : NAND4_X1 port map( A1 => n364, A2 => n363, A3 => n362, A4 => n361, ZN
                           => Y(52));
   U309 : NAND2_X1 port map( A1 => E(53), A2 => net146809, ZN => n368);
   U310 : NAND2_X1 port map( A1 => B(53), A2 => net146803, ZN => n367);
   U311 : NAND2_X1 port map( A1 => D(53), A2 => net146785, ZN => n366);
   U312 : AOI22_X1 port map( A1 => C(53), A2 => net146767, B1 => A(53), B2 => 
                           net146779, ZN => n365);
   U313 : NAND4_X1 port map( A1 => n368, A2 => n367, A3 => n366, A4 => n365, ZN
                           => Y(53));
   U314 : NAND2_X1 port map( A1 => E(54), A2 => net146811, ZN => n372);
   U315 : NAND2_X1 port map( A1 => B(54), A2 => net146803, ZN => n371);
   U316 : NAND2_X1 port map( A1 => D(54), A2 => net146793, ZN => n370);
   U317 : AOI22_X1 port map( A1 => C(54), A2 => net146767, B1 => A(54), B2 => 
                           net146781, ZN => n369);
   U318 : NAND4_X1 port map( A1 => n372, A2 => n371, A3 => n370, A4 => n369, ZN
                           => Y(54));
   U319 : NAND2_X1 port map( A1 => E(55), A2 => net146813, ZN => n376);
   U320 : NAND2_X1 port map( A1 => B(55), A2 => net146803, ZN => n375);
   U321 : NAND2_X1 port map( A1 => D(55), A2 => net146791, ZN => n374);
   U322 : AOI22_X1 port map( A1 => C(55), A2 => net146765, B1 => A(55), B2 => 
                           net146777, ZN => n373);
   U323 : NAND4_X1 port map( A1 => n376, A2 => n375, A3 => n374, A4 => n373, ZN
                           => Y(55));
   U324 : NAND2_X1 port map( A1 => E(56), A2 => net146817, ZN => n380);
   U325 : NAND2_X1 port map( A1 => B(56), A2 => net146803, ZN => n379);
   U326 : NAND2_X1 port map( A1 => D(56), A2 => net146789, ZN => n378);
   U327 : AOI22_X1 port map( A1 => C(56), A2 => net146767, B1 => A(56), B2 => 
                           net146779, ZN => n377);
   U328 : NAND4_X1 port map( A1 => n380, A2 => n379, A3 => n378, A4 => n377, ZN
                           => Y(56));
   U329 : NAND2_X1 port map( A1 => E(57), A2 => net146809, ZN => n384);
   U330 : NAND2_X1 port map( A1 => B(57), A2 => net146803, ZN => n383);
   U331 : NAND2_X1 port map( A1 => D(57), A2 => net146787, ZN => n382);
   U332 : AOI22_X1 port map( A1 => C(57), A2 => net146765, B1 => A(57), B2 => 
                           net146779, ZN => n381);
   U333 : NAND4_X1 port map( A1 => n384, A2 => n383, A3 => n382, A4 => n381, ZN
                           => Y(57));
   U334 : NAND2_X1 port map( A1 => E(58), A2 => net146811, ZN => n388);
   U335 : NAND2_X1 port map( A1 => B(58), A2 => net146803, ZN => n387);
   U336 : NAND2_X1 port map( A1 => D(58), A2 => net146785, ZN => n386);
   U337 : AOI22_X1 port map( A1 => C(58), A2 => net146767, B1 => A(58), B2 => 
                           net146779, ZN => n385);
   U338 : NAND4_X1 port map( A1 => n388, A2 => n387, A3 => n386, A4 => n385, ZN
                           => Y(58));
   U339 : NAND2_X1 port map( A1 => E(59), A2 => net146813, ZN => n392);
   U340 : NAND2_X1 port map( A1 => B(59), A2 => net146803, ZN => n391);
   U341 : NAND2_X1 port map( A1 => D(59), A2 => net146793, ZN => n390);
   U342 : AOI22_X1 port map( A1 => C(59), A2 => net146767, B1 => A(59), B2 => 
                           net146777, ZN => n389);
   U343 : NAND4_X1 port map( A1 => n392, A2 => n391, A3 => n390, A4 => n389, ZN
                           => Y(59));
   U344 : NAND2_X1 port map( A1 => E(60), A2 => net146813, ZN => n396);
   U345 : NAND2_X1 port map( A1 => B(60), A2 => net146805, ZN => n395);
   U346 : NAND2_X1 port map( A1 => D(60), A2 => net146791, ZN => n394);
   U347 : AOI22_X1 port map( A1 => C(60), A2 => net146765, B1 => A(60), B2 => 
                           net146781, ZN => n393);
   U348 : NAND4_X1 port map( A1 => n396, A2 => n395, A3 => n394, A4 => n393, ZN
                           => Y(60));
   U349 : NAND2_X1 port map( A1 => E(61), A2 => net146817, ZN => n400);
   U350 : NAND2_X1 port map( A1 => B(61), A2 => net146805, ZN => n399);
   U351 : NAND2_X1 port map( A1 => D(61), A2 => net146789, ZN => n398);
   U352 : AOI22_X1 port map( A1 => C(61), A2 => net146767, B1 => A(61), B2 => 
                           net146779, ZN => n397);
   U353 : NAND4_X1 port map( A1 => n400, A2 => n399, A3 => n398, A4 => n397, ZN
                           => Y(61));
   U354 : NAND2_X1 port map( A1 => E(62), A2 => net146809, ZN => n404);
   U355 : NAND2_X1 port map( A1 => B(62), A2 => net146805, ZN => n403);
   U356 : NAND2_X1 port map( A1 => D(62), A2 => net146787, ZN => n402);
   U357 : AOI22_X1 port map( A1 => C(62), A2 => net146765, B1 => A(62), B2 => 
                           net146777, ZN => n401);
   U358 : NAND4_X1 port map( A1 => n404, A2 => n403, A3 => n402, A4 => n401, ZN
                           => Y(62));
   U359 : NAND2_X1 port map( A1 => E(63), A2 => net146813, ZN => n408);
   U360 : NAND2_X1 port map( A1 => B(63), A2 => net146805, ZN => n407);
   U361 : NAND2_X1 port map( A1 => D(63), A2 => net146785, ZN => n406);
   U362 : AOI22_X1 port map( A1 => C(63), A2 => net146767, B1 => A(63), B2 => 
                           net146779, ZN => n405);
   U363 : NAND4_X1 port map( A1 => n408, A2 => n407, A3 => n406, A4 => n405, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_14 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_14;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_14 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438, n439, n440, n441 : std_logic;

begin
   
   U1 : BUF_X2 port map( A => n434, Z => n150);
   U2 : BUF_X2 port map( A => n437, Z => n140);
   U3 : BUF_X2 port map( A => n437, Z => n139);
   U4 : OR2_X2 port map( A1 => n176, A2 => n142, ZN => n180);
   U5 : NAND4_X1 port map( A1 => n209, A2 => n208, A3 => n207, A4 => n206, ZN 
                           => Y(6));
   U6 : NAND4_X1 port map( A1 => n201, A2 => n200, A3 => n199, A4 => n198, ZN 
                           => Y(4));
   U7 : NAND4_X1 port map( A1 => n213, A2 => n212, A3 => n211, A4 => n210, ZN 
                           => Y(7));
   U8 : CLKBUF_X1 port map( A => n436, Z => n162);
   U9 : BUF_X1 port map( A => n436, Z => n163);
   U10 : BUF_X2 port map( A => n436, Z => n164);
   U11 : INV_X1 port map( A => n181, ZN => n141);
   U12 : CLKBUF_X1 port map( A => n143, Z => n144);
   U13 : BUF_X2 port map( A => n143, Z => n146);
   U14 : BUF_X2 port map( A => n437, Z => n168);
   U15 : AND4_X2 port map( A1 => n178, A2 => n179, A3 => n181, A4 => n180, ZN 
                           => n143);
   U16 : NAND2_X1 port map( A1 => n177, A2 => n174, ZN => n142);
   U17 : CLKBUF_X1 port map( A => n437, Z => n169);
   U18 : BUF_X1 port map( A => n435, Z => n156);
   U19 : CLKBUF_X1 port map( A => n435, Z => n157);
   U20 : CLKBUF_X1 port map( A => n434, Z => n151);
   U21 : CLKBUF_X1 port map( A => n143, Z => n145);
   U22 : CLKBUF_X1 port map( A => n437, Z => n170);
   U23 : CLKBUF_X1 port map( A => n435, Z => n158);
   U24 : CLKBUF_X1 port map( A => n434, Z => n152);
   U25 : CLKBUF_X1 port map( A => n437, Z => n171);
   U26 : CLKBUF_X1 port map( A => n435, Z => n159);
   U27 : CLKBUF_X1 port map( A => n434, Z => n153);
   U28 : CLKBUF_X1 port map( A => n143, Z => n147);
   U29 : CLKBUF_X1 port map( A => n141, Z => n165);
   U30 : CLKBUF_X1 port map( A => n437, Z => n172);
   U31 : CLKBUF_X1 port map( A => n435, Z => n160);
   U32 : CLKBUF_X1 port map( A => n434, Z => n154);
   U33 : CLKBUF_X1 port map( A => n143, Z => n148);
   U34 : CLKBUF_X1 port map( A => n141, Z => n166);
   U35 : NAND2_X1 port map( A1 => n177, A2 => n175, ZN => n181);
   U36 : CLKBUF_X1 port map( A => n143, Z => n149);
   U37 : CLKBUF_X1 port map( A => n434, Z => n155);
   U38 : CLKBUF_X1 port map( A => n435, Z => n161);
   U39 : CLKBUF_X1 port map( A => n141, Z => n167);
   U40 : CLKBUF_X1 port map( A => n437, Z => n173);
   U41 : INV_X1 port map( A => SEL(1), ZN => n176);
   U42 : INV_X1 port map( A => SEL(2), ZN => n174);
   U43 : NAND3_X1 port map( A1 => SEL(0), A2 => n176, A3 => n174, ZN => n178);
   U44 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n174, ZN => n179)
                           ;
   U45 : INV_X1 port map( A => SEL(0), ZN => n177);
   U46 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n175);
   U47 : NAND2_X1 port map( A1 => E(0), A2 => n144, ZN => n185);
   U48 : INV_X1 port map( A => n178, ZN => n434);
   U49 : NAND2_X1 port map( A1 => B(0), A2 => n150, ZN => n184);
   U50 : INV_X1 port map( A => n179, ZN => n435);
   U51 : NAND2_X1 port map( A1 => D(0), A2 => n156, ZN => n183);
   U52 : INV_X1 port map( A => n180, ZN => n437);
   U53 : INV_X1 port map( A => n181, ZN => n436);
   U54 : AOI22_X1 port map( A1 => C(0), A2 => n168, B1 => A(0), B2 => n162, ZN 
                           => n182);
   U55 : NAND4_X1 port map( A1 => n185, A2 => n184, A3 => n183, A4 => n182, ZN 
                           => Y(0));
   U56 : NAND2_X1 port map( A1 => E(1), A2 => n144, ZN => n189);
   U57 : NAND2_X1 port map( A1 => B(1), A2 => n150, ZN => n188);
   U58 : NAND2_X1 port map( A1 => D(1), A2 => n156, ZN => n187);
   U59 : AOI22_X1 port map( A1 => C(1), A2 => n140, B1 => A(1), B2 => n162, ZN 
                           => n186);
   U60 : NAND4_X1 port map( A1 => n189, A2 => n188, A3 => n187, A4 => n186, ZN 
                           => Y(1));
   U61 : NAND2_X1 port map( A1 => E(2), A2 => n146, ZN => n193);
   U62 : NAND2_X1 port map( A1 => B(2), A2 => n150, ZN => n192);
   U63 : NAND2_X1 port map( A1 => D(2), A2 => n156, ZN => n191);
   U64 : AOI22_X1 port map( A1 => C(2), A2 => n139, B1 => A(2), B2 => n164, ZN 
                           => n190);
   U65 : NAND4_X1 port map( A1 => n193, A2 => n192, A3 => n191, A4 => n190, ZN 
                           => Y(2));
   U66 : NAND2_X1 port map( A1 => E(3), A2 => n145, ZN => n197);
   U67 : NAND2_X1 port map( A1 => B(3), A2 => n150, ZN => n196);
   U68 : NAND2_X1 port map( A1 => D(3), A2 => n156, ZN => n195);
   U69 : AOI22_X1 port map( A1 => C(3), A2 => n173, B1 => A(3), B2 => n163, ZN 
                           => n194);
   U70 : NAND4_X1 port map( A1 => n197, A2 => n196, A3 => n195, A4 => n194, ZN 
                           => Y(3));
   U71 : NAND2_X1 port map( A1 => E(4), A2 => n149, ZN => n201);
   U72 : NAND2_X1 port map( A1 => B(4), A2 => n150, ZN => n200);
   U73 : NAND2_X1 port map( A1 => D(4), A2 => n156, ZN => n199);
   U74 : AOI22_X1 port map( A1 => C(4), A2 => n172, B1 => A(4), B2 => n164, ZN 
                           => n198);
   U75 : NAND2_X1 port map( A1 => E(5), A2 => n148, ZN => n205);
   U76 : NAND2_X1 port map( A1 => B(5), A2 => n150, ZN => n204);
   U77 : NAND2_X1 port map( A1 => D(5), A2 => n156, ZN => n203);
   U78 : AOI22_X1 port map( A1 => C(5), A2 => n171, B1 => A(5), B2 => n163, ZN 
                           => n202);
   U79 : NAND4_X1 port map( A1 => n205, A2 => n204, A3 => n203, A4 => n202, ZN 
                           => Y(5));
   U80 : NAND2_X1 port map( A1 => E(6), A2 => n147, ZN => n209);
   U81 : NAND2_X1 port map( A1 => B(6), A2 => n150, ZN => n208);
   U82 : NAND2_X1 port map( A1 => D(6), A2 => n156, ZN => n207);
   U83 : AOI22_X1 port map( A1 => C(6), A2 => n170, B1 => A(6), B2 => n164, ZN 
                           => n206);
   U84 : NAND2_X1 port map( A1 => E(7), A2 => n146, ZN => n213);
   U85 : NAND2_X1 port map( A1 => B(7), A2 => n150, ZN => n212);
   U86 : NAND2_X1 port map( A1 => D(7), A2 => n156, ZN => n211);
   U87 : AOI22_X1 port map( A1 => C(7), A2 => n169, B1 => A(7), B2 => n163, ZN 
                           => n210);
   U88 : NAND2_X1 port map( A1 => E(8), A2 => n145, ZN => n217);
   U89 : NAND2_X1 port map( A1 => B(8), A2 => n150, ZN => n216);
   U90 : NAND2_X1 port map( A1 => D(8), A2 => n156, ZN => n215);
   U91 : AOI22_X1 port map( A1 => C(8), A2 => n173, B1 => A(8), B2 => n164, ZN 
                           => n214);
   U92 : NAND4_X1 port map( A1 => n217, A2 => n216, A3 => n215, A4 => n214, ZN 
                           => Y(8));
   U93 : NAND2_X1 port map( A1 => E(9), A2 => n149, ZN => n221);
   U94 : NAND2_X1 port map( A1 => B(9), A2 => n150, ZN => n220);
   U95 : NAND2_X1 port map( A1 => D(9), A2 => n156, ZN => n219);
   U96 : AOI22_X1 port map( A1 => C(9), A2 => n172, B1 => A(9), B2 => n163, ZN 
                           => n218);
   U97 : NAND4_X1 port map( A1 => n221, A2 => n220, A3 => n219, A4 => n218, ZN 
                           => Y(9));
   U98 : NAND2_X1 port map( A1 => E(10), A2 => n148, ZN => n225);
   U99 : NAND2_X1 port map( A1 => B(10), A2 => n150, ZN => n224);
   U100 : NAND2_X1 port map( A1 => D(10), A2 => n156, ZN => n223);
   U101 : AOI22_X1 port map( A1 => C(10), A2 => n171, B1 => A(10), B2 => n164, 
                           ZN => n222);
   U102 : NAND4_X1 port map( A1 => n225, A2 => n224, A3 => n223, A4 => n222, ZN
                           => Y(10));
   U103 : NAND2_X1 port map( A1 => E(11), A2 => n147, ZN => n229);
   U104 : NAND2_X1 port map( A1 => B(11), A2 => n150, ZN => n228);
   U105 : NAND2_X1 port map( A1 => D(11), A2 => n156, ZN => n227);
   U106 : AOI22_X1 port map( A1 => C(11), A2 => n170, B1 => A(11), B2 => n163, 
                           ZN => n226);
   U107 : NAND4_X1 port map( A1 => n229, A2 => n228, A3 => n227, A4 => n226, ZN
                           => Y(11));
   U108 : NAND2_X1 port map( A1 => E(12), A2 => n146, ZN => n233);
   U109 : NAND2_X1 port map( A1 => B(12), A2 => n151, ZN => n232);
   U110 : NAND2_X1 port map( A1 => D(12), A2 => n157, ZN => n231);
   U111 : AOI22_X1 port map( A1 => C(12), A2 => n169, B1 => A(12), B2 => n164, 
                           ZN => n230);
   U112 : NAND4_X1 port map( A1 => n233, A2 => n232, A3 => n231, A4 => n230, ZN
                           => Y(12));
   U113 : NAND2_X1 port map( A1 => E(13), A2 => n145, ZN => n237);
   U114 : NAND2_X1 port map( A1 => B(13), A2 => n151, ZN => n236);
   U115 : NAND2_X1 port map( A1 => D(13), A2 => n157, ZN => n235);
   U116 : AOI22_X1 port map( A1 => C(13), A2 => n140, B1 => A(13), B2 => n163, 
                           ZN => n234);
   U117 : NAND4_X1 port map( A1 => n237, A2 => n236, A3 => n235, A4 => n234, ZN
                           => Y(13));
   U118 : NAND2_X1 port map( A1 => E(14), A2 => n149, ZN => n241);
   U119 : NAND2_X1 port map( A1 => B(14), A2 => n151, ZN => n240);
   U120 : NAND2_X1 port map( A1 => D(14), A2 => n157, ZN => n239);
   U121 : AOI22_X1 port map( A1 => C(14), A2 => n139, B1 => A(14), B2 => n164, 
                           ZN => n238);
   U122 : NAND4_X1 port map( A1 => n241, A2 => n240, A3 => n239, A4 => n238, ZN
                           => Y(14));
   U123 : NAND2_X1 port map( A1 => E(15), A2 => n148, ZN => n245);
   U124 : NAND2_X1 port map( A1 => B(15), A2 => n151, ZN => n244);
   U125 : NAND2_X1 port map( A1 => D(15), A2 => n157, ZN => n243);
   U126 : AOI22_X1 port map( A1 => C(15), A2 => n140, B1 => A(15), B2 => n163, 
                           ZN => n242);
   U127 : NAND4_X1 port map( A1 => n245, A2 => n244, A3 => n243, A4 => n242, ZN
                           => Y(15));
   U128 : NAND2_X1 port map( A1 => E(16), A2 => n147, ZN => n249);
   U129 : NAND2_X1 port map( A1 => B(16), A2 => n151, ZN => n248);
   U130 : NAND2_X1 port map( A1 => D(16), A2 => n157, ZN => n247);
   U131 : AOI22_X1 port map( A1 => C(16), A2 => n139, B1 => A(16), B2 => n164, 
                           ZN => n246);
   U132 : NAND4_X1 port map( A1 => n249, A2 => n248, A3 => n247, A4 => n246, ZN
                           => Y(16));
   U133 : NAND2_X1 port map( A1 => E(17), A2 => n146, ZN => n253);
   U134 : NAND2_X1 port map( A1 => B(17), A2 => n151, ZN => n252);
   U135 : NAND2_X1 port map( A1 => D(17), A2 => n157, ZN => n251);
   U136 : AOI22_X1 port map( A1 => C(17), A2 => n173, B1 => A(17), B2 => n163, 
                           ZN => n250);
   U137 : NAND4_X1 port map( A1 => n253, A2 => n252, A3 => n251, A4 => n250, ZN
                           => Y(17));
   U138 : NAND2_X1 port map( A1 => E(18), A2 => n145, ZN => n257);
   U139 : NAND2_X1 port map( A1 => B(18), A2 => n151, ZN => n256);
   U140 : NAND2_X1 port map( A1 => D(18), A2 => n157, ZN => n255);
   U141 : AOI22_X1 port map( A1 => C(18), A2 => n172, B1 => A(18), B2 => n164, 
                           ZN => n254);
   U142 : NAND4_X1 port map( A1 => n257, A2 => n256, A3 => n255, A4 => n254, ZN
                           => Y(18));
   U143 : NAND2_X1 port map( A1 => E(19), A2 => n149, ZN => n261);
   U144 : NAND2_X1 port map( A1 => B(19), A2 => n151, ZN => n260);
   U145 : NAND2_X1 port map( A1 => D(19), A2 => n157, ZN => n259);
   U146 : AOI22_X1 port map( A1 => C(19), A2 => n171, B1 => A(19), B2 => n163, 
                           ZN => n258);
   U147 : NAND4_X1 port map( A1 => n261, A2 => n260, A3 => n259, A4 => n258, ZN
                           => Y(19));
   U148 : NAND2_X1 port map( A1 => E(20), A2 => n148, ZN => n265);
   U149 : NAND2_X1 port map( A1 => B(20), A2 => n151, ZN => n264);
   U150 : NAND2_X1 port map( A1 => D(20), A2 => n157, ZN => n263);
   U151 : AOI22_X1 port map( A1 => C(20), A2 => n170, B1 => A(20), B2 => n164, 
                           ZN => n262);
   U152 : NAND4_X1 port map( A1 => n265, A2 => n264, A3 => n263, A4 => n262, ZN
                           => Y(20));
   U153 : NAND2_X1 port map( A1 => E(21), A2 => n147, ZN => n269);
   U154 : NAND2_X1 port map( A1 => B(21), A2 => n151, ZN => n268);
   U155 : NAND2_X1 port map( A1 => D(21), A2 => n157, ZN => n267);
   U156 : AOI22_X1 port map( A1 => C(21), A2 => n169, B1 => A(21), B2 => n163, 
                           ZN => n266);
   U157 : NAND4_X1 port map( A1 => n269, A2 => n268, A3 => n267, A4 => n266, ZN
                           => Y(21));
   U158 : NAND2_X1 port map( A1 => E(22), A2 => n146, ZN => n273);
   U159 : NAND2_X1 port map( A1 => B(22), A2 => n151, ZN => n272);
   U160 : NAND2_X1 port map( A1 => D(22), A2 => n157, ZN => n271);
   U161 : AOI22_X1 port map( A1 => C(22), A2 => n140, B1 => A(22), B2 => n164, 
                           ZN => n270);
   U162 : NAND4_X1 port map( A1 => n273, A2 => n272, A3 => n271, A4 => n270, ZN
                           => Y(22));
   U163 : NAND2_X1 port map( A1 => E(23), A2 => n145, ZN => n277);
   U164 : NAND2_X1 port map( A1 => B(23), A2 => n151, ZN => n276);
   U165 : NAND2_X1 port map( A1 => D(23), A2 => n157, ZN => n275);
   U166 : AOI22_X1 port map( A1 => C(23), A2 => n140, B1 => A(23), B2 => n163, 
                           ZN => n274);
   U167 : NAND4_X1 port map( A1 => n277, A2 => n276, A3 => n275, A4 => n274, ZN
                           => Y(23));
   U168 : NAND2_X1 port map( A1 => E(24), A2 => n149, ZN => n281);
   U169 : NAND2_X1 port map( A1 => B(24), A2 => n152, ZN => n280);
   U170 : NAND2_X1 port map( A1 => D(24), A2 => n158, ZN => n279);
   U171 : AOI22_X1 port map( A1 => C(24), A2 => n140, B1 => A(24), B2 => n164, 
                           ZN => n278);
   U172 : NAND4_X1 port map( A1 => n281, A2 => n280, A3 => n279, A4 => n278, ZN
                           => Y(24));
   U173 : NAND2_X1 port map( A1 => E(25), A2 => n148, ZN => n285);
   U174 : NAND2_X1 port map( A1 => B(25), A2 => n152, ZN => n284);
   U175 : NAND2_X1 port map( A1 => D(25), A2 => n158, ZN => n283);
   U176 : AOI22_X1 port map( A1 => C(25), A2 => n139, B1 => A(25), B2 => n163, 
                           ZN => n282);
   U177 : NAND4_X1 port map( A1 => n285, A2 => n284, A3 => n283, A4 => n282, ZN
                           => Y(25));
   U178 : NAND2_X1 port map( A1 => E(26), A2 => n147, ZN => n289);
   U179 : NAND2_X1 port map( A1 => B(26), A2 => n152, ZN => n288);
   U180 : NAND2_X1 port map( A1 => D(26), A2 => n158, ZN => n287);
   U181 : AOI22_X1 port map( A1 => C(26), A2 => n139, B1 => A(26), B2 => n164, 
                           ZN => n286);
   U182 : NAND4_X1 port map( A1 => n289, A2 => n288, A3 => n287, A4 => n286, ZN
                           => Y(26));
   U183 : NAND2_X1 port map( A1 => E(27), A2 => n146, ZN => n293);
   U184 : NAND2_X1 port map( A1 => B(27), A2 => n152, ZN => n292);
   U185 : NAND2_X1 port map( A1 => D(27), A2 => n158, ZN => n291);
   U186 : AOI22_X1 port map( A1 => C(27), A2 => n139, B1 => A(27), B2 => n163, 
                           ZN => n290);
   U187 : NAND4_X1 port map( A1 => n293, A2 => n292, A3 => n291, A4 => n290, ZN
                           => Y(27));
   U188 : NAND2_X1 port map( A1 => E(28), A2 => n145, ZN => n297);
   U189 : NAND2_X1 port map( A1 => B(28), A2 => n152, ZN => n296);
   U190 : NAND2_X1 port map( A1 => D(28), A2 => n158, ZN => n295);
   U191 : AOI22_X1 port map( A1 => C(28), A2 => n140, B1 => A(28), B2 => n164, 
                           ZN => n294);
   U192 : NAND4_X1 port map( A1 => n297, A2 => n296, A3 => n295, A4 => n294, ZN
                           => Y(28));
   U193 : NAND2_X1 port map( A1 => E(29), A2 => n149, ZN => n301);
   U194 : NAND2_X1 port map( A1 => B(29), A2 => n152, ZN => n300);
   U195 : NAND2_X1 port map( A1 => D(29), A2 => n158, ZN => n299);
   U196 : AOI22_X1 port map( A1 => C(29), A2 => n139, B1 => A(29), B2 => n163, 
                           ZN => n298);
   U197 : NAND4_X1 port map( A1 => n301, A2 => n300, A3 => n299, A4 => n298, ZN
                           => Y(29));
   U198 : NAND2_X1 port map( A1 => E(30), A2 => n148, ZN => n305);
   U199 : NAND2_X1 port map( A1 => B(30), A2 => n152, ZN => n304);
   U200 : NAND2_X1 port map( A1 => D(30), A2 => n158, ZN => n303);
   U201 : AOI22_X1 port map( A1 => C(30), A2 => n140, B1 => A(30), B2 => n164, 
                           ZN => n302);
   U202 : NAND4_X1 port map( A1 => n305, A2 => n304, A3 => n303, A4 => n302, ZN
                           => Y(30));
   U203 : NAND2_X1 port map( A1 => E(31), A2 => n147, ZN => n309);
   U204 : NAND2_X1 port map( A1 => B(31), A2 => n152, ZN => n308);
   U205 : NAND2_X1 port map( A1 => D(31), A2 => n158, ZN => n307);
   U206 : AOI22_X1 port map( A1 => C(31), A2 => n139, B1 => A(31), B2 => n163, 
                           ZN => n306);
   U207 : NAND4_X1 port map( A1 => n309, A2 => n308, A3 => n307, A4 => n306, ZN
                           => Y(31));
   U208 : NAND2_X1 port map( A1 => E(32), A2 => n146, ZN => n313);
   U209 : NAND2_X1 port map( A1 => B(32), A2 => n152, ZN => n312);
   U210 : NAND2_X1 port map( A1 => D(32), A2 => n158, ZN => n311);
   U211 : AOI22_X1 port map( A1 => C(32), A2 => n173, B1 => A(32), B2 => n164, 
                           ZN => n310);
   U212 : NAND4_X1 port map( A1 => n313, A2 => n312, A3 => n311, A4 => n310, ZN
                           => Y(32));
   U213 : NAND2_X1 port map( A1 => E(33), A2 => n145, ZN => n317);
   U214 : NAND2_X1 port map( A1 => B(33), A2 => n152, ZN => n316);
   U215 : NAND2_X1 port map( A1 => D(33), A2 => n158, ZN => n315);
   U216 : AOI22_X1 port map( A1 => C(33), A2 => n172, B1 => A(33), B2 => n163, 
                           ZN => n314);
   U217 : NAND4_X1 port map( A1 => n317, A2 => n316, A3 => n315, A4 => n314, ZN
                           => Y(33));
   U218 : NAND2_X1 port map( A1 => E(34), A2 => n149, ZN => n321);
   U219 : NAND2_X1 port map( A1 => B(34), A2 => n152, ZN => n320);
   U220 : NAND2_X1 port map( A1 => D(34), A2 => n158, ZN => n319);
   U221 : AOI22_X1 port map( A1 => C(34), A2 => n171, B1 => A(34), B2 => n164, 
                           ZN => n318);
   U222 : NAND4_X1 port map( A1 => n321, A2 => n320, A3 => n319, A4 => n318, ZN
                           => Y(34));
   U223 : NAND2_X1 port map( A1 => E(35), A2 => n148, ZN => n325);
   U224 : NAND2_X1 port map( A1 => B(35), A2 => n152, ZN => n324);
   U225 : NAND2_X1 port map( A1 => D(35), A2 => n158, ZN => n323);
   U226 : AOI22_X1 port map( A1 => C(35), A2 => n170, B1 => A(35), B2 => n163, 
                           ZN => n322);
   U227 : NAND4_X1 port map( A1 => n325, A2 => n324, A3 => n323, A4 => n322, ZN
                           => Y(35));
   U228 : NAND2_X1 port map( A1 => E(36), A2 => n147, ZN => n329);
   U229 : NAND2_X1 port map( A1 => B(36), A2 => n153, ZN => n328);
   U230 : NAND2_X1 port map( A1 => D(36), A2 => n159, ZN => n327);
   U231 : AOI22_X1 port map( A1 => C(36), A2 => n169, B1 => A(36), B2 => n165, 
                           ZN => n326);
   U232 : NAND4_X1 port map( A1 => n329, A2 => n328, A3 => n327, A4 => n326, ZN
                           => Y(36));
   U233 : NAND2_X1 port map( A1 => E(37), A2 => n146, ZN => n333);
   U234 : NAND2_X1 port map( A1 => B(37), A2 => n153, ZN => n332);
   U235 : NAND2_X1 port map( A1 => D(37), A2 => n159, ZN => n331);
   U236 : AOI22_X1 port map( A1 => C(37), A2 => n140, B1 => A(37), B2 => n165, 
                           ZN => n330);
   U237 : NAND4_X1 port map( A1 => n333, A2 => n332, A3 => n331, A4 => n330, ZN
                           => Y(37));
   U238 : NAND2_X1 port map( A1 => E(38), A2 => n145, ZN => n337);
   U239 : NAND2_X1 port map( A1 => B(38), A2 => n153, ZN => n336);
   U240 : NAND2_X1 port map( A1 => D(38), A2 => n159, ZN => n335);
   U241 : AOI22_X1 port map( A1 => C(38), A2 => n139, B1 => A(38), B2 => n165, 
                           ZN => n334);
   U242 : NAND4_X1 port map( A1 => n337, A2 => n336, A3 => n335, A4 => n334, ZN
                           => Y(38));
   U243 : NAND2_X1 port map( A1 => E(39), A2 => n149, ZN => n341);
   U244 : NAND2_X1 port map( A1 => B(39), A2 => n153, ZN => n340);
   U245 : NAND2_X1 port map( A1 => D(39), A2 => n159, ZN => n339);
   U246 : AOI22_X1 port map( A1 => C(39), A2 => n140, B1 => A(39), B2 => n165, 
                           ZN => n338);
   U247 : NAND4_X1 port map( A1 => n341, A2 => n340, A3 => n339, A4 => n338, ZN
                           => Y(39));
   U248 : NAND2_X1 port map( A1 => E(40), A2 => n148, ZN => n345);
   U249 : NAND2_X1 port map( A1 => B(40), A2 => n153, ZN => n344);
   U250 : NAND2_X1 port map( A1 => D(40), A2 => n159, ZN => n343);
   U251 : AOI22_X1 port map( A1 => C(40), A2 => n139, B1 => A(40), B2 => n165, 
                           ZN => n342);
   U252 : NAND4_X1 port map( A1 => n345, A2 => n344, A3 => n343, A4 => n342, ZN
                           => Y(40));
   U253 : NAND2_X1 port map( A1 => E(41), A2 => n147, ZN => n349);
   U254 : NAND2_X1 port map( A1 => B(41), A2 => n153, ZN => n348);
   U255 : NAND2_X1 port map( A1 => D(41), A2 => n159, ZN => n347);
   U256 : AOI22_X1 port map( A1 => C(41), A2 => n173, B1 => A(41), B2 => n165, 
                           ZN => n346);
   U257 : NAND4_X1 port map( A1 => n349, A2 => n348, A3 => n347, A4 => n346, ZN
                           => Y(41));
   U258 : NAND2_X1 port map( A1 => E(42), A2 => n146, ZN => n353);
   U259 : NAND2_X1 port map( A1 => B(42), A2 => n153, ZN => n352);
   U260 : NAND2_X1 port map( A1 => D(42), A2 => n159, ZN => n351);
   U261 : AOI22_X1 port map( A1 => C(42), A2 => n172, B1 => A(42), B2 => n165, 
                           ZN => n350);
   U262 : NAND4_X1 port map( A1 => n353, A2 => n352, A3 => n351, A4 => n350, ZN
                           => Y(42));
   U263 : NAND2_X1 port map( A1 => E(43), A2 => n145, ZN => n357);
   U264 : NAND2_X1 port map( A1 => B(43), A2 => n153, ZN => n356);
   U265 : NAND2_X1 port map( A1 => D(43), A2 => n159, ZN => n355);
   U266 : AOI22_X1 port map( A1 => C(43), A2 => n171, B1 => A(43), B2 => n165, 
                           ZN => n354);
   U267 : NAND4_X1 port map( A1 => n357, A2 => n356, A3 => n355, A4 => n354, ZN
                           => Y(43));
   U268 : NAND2_X1 port map( A1 => E(44), A2 => n149, ZN => n361);
   U269 : NAND2_X1 port map( A1 => B(44), A2 => n153, ZN => n360);
   U270 : NAND2_X1 port map( A1 => D(44), A2 => n159, ZN => n359);
   U271 : AOI22_X1 port map( A1 => C(44), A2 => n170, B1 => A(44), B2 => n165, 
                           ZN => n358);
   U272 : NAND4_X1 port map( A1 => n361, A2 => n360, A3 => n359, A4 => n358, ZN
                           => Y(44));
   U273 : NAND2_X1 port map( A1 => E(45), A2 => n148, ZN => n365);
   U274 : NAND2_X1 port map( A1 => B(45), A2 => n153, ZN => n364);
   U275 : NAND2_X1 port map( A1 => D(45), A2 => n159, ZN => n363);
   U276 : AOI22_X1 port map( A1 => C(45), A2 => n169, B1 => A(45), B2 => n165, 
                           ZN => n362);
   U277 : NAND4_X1 port map( A1 => n365, A2 => n364, A3 => n363, A4 => n362, ZN
                           => Y(45));
   U278 : NAND2_X1 port map( A1 => E(46), A2 => n147, ZN => n369);
   U279 : NAND2_X1 port map( A1 => B(46), A2 => n153, ZN => n368);
   U280 : NAND2_X1 port map( A1 => D(46), A2 => n159, ZN => n367);
   U281 : AOI22_X1 port map( A1 => C(46), A2 => n140, B1 => A(46), B2 => n165, 
                           ZN => n366);
   U282 : NAND4_X1 port map( A1 => n369, A2 => n368, A3 => n367, A4 => n366, ZN
                           => Y(46));
   U283 : NAND2_X1 port map( A1 => E(47), A2 => n146, ZN => n373);
   U284 : NAND2_X1 port map( A1 => B(47), A2 => n153, ZN => n372);
   U285 : NAND2_X1 port map( A1 => D(47), A2 => n159, ZN => n371);
   U286 : AOI22_X1 port map( A1 => C(47), A2 => n139, B1 => A(47), B2 => n165, 
                           ZN => n370);
   U287 : NAND4_X1 port map( A1 => n373, A2 => n372, A3 => n371, A4 => n370, ZN
                           => Y(47));
   U288 : NAND2_X1 port map( A1 => E(48), A2 => n145, ZN => n377);
   U289 : NAND2_X1 port map( A1 => B(48), A2 => n154, ZN => n376);
   U290 : NAND2_X1 port map( A1 => D(48), A2 => n160, ZN => n375);
   U291 : AOI22_X1 port map( A1 => C(48), A2 => n140, B1 => A(48), B2 => n166, 
                           ZN => n374);
   U292 : NAND4_X1 port map( A1 => n377, A2 => n376, A3 => n375, A4 => n374, ZN
                           => Y(48));
   U293 : NAND2_X1 port map( A1 => E(49), A2 => n149, ZN => n381);
   U294 : NAND2_X1 port map( A1 => B(49), A2 => n154, ZN => n380);
   U295 : NAND2_X1 port map( A1 => D(49), A2 => n160, ZN => n379);
   U296 : AOI22_X1 port map( A1 => C(49), A2 => n139, B1 => A(49), B2 => n166, 
                           ZN => n378);
   U297 : NAND4_X1 port map( A1 => n381, A2 => n380, A3 => n379, A4 => n378, ZN
                           => Y(49));
   U298 : NAND2_X1 port map( A1 => E(50), A2 => n148, ZN => n385);
   U299 : NAND2_X1 port map( A1 => B(50), A2 => n154, ZN => n384);
   U300 : NAND2_X1 port map( A1 => D(50), A2 => n160, ZN => n383);
   U301 : AOI22_X1 port map( A1 => C(50), A2 => n140, B1 => A(50), B2 => n166, 
                           ZN => n382);
   U302 : NAND4_X1 port map( A1 => n385, A2 => n384, A3 => n383, A4 => n382, ZN
                           => Y(50));
   U303 : NAND2_X1 port map( A1 => E(51), A2 => n147, ZN => n389);
   U304 : NAND2_X1 port map( A1 => B(51), A2 => n154, ZN => n388);
   U305 : NAND2_X1 port map( A1 => D(51), A2 => n160, ZN => n387);
   U306 : AOI22_X1 port map( A1 => C(51), A2 => n139, B1 => A(51), B2 => n166, 
                           ZN => n386);
   U307 : NAND4_X1 port map( A1 => n389, A2 => n388, A3 => n387, A4 => n386, ZN
                           => Y(51));
   U308 : NAND2_X1 port map( A1 => E(52), A2 => n146, ZN => n393);
   U309 : NAND2_X1 port map( A1 => B(52), A2 => n154, ZN => n392);
   U310 : NAND2_X1 port map( A1 => D(52), A2 => n160, ZN => n391);
   U311 : AOI22_X1 port map( A1 => C(52), A2 => n173, B1 => A(52), B2 => n166, 
                           ZN => n390);
   U312 : NAND4_X1 port map( A1 => n393, A2 => n392, A3 => n391, A4 => n390, ZN
                           => Y(52));
   U313 : NAND2_X1 port map( A1 => E(53), A2 => n145, ZN => n397);
   U314 : NAND2_X1 port map( A1 => B(53), A2 => n154, ZN => n396);
   U315 : NAND2_X1 port map( A1 => D(53), A2 => n160, ZN => n395);
   U316 : AOI22_X1 port map( A1 => C(53), A2 => n172, B1 => A(53), B2 => n166, 
                           ZN => n394);
   U317 : NAND4_X1 port map( A1 => n397, A2 => n396, A3 => n395, A4 => n394, ZN
                           => Y(53));
   U318 : NAND2_X1 port map( A1 => E(54), A2 => n149, ZN => n401);
   U319 : NAND2_X1 port map( A1 => B(54), A2 => n154, ZN => n400);
   U320 : NAND2_X1 port map( A1 => D(54), A2 => n160, ZN => n399);
   U321 : AOI22_X1 port map( A1 => C(54), A2 => n171, B1 => A(54), B2 => n166, 
                           ZN => n398);
   U322 : NAND4_X1 port map( A1 => n401, A2 => n400, A3 => n399, A4 => n398, ZN
                           => Y(54));
   U323 : NAND2_X1 port map( A1 => E(55), A2 => n148, ZN => n405);
   U324 : NAND2_X1 port map( A1 => B(55), A2 => n154, ZN => n404);
   U325 : NAND2_X1 port map( A1 => D(55), A2 => n160, ZN => n403);
   U326 : AOI22_X1 port map( A1 => C(55), A2 => n170, B1 => A(55), B2 => n166, 
                           ZN => n402);
   U327 : NAND4_X1 port map( A1 => n405, A2 => n404, A3 => n403, A4 => n402, ZN
                           => Y(55));
   U328 : NAND2_X1 port map( A1 => E(56), A2 => n147, ZN => n409);
   U329 : NAND2_X1 port map( A1 => B(56), A2 => n154, ZN => n408);
   U330 : NAND2_X1 port map( A1 => D(56), A2 => n160, ZN => n407);
   U331 : AOI22_X1 port map( A1 => C(56), A2 => n169, B1 => A(56), B2 => n166, 
                           ZN => n406);
   U332 : NAND4_X1 port map( A1 => n409, A2 => n408, A3 => n407, A4 => n406, ZN
                           => Y(56));
   U333 : NAND2_X1 port map( A1 => E(57), A2 => n146, ZN => n413);
   U334 : NAND2_X1 port map( A1 => B(57), A2 => n154, ZN => n412);
   U335 : NAND2_X1 port map( A1 => D(57), A2 => n160, ZN => n411);
   U336 : AOI22_X1 port map( A1 => C(57), A2 => n173, B1 => A(57), B2 => n166, 
                           ZN => n410);
   U337 : NAND4_X1 port map( A1 => n413, A2 => n412, A3 => n411, A4 => n410, ZN
                           => Y(57));
   U338 : NAND2_X1 port map( A1 => E(58), A2 => n145, ZN => n417);
   U339 : NAND2_X1 port map( A1 => B(58), A2 => n154, ZN => n416);
   U340 : NAND2_X1 port map( A1 => D(58), A2 => n160, ZN => n415);
   U341 : AOI22_X1 port map( A1 => C(58), A2 => n172, B1 => A(58), B2 => n166, 
                           ZN => n414);
   U342 : NAND4_X1 port map( A1 => n417, A2 => n416, A3 => n415, A4 => n414, ZN
                           => Y(58));
   U343 : NAND2_X1 port map( A1 => E(59), A2 => n149, ZN => n421);
   U344 : NAND2_X1 port map( A1 => B(59), A2 => n154, ZN => n420);
   U345 : NAND2_X1 port map( A1 => D(59), A2 => n160, ZN => n419);
   U346 : AOI22_X1 port map( A1 => C(59), A2 => n171, B1 => A(59), B2 => n166, 
                           ZN => n418);
   U347 : NAND4_X1 port map( A1 => n421, A2 => n420, A3 => n419, A4 => n418, ZN
                           => Y(59));
   U348 : NAND2_X1 port map( A1 => E(60), A2 => n148, ZN => n425);
   U349 : NAND2_X1 port map( A1 => B(60), A2 => n155, ZN => n424);
   U350 : NAND2_X1 port map( A1 => D(60), A2 => n161, ZN => n423);
   U351 : AOI22_X1 port map( A1 => C(60), A2 => n170, B1 => A(60), B2 => n167, 
                           ZN => n422);
   U352 : NAND4_X1 port map( A1 => n425, A2 => n424, A3 => n423, A4 => n422, ZN
                           => Y(60));
   U353 : NAND2_X1 port map( A1 => E(61), A2 => n147, ZN => n429);
   U354 : NAND2_X1 port map( A1 => B(61), A2 => n155, ZN => n428);
   U355 : NAND2_X1 port map( A1 => D(61), A2 => n161, ZN => n427);
   U356 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n167, 
                           ZN => n426);
   U357 : NAND4_X1 port map( A1 => n429, A2 => n428, A3 => n427, A4 => n426, ZN
                           => Y(61));
   U358 : NAND2_X1 port map( A1 => E(62), A2 => n146, ZN => n433);
   U359 : NAND2_X1 port map( A1 => B(62), A2 => n155, ZN => n432);
   U360 : NAND2_X1 port map( A1 => D(62), A2 => n161, ZN => n431);
   U361 : AOI22_X1 port map( A1 => C(62), A2 => n140, B1 => A(62), B2 => n167, 
                           ZN => n430);
   U362 : NAND4_X1 port map( A1 => n433, A2 => n432, A3 => n431, A4 => n430, ZN
                           => Y(62));
   U363 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n441);
   U364 : NAND2_X1 port map( A1 => B(63), A2 => n155, ZN => n440);
   U365 : NAND2_X1 port map( A1 => D(63), A2 => n161, ZN => n439);
   U366 : AOI22_X1 port map( A1 => C(63), A2 => n139, B1 => A(63), B2 => n167, 
                           ZN => n438);
   U367 : NAND4_X1 port map( A1 => n441, A2 => n440, A3 => n439, A4 => n438, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_13 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_13;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_13 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U2 : NAND4_X2 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U3 : NAND4_X2 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN 
                           => Y(11));
   U4 : NAND4_X2 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U5 : NAND4_X2 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U6 : BUF_X2 port map( A => n434, Z => n164);
   U7 : CLKBUF_X1 port map( A => n434, Z => n165);
   U8 : BUF_X2 port map( A => n432, Z => n152);
   U9 : BUF_X2 port map( A => n431, Z => n146);
   U10 : BUF_X2 port map( A => n139, Z => n140);
   U11 : CLKBUF_X1 port map( A => n139, Z => n141);
   U12 : BUF_X2 port map( A => n433, Z => n158);
   U13 : CLKBUF_X1 port map( A => n434, Z => n166);
   U14 : CLKBUF_X1 port map( A => n432, Z => n153);
   U15 : CLKBUF_X1 port map( A => n432, Z => n154);
   U16 : CLKBUF_X1 port map( A => n431, Z => n147);
   U17 : CLKBUF_X1 port map( A => n431, Z => n148);
   U18 : CLKBUF_X1 port map( A => n139, Z => n142);
   U19 : CLKBUF_X1 port map( A => n433, Z => n159);
   U20 : CLKBUF_X1 port map( A => n433, Z => n160);
   U21 : CLKBUF_X1 port map( A => n434, Z => n167);
   U22 : CLKBUF_X1 port map( A => n432, Z => n155);
   U23 : CLKBUF_X1 port map( A => n431, Z => n149);
   U24 : CLKBUF_X1 port map( A => n139, Z => n143);
   U25 : CLKBUF_X1 port map( A => n433, Z => n161);
   U26 : CLKBUF_X1 port map( A => n434, Z => n168);
   U27 : CLKBUF_X1 port map( A => n432, Z => n156);
   U28 : CLKBUF_X1 port map( A => n431, Z => n150);
   U29 : CLKBUF_X1 port map( A => n139, Z => n144);
   U30 : CLKBUF_X1 port map( A => n433, Z => n162);
   U31 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U32 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U33 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U34 : CLKBUF_X1 port map( A => n139, Z => n145);
   U35 : CLKBUF_X1 port map( A => n431, Z => n151);
   U36 : CLKBUF_X1 port map( A => n432, Z => n157);
   U37 : CLKBUF_X1 port map( A => n433, Z => n163);
   U38 : CLKBUF_X1 port map( A => n434, Z => n169);
   U39 : INV_X1 port map( A => SEL(1), ZN => n172);
   U40 : INV_X1 port map( A => SEL(2), ZN => n170);
   U41 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U42 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U43 : INV_X1 port map( A => SEL(0), ZN => n174);
   U44 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U45 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U46 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U47 : INV_X1 port map( A => n175, ZN => n431);
   U48 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U49 : INV_X1 port map( A => n176, ZN => n432);
   U50 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U51 : INV_X1 port map( A => n177, ZN => n434);
   U52 : INV_X1 port map( A => n178, ZN => n433);
   U53 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U54 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U55 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U56 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U57 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U58 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U59 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U60 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U61 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U62 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U63 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U64 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U65 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U66 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U67 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U68 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U69 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U70 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U71 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U72 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U73 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U74 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U75 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U76 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U77 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U78 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U79 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U80 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U81 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U82 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U83 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U84 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U85 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U86 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U87 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U88 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U89 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U90 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U91 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U92 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U93 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U94 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U95 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U96 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U97 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U98 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U99 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U100 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(10));
   U101 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U102 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U103 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U104 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U105 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U106 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U107 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U108 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U109 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U110 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U111 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U112 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U113 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U114 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U115 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U116 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U117 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U118 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U119 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U120 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U121 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U122 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U123 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U124 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U125 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U126 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U127 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U128 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U129 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U130 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U131 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U132 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U133 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U134 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U135 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U136 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U137 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U138 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U139 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U140 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U141 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U142 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U143 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U144 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U145 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U146 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U147 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U148 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U149 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U150 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U151 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U152 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U153 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U154 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U155 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U156 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U157 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U158 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U159 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U160 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U161 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U162 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U163 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U164 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U165 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U166 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U167 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U168 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U169 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U170 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U171 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U172 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U173 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U174 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U175 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U176 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U177 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U178 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U179 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U180 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U181 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U182 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U183 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U184 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U185 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U186 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U187 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U188 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U189 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U190 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U191 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U192 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U193 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U194 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U195 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U196 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U197 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U198 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U199 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U200 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U201 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U202 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U203 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U204 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U205 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U206 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U207 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U208 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U209 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U210 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U211 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U212 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U213 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U214 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U215 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U216 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U217 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U218 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U219 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U220 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U221 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U222 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U223 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U224 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U225 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U226 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U227 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U228 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U229 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U230 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U231 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U232 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U233 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U234 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U235 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U236 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U237 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U238 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U239 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U240 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U241 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U242 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U243 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U244 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U245 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U246 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U247 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U248 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U249 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U250 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U251 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U252 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U253 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U254 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U255 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U256 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U257 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U258 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U259 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U260 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U261 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U262 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U263 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U264 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U265 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U266 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U267 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U268 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U269 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U270 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U271 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U272 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U273 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U274 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U275 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U276 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U277 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U278 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U279 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U280 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U281 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U282 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U283 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U284 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U285 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U286 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U287 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U288 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U289 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U290 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U291 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U292 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U293 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U294 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U295 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U296 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U297 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U298 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U299 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U300 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U301 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U302 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U303 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U304 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U305 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U306 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U307 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U308 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U309 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U310 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U311 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U312 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U313 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U314 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U315 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U316 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U317 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U318 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U319 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U320 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U321 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U322 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U323 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U324 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U325 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U326 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U327 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U328 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U329 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U330 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U331 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U332 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U333 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U334 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U335 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U336 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U337 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U338 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U339 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U340 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U341 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U342 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U343 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U344 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U345 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U346 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U347 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U348 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U349 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U350 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U351 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U352 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U353 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U354 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => Y(61));
   U355 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U356 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U357 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U358 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U359 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => Y(62));
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_12 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_12;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_12 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X2 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U2 : NAND4_X2 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U3 : BUF_X1 port map( A => n434, Z => n164);
   U4 : BUF_X1 port map( A => n432, Z => n152);
   U5 : BUF_X1 port map( A => n431, Z => n146);
   U6 : BUF_X1 port map( A => n139, Z => n140);
   U7 : BUF_X1 port map( A => n433, Z => n158);
   U8 : CLKBUF_X1 port map( A => n434, Z => n165);
   U9 : CLKBUF_X1 port map( A => n434, Z => n166);
   U10 : CLKBUF_X1 port map( A => n432, Z => n153);
   U11 : CLKBUF_X1 port map( A => n432, Z => n154);
   U12 : CLKBUF_X1 port map( A => n431, Z => n147);
   U13 : CLKBUF_X1 port map( A => n431, Z => n148);
   U14 : CLKBUF_X1 port map( A => n139, Z => n141);
   U15 : CLKBUF_X1 port map( A => n139, Z => n142);
   U16 : CLKBUF_X1 port map( A => n433, Z => n159);
   U17 : CLKBUF_X1 port map( A => n433, Z => n160);
   U18 : CLKBUF_X1 port map( A => n434, Z => n167);
   U19 : CLKBUF_X1 port map( A => n432, Z => n155);
   U20 : CLKBUF_X1 port map( A => n431, Z => n149);
   U21 : CLKBUF_X1 port map( A => n139, Z => n143);
   U22 : CLKBUF_X1 port map( A => n433, Z => n161);
   U23 : CLKBUF_X1 port map( A => n434, Z => n168);
   U24 : CLKBUF_X1 port map( A => n432, Z => n156);
   U25 : CLKBUF_X1 port map( A => n431, Z => n150);
   U26 : CLKBUF_X1 port map( A => n139, Z => n144);
   U27 : CLKBUF_X1 port map( A => n433, Z => n162);
   U28 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U29 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U30 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U31 : CLKBUF_X1 port map( A => n139, Z => n145);
   U32 : CLKBUF_X1 port map( A => n431, Z => n151);
   U33 : CLKBUF_X1 port map( A => n432, Z => n157);
   U34 : CLKBUF_X1 port map( A => n433, Z => n163);
   U35 : CLKBUF_X1 port map( A => n434, Z => n169);
   U36 : INV_X1 port map( A => SEL(1), ZN => n172);
   U37 : INV_X1 port map( A => SEL(2), ZN => n170);
   U38 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U39 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U40 : INV_X1 port map( A => SEL(0), ZN => n174);
   U41 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U42 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U43 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U44 : INV_X1 port map( A => n175, ZN => n431);
   U45 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U46 : INV_X1 port map( A => n176, ZN => n432);
   U47 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U48 : INV_X1 port map( A => n177, ZN => n434);
   U49 : INV_X1 port map( A => n178, ZN => n433);
   U50 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U51 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U52 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U53 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U54 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U55 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U56 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U57 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U58 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U59 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U60 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U61 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U62 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U63 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U64 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U65 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U66 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U67 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U68 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U69 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U70 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U71 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U72 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U73 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U74 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U75 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U76 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U77 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U78 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U79 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U80 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U81 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U82 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U83 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U84 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U85 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U86 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U87 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U88 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U89 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U90 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U91 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U92 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U93 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U94 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U95 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U96 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U97 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U98 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U99 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN 
                           => Y(10));
   U100 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U101 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U102 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U103 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U104 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN
                           => Y(11));
   U105 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U106 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U107 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U108 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U109 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U110 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U111 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U112 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U113 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U114 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U115 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U116 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U117 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U118 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U119 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U120 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U121 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U122 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U123 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U124 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U125 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U126 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U127 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U128 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U129 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U130 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U131 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U132 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U133 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U134 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U135 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U136 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U137 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U138 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U139 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U140 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U141 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U142 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U143 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U144 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U145 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U146 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U147 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U148 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U149 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U150 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U151 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U152 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U153 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U154 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U155 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U156 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U157 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U158 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U159 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U160 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U161 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U162 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U163 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U164 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U165 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U166 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U167 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U168 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U169 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U170 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U171 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U172 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U173 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U174 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U175 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U176 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U177 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U178 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U179 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U180 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U181 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U182 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U183 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U184 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U185 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U186 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U187 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U188 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U189 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U190 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U191 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U192 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U193 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U194 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U195 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U196 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U197 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U198 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U199 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U200 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U201 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U202 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U203 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U204 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U205 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U206 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U207 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U208 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U209 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U210 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U211 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U212 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U213 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U214 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U215 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U216 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U217 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U218 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U219 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U220 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U221 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U222 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U223 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U224 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U225 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U226 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U227 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U228 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U229 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U230 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U231 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U232 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U233 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U234 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U235 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U236 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U237 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U238 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U239 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U240 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U241 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U242 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U243 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U244 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U245 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U246 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U247 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U248 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U249 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U250 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U251 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U252 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U253 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U254 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U255 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U256 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U257 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U258 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U259 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U260 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U261 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U262 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U263 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U264 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U265 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U266 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U267 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U268 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U269 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U270 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U271 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U272 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U273 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U274 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U275 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U276 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U277 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U278 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U279 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U280 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U281 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U282 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U283 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U284 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U285 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U286 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U287 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U288 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U289 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U290 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U291 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U292 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U293 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U294 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U295 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U296 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U297 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U298 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U299 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U300 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U301 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U302 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U303 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U304 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U305 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U306 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U307 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U308 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U309 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U310 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U311 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U312 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U313 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U314 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U315 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U316 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U317 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U318 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U319 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U320 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U321 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U322 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U323 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U324 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U325 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U326 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U327 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U328 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U329 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U330 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U331 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U332 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U333 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U334 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U335 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U336 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U337 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U338 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U339 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U340 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U341 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U342 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U343 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U344 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U345 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U346 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U347 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U348 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U349 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U350 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U351 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U352 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U353 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U354 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => Y(61));
   U355 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U356 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U357 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U358 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U359 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => Y(62));
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_11 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_11;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_11 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X2 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U2 : NAND4_X2 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN 
                           => Y(10));
   U3 : NAND4_X2 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U4 : NAND4_X2 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U5 : BUF_X2 port map( A => n434, Z => n164);
   U6 : BUF_X2 port map( A => n432, Z => n152);
   U7 : BUF_X1 port map( A => n431, Z => n146);
   U8 : BUF_X1 port map( A => n139, Z => n140);
   U9 : BUF_X1 port map( A => n433, Z => n158);
   U10 : CLKBUF_X1 port map( A => n434, Z => n165);
   U11 : CLKBUF_X1 port map( A => n432, Z => n153);
   U12 : CLKBUF_X1 port map( A => n431, Z => n147);
   U13 : CLKBUF_X1 port map( A => n139, Z => n141);
   U14 : CLKBUF_X1 port map( A => n433, Z => n159);
   U15 : CLKBUF_X1 port map( A => n434, Z => n167);
   U16 : CLKBUF_X1 port map( A => n434, Z => n166);
   U17 : CLKBUF_X1 port map( A => n432, Z => n155);
   U18 : CLKBUF_X1 port map( A => n432, Z => n154);
   U19 : CLKBUF_X1 port map( A => n431, Z => n149);
   U20 : CLKBUF_X1 port map( A => n431, Z => n148);
   U21 : CLKBUF_X1 port map( A => n139, Z => n143);
   U22 : CLKBUF_X1 port map( A => n139, Z => n142);
   U23 : CLKBUF_X1 port map( A => n433, Z => n161);
   U24 : CLKBUF_X1 port map( A => n433, Z => n160);
   U25 : CLKBUF_X1 port map( A => n434, Z => n168);
   U26 : CLKBUF_X1 port map( A => n432, Z => n156);
   U27 : CLKBUF_X1 port map( A => n431, Z => n150);
   U28 : CLKBUF_X1 port map( A => n139, Z => n144);
   U29 : CLKBUF_X1 port map( A => n433, Z => n162);
   U30 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U31 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U32 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U33 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U34 : CLKBUF_X1 port map( A => n139, Z => n145);
   U35 : CLKBUF_X1 port map( A => n431, Z => n151);
   U36 : CLKBUF_X1 port map( A => n432, Z => n157);
   U37 : CLKBUF_X1 port map( A => n433, Z => n163);
   U38 : CLKBUF_X1 port map( A => n434, Z => n169);
   U39 : INV_X1 port map( A => SEL(1), ZN => n172);
   U40 : INV_X1 port map( A => SEL(2), ZN => n170);
   U41 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U42 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U43 : INV_X1 port map( A => SEL(0), ZN => n174);
   U44 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U45 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U46 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U47 : INV_X1 port map( A => n175, ZN => n431);
   U48 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U49 : INV_X1 port map( A => n176, ZN => n432);
   U50 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U51 : INV_X1 port map( A => n177, ZN => n434);
   U52 : INV_X1 port map( A => n178, ZN => n433);
   U53 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U54 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U55 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U56 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U57 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U58 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U59 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U60 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U61 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U62 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U63 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U64 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U65 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U66 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U67 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U68 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U69 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U70 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U71 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U72 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U73 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U74 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U75 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U76 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U77 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U78 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U79 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U80 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U81 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U82 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U83 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U84 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U85 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U86 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U87 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U88 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U89 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U90 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U91 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U92 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U93 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U94 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U95 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U96 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U97 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U98 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U99 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U100 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U101 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U102 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U103 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U104 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN
                           => Y(11));
   U105 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U106 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U107 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U108 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U109 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U110 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U111 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U112 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U113 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U114 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U115 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U116 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U117 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U118 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U119 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U120 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U121 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U122 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U123 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U124 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U125 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U126 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U127 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U128 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U129 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U130 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U131 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U132 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U133 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U134 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U135 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U136 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U137 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U138 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U139 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U140 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U141 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U142 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U143 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U144 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U145 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U146 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U147 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U148 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U149 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U150 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U151 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U152 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U153 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U154 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U155 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U156 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U157 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U158 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U159 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U160 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U161 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U162 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U163 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U164 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U165 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U166 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U167 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U168 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U169 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U170 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U171 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U172 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U173 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U174 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U175 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U176 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U177 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U178 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U179 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U180 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U181 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U182 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U183 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U184 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U185 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U186 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U187 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U188 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U189 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U190 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U191 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U192 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U193 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U194 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U195 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U196 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U197 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U198 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U199 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U200 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U201 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U202 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U203 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U204 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U205 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U206 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U207 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U208 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U209 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U210 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U211 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U212 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U213 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U214 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U215 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U216 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U217 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U218 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U219 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U220 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U221 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U222 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U223 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U224 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U225 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U226 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U227 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U228 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U229 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U230 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U231 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U232 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U233 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U234 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U235 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U236 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U237 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U238 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U239 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U240 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U241 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U242 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U243 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U244 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U245 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U246 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U247 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U248 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U249 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U250 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U251 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U252 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U253 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U254 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U255 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U256 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U257 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U258 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U259 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U260 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U261 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U262 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U263 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U264 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U265 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U266 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U267 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U268 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U269 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U270 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U271 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U272 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U273 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U274 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U275 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U276 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U277 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U278 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U279 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U280 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U281 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U282 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U283 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U284 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U285 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U286 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U287 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U288 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U289 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U290 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U291 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U292 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U293 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U294 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U295 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U296 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U297 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U298 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U299 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U300 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U301 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U302 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U303 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U304 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U305 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U306 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U307 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U308 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U309 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U310 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U311 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U312 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U313 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U314 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U315 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U316 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U317 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U318 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U319 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U320 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U321 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U322 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U323 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U324 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U325 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U326 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U327 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U328 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U329 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U330 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U331 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U332 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U333 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U334 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U335 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U336 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U337 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U338 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U339 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U340 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U341 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U342 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U343 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U344 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U345 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U346 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U347 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U348 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U349 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U350 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U351 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U352 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U353 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U354 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => Y(61));
   U355 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U356 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U357 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U358 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U359 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => Y(62));
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_10 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_10;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_10 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X2 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U2 : NAND4_X2 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN 
                           => Y(60));
   U3 : BUF_X2 port map( A => n431, Z => n146);
   U4 : BUF_X2 port map( A => n434, Z => n164);
   U5 : BUF_X2 port map( A => n432, Z => n152);
   U6 : BUF_X1 port map( A => n139, Z => n140);
   U7 : BUF_X1 port map( A => n433, Z => n158);
   U8 : CLKBUF_X1 port map( A => n434, Z => n165);
   U9 : CLKBUF_X1 port map( A => n432, Z => n153);
   U10 : CLKBUF_X1 port map( A => n431, Z => n147);
   U11 : CLKBUF_X1 port map( A => n139, Z => n141);
   U12 : CLKBUF_X1 port map( A => n433, Z => n159);
   U13 : CLKBUF_X1 port map( A => n434, Z => n166);
   U14 : CLKBUF_X1 port map( A => n432, Z => n154);
   U15 : CLKBUF_X1 port map( A => n431, Z => n148);
   U16 : CLKBUF_X1 port map( A => n139, Z => n143);
   U17 : CLKBUF_X1 port map( A => n139, Z => n142);
   U18 : CLKBUF_X1 port map( A => n433, Z => n160);
   U19 : CLKBUF_X1 port map( A => n434, Z => n168);
   U20 : CLKBUF_X1 port map( A => n434, Z => n167);
   U21 : CLKBUF_X1 port map( A => n432, Z => n156);
   U22 : CLKBUF_X1 port map( A => n432, Z => n155);
   U23 : CLKBUF_X1 port map( A => n431, Z => n150);
   U24 : CLKBUF_X1 port map( A => n431, Z => n149);
   U25 : CLKBUF_X1 port map( A => n139, Z => n144);
   U26 : CLKBUF_X1 port map( A => n433, Z => n162);
   U27 : CLKBUF_X1 port map( A => n433, Z => n161);
   U28 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U29 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U30 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U31 : CLKBUF_X1 port map( A => n139, Z => n145);
   U32 : CLKBUF_X1 port map( A => n431, Z => n151);
   U33 : CLKBUF_X1 port map( A => n432, Z => n157);
   U34 : CLKBUF_X1 port map( A => n433, Z => n163);
   U35 : CLKBUF_X1 port map( A => n434, Z => n169);
   U36 : INV_X1 port map( A => SEL(1), ZN => n172);
   U37 : INV_X1 port map( A => SEL(2), ZN => n170);
   U38 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U39 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U40 : INV_X1 port map( A => SEL(0), ZN => n174);
   U41 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U42 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U43 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U44 : INV_X1 port map( A => n175, ZN => n431);
   U45 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U46 : INV_X1 port map( A => n176, ZN => n432);
   U47 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U48 : INV_X1 port map( A => n177, ZN => n434);
   U49 : INV_X1 port map( A => n178, ZN => n433);
   U50 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U51 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U52 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U53 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U54 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U55 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U56 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U57 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U58 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U59 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U60 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U61 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U62 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U63 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U64 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U65 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U66 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U67 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U68 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U69 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U70 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U71 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U72 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U73 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U74 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U75 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U76 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U77 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U78 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U79 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U80 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U81 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U82 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U83 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U84 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U85 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U86 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U87 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U88 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U89 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U90 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U91 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U92 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U93 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U94 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U95 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U96 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U97 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U98 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U99 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U100 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(10));
   U101 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U102 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U103 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U104 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U105 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN
                           => Y(11));
   U106 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U107 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U108 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U109 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U110 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U111 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U112 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U113 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U114 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U115 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U116 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U117 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U118 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U119 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U120 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U121 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U122 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U123 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U124 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U125 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U126 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U127 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U128 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U129 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U130 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U131 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U132 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U133 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U134 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U135 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U136 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U138 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U139 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U140 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U141 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U142 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U143 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U144 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U145 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U146 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U147 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U148 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U149 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U150 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U151 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U152 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U153 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U154 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U155 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U156 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U157 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U158 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U159 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U160 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U161 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U162 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U163 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U164 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U165 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U166 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U167 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U168 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U169 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U170 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U171 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U172 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U173 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U174 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U175 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U176 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U177 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U178 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U179 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U180 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U181 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U182 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U183 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U184 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U185 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U186 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U187 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U188 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U189 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U190 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U191 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U192 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U193 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U194 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U195 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U196 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U197 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U198 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U199 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U200 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U201 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U202 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U203 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U204 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U205 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U206 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U207 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U208 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U209 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U210 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U211 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U212 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U213 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U214 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U215 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U216 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U217 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U218 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U219 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U220 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U221 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U222 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U223 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U224 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U225 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U226 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U227 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U228 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U229 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U230 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U231 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U232 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U233 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U234 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U235 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U236 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U237 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U238 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U239 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U240 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U241 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U242 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U243 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U244 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U245 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U246 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U247 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U248 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U249 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U250 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U251 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U252 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U253 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U254 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U255 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U256 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U257 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U258 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U259 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U260 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U261 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U262 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U263 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U264 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U265 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U266 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U267 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U268 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U269 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U270 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U271 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U272 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U273 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U274 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U275 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U276 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U277 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U278 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U279 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U280 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U281 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U282 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U283 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U284 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U285 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U286 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U287 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U288 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U289 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U290 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U291 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U292 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U293 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U294 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U295 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U296 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U297 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U298 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U299 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U300 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U301 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U302 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U303 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U304 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U305 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U306 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U307 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U308 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U309 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U310 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U311 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U312 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U313 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U314 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U315 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U316 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U317 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U318 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U319 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U320 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U321 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U322 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U323 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U324 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U325 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U326 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U327 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U328 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U329 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U330 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U331 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U332 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U333 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U334 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U335 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U336 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U337 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U338 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U339 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U340 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U341 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U342 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U343 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U344 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U345 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U346 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U347 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U348 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U349 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U350 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U351 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U352 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U353 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U354 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => Y(61));
   U355 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U356 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U357 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U358 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U359 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => Y(62));
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_9 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_9;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_9 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X2 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN 
                           => Y(62));
   U2 : NAND4_X2 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U3 : NAND4_X2 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U4 : NAND4_X2 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN 
                           => Y(11));
   U5 : NAND4_X2 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U6 : BUF_X2 port map( A => n434, Z => n164);
   U7 : BUF_X2 port map( A => n432, Z => n152);
   U8 : BUF_X2 port map( A => n431, Z => n146);
   U9 : BUF_X2 port map( A => n139, Z => n140);
   U10 : BUF_X2 port map( A => n433, Z => n158);
   U11 : CLKBUF_X1 port map( A => n434, Z => n165);
   U12 : CLKBUF_X1 port map( A => n432, Z => n153);
   U13 : CLKBUF_X1 port map( A => n431, Z => n147);
   U14 : CLKBUF_X1 port map( A => n139, Z => n141);
   U15 : CLKBUF_X1 port map( A => n433, Z => n159);
   U16 : CLKBUF_X1 port map( A => n434, Z => n166);
   U17 : CLKBUF_X1 port map( A => n432, Z => n154);
   U18 : CLKBUF_X1 port map( A => n431, Z => n148);
   U19 : CLKBUF_X1 port map( A => n139, Z => n142);
   U20 : CLKBUF_X1 port map( A => n433, Z => n160);
   U21 : CLKBUF_X1 port map( A => n434, Z => n168);
   U22 : CLKBUF_X1 port map( A => n434, Z => n167);
   U23 : CLKBUF_X1 port map( A => n432, Z => n155);
   U24 : CLKBUF_X1 port map( A => n431, Z => n149);
   U25 : CLKBUF_X1 port map( A => n139, Z => n144);
   U26 : CLKBUF_X1 port map( A => n139, Z => n143);
   U27 : CLKBUF_X1 port map( A => n433, Z => n162);
   U28 : CLKBUF_X1 port map( A => n433, Z => n161);
   U29 : CLKBUF_X1 port map( A => n432, Z => n156);
   U30 : CLKBUF_X1 port map( A => n431, Z => n150);
   U31 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U32 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U33 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U34 : CLKBUF_X1 port map( A => n139, Z => n145);
   U35 : CLKBUF_X1 port map( A => n431, Z => n151);
   U36 : CLKBUF_X1 port map( A => n432, Z => n157);
   U37 : CLKBUF_X1 port map( A => n433, Z => n163);
   U38 : CLKBUF_X1 port map( A => n434, Z => n169);
   U39 : INV_X1 port map( A => SEL(1), ZN => n172);
   U40 : INV_X1 port map( A => SEL(2), ZN => n170);
   U41 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U42 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U43 : INV_X1 port map( A => SEL(0), ZN => n174);
   U44 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U45 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U46 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U47 : INV_X1 port map( A => n175, ZN => n431);
   U48 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U49 : INV_X1 port map( A => n176, ZN => n432);
   U50 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U51 : INV_X1 port map( A => n177, ZN => n434);
   U52 : INV_X1 port map( A => n178, ZN => n433);
   U53 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U54 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U55 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U56 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U57 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U58 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U59 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U60 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U61 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U62 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U63 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U64 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U65 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U66 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U67 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U68 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U69 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U70 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U71 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U72 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U73 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U74 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U75 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U76 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U77 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U78 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U79 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U80 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U81 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U82 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U83 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U84 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U85 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U86 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U87 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U88 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U89 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U90 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U91 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U92 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U93 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U94 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U95 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U96 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U97 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U98 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U99 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U100 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U101 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(10));
   U102 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U103 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U104 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U105 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U106 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U107 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U108 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U109 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U110 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U111 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U112 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U113 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U114 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U115 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U116 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U117 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U118 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U119 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U120 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U121 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U122 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U123 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U124 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U125 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U126 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U127 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U128 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U129 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U130 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U131 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U132 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U133 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U134 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U135 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U136 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U138 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U139 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U140 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U141 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U142 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U143 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U144 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U145 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U146 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U147 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U148 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U149 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U150 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U151 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U152 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U153 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U154 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U155 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U156 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U157 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U158 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U159 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U160 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U161 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U162 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U163 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U164 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U165 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U166 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U167 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U168 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U169 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U170 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U171 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U172 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U173 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U174 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U175 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U176 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U177 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U178 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U179 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U180 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U181 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U182 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U183 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U184 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U185 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U186 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U187 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U188 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U189 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U190 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U191 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U192 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U193 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U194 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U195 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U196 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U197 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U198 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U199 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U200 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U201 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U202 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U203 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U204 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U205 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U206 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U207 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U208 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U209 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U210 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U211 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U212 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U213 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U214 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U215 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U216 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U217 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U218 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U219 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U220 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U221 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U222 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U223 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U224 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U225 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U226 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U227 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U228 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U229 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U230 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U231 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U232 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U233 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U234 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U235 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U236 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U237 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U238 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U239 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U240 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U241 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U242 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U243 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U244 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U245 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U246 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U247 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U248 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U249 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U250 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U251 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U252 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U253 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U254 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U255 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U256 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U257 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U258 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U259 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U260 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U261 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U262 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U263 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U264 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U265 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U266 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U267 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U268 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U269 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U270 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U271 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U272 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U273 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U274 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U275 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U276 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U277 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U278 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U279 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U280 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U281 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U282 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U283 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U284 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U285 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U286 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U287 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U288 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U289 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U290 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U291 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U292 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U293 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U294 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U295 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U296 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U297 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U298 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U299 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U300 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U301 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U302 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U303 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U304 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U305 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U306 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U307 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U308 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U309 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U310 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U311 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U312 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U313 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U314 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U315 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U316 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U317 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U318 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U319 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U320 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U321 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U322 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U323 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U324 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U325 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U326 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U327 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U328 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U329 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U330 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U331 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U332 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U333 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U334 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U335 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U336 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U337 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U338 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U339 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U340 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U341 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U342 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U343 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U344 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U345 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U346 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U347 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U348 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U349 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U350 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U351 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U352 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U353 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U354 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U355 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => Y(61));
   U356 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U357 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U358 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U359 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_8 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_8;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_8 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN =>
                           n139);
   U2 : BUF_X2 port map( A => n139, Z => n140);
   U3 : BUF_X2 port map( A => n434, Z => n164);
   U4 : CLKBUF_X1 port map( A => n434, Z => n165);
   U5 : BUF_X2 port map( A => n432, Z => n152);
   U6 : CLKBUF_X1 port map( A => n432, Z => n153);
   U7 : BUF_X2 port map( A => n431, Z => n146);
   U8 : CLKBUF_X1 port map( A => n431, Z => n147);
   U9 : CLKBUF_X1 port map( A => n139, Z => n141);
   U10 : BUF_X2 port map( A => n433, Z => n158);
   U11 : CLKBUF_X1 port map( A => n433, Z => n159);
   U12 : CLKBUF_X1 port map( A => n434, Z => n166);
   U13 : CLKBUF_X1 port map( A => n432, Z => n154);
   U14 : CLKBUF_X1 port map( A => n431, Z => n148);
   U15 : CLKBUF_X1 port map( A => n139, Z => n142);
   U16 : CLKBUF_X1 port map( A => n433, Z => n160);
   U17 : CLKBUF_X1 port map( A => n434, Z => n167);
   U18 : CLKBUF_X1 port map( A => n432, Z => n155);
   U19 : CLKBUF_X1 port map( A => n431, Z => n149);
   U20 : CLKBUF_X1 port map( A => n139, Z => n143);
   U21 : CLKBUF_X1 port map( A => n433, Z => n161);
   U22 : CLKBUF_X1 port map( A => n434, Z => n168);
   U23 : CLKBUF_X1 port map( A => n432, Z => n156);
   U24 : CLKBUF_X1 port map( A => n431, Z => n150);
   U25 : CLKBUF_X1 port map( A => n139, Z => n144);
   U26 : CLKBUF_X1 port map( A => n433, Z => n162);
   U27 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U28 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U29 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN 
                           => Y(43));
   U30 : CLKBUF_X1 port map( A => n139, Z => n145);
   U31 : CLKBUF_X1 port map( A => n431, Z => n151);
   U32 : CLKBUF_X1 port map( A => n432, Z => n157);
   U33 : CLKBUF_X1 port map( A => n433, Z => n163);
   U34 : CLKBUF_X1 port map( A => n434, Z => n169);
   U35 : INV_X1 port map( A => SEL(1), ZN => n172);
   U36 : INV_X1 port map( A => SEL(2), ZN => n170);
   U37 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U38 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U39 : INV_X1 port map( A => SEL(0), ZN => n174);
   U40 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U41 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U42 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U43 : INV_X1 port map( A => n175, ZN => n431);
   U44 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U45 : INV_X1 port map( A => n176, ZN => n432);
   U46 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U47 : INV_X1 port map( A => n177, ZN => n434);
   U48 : INV_X1 port map( A => n178, ZN => n433);
   U49 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U50 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U51 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U52 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U53 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U54 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U55 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U56 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U57 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U58 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U59 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U60 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U61 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U62 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U63 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U64 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U65 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U66 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U67 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U68 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U69 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U70 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U71 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U72 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U73 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U74 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U75 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U76 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U77 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U78 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U79 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U80 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U81 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U82 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U83 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U84 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U85 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U86 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U87 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U88 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U89 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U90 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U91 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U92 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U93 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U94 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U95 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U96 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U97 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U98 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U99 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U100 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(10));
   U101 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U102 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U103 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U104 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U105 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN
                           => Y(11));
   U106 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U107 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U108 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U109 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U110 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U111 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U112 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U113 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U114 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U115 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U116 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U117 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U118 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U119 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U120 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U121 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U122 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U123 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U124 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U125 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U126 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U127 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U128 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U129 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U130 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U131 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U132 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U133 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U134 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U135 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U136 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U138 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U139 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U140 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U141 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U142 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U143 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U144 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U145 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U146 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U147 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U148 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U149 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U150 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U151 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U152 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U153 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U154 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U155 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U156 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U157 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U158 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U159 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U160 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U161 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U162 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U163 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U164 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U165 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U166 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U167 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U168 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U169 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U170 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U171 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U172 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U173 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U174 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U175 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U176 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U177 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U178 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U179 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U180 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U181 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U182 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U183 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U184 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U185 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U186 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U187 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U188 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U189 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U190 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U191 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U192 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U193 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U194 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U195 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U196 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U197 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U198 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U199 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U200 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U201 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U202 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U203 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U204 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U205 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U206 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U207 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U208 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U209 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U210 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U211 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U212 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U213 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U214 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U215 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U216 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U217 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U218 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U219 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U220 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U221 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U222 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U223 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U224 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U225 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U226 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U227 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U228 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U229 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U230 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U231 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U232 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U233 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U234 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U235 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U236 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U237 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U238 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U239 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U240 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U241 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U242 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U243 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U244 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U245 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U246 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U247 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U248 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U249 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U250 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U251 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U252 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U253 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U254 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U255 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U256 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U257 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U258 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U259 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U260 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U261 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U262 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U263 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U264 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U265 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U266 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U267 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U268 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U269 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U270 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U271 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U272 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U273 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U274 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U275 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U276 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U277 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U278 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U279 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U280 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U281 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U282 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U283 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U284 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U285 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U286 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U287 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U288 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U289 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U290 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U291 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U292 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U293 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U294 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U295 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U296 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U297 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U298 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U299 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U300 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U301 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U302 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U303 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U304 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U305 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U306 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U307 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U308 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U309 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U310 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U311 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U312 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U313 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U314 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U315 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U316 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U317 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U318 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U319 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U320 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U321 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U322 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U323 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U324 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U325 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U326 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U327 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U328 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U329 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U330 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U331 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U332 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U333 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U334 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U335 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U336 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U337 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U338 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U339 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U340 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U341 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U342 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U343 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U344 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U345 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U346 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U347 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U348 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U349 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U350 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U351 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U352 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U353 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U354 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => Y(61));
   U355 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U356 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U357 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U358 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U359 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => Y(62));
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_7 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_7;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_7 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X2 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U2 : NAND4_X2 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN 
                           => Y(62));
   U3 : BUF_X2 port map( A => n434, Z => n164);
   U4 : CLKBUF_X1 port map( A => n434, Z => n165);
   U5 : BUF_X2 port map( A => n432, Z => n152);
   U6 : BUF_X2 port map( A => n431, Z => n146);
   U7 : BUF_X2 port map( A => n139, Z => n140);
   U8 : CLKBUF_X1 port map( A => n139, Z => n141);
   U9 : BUF_X2 port map( A => n433, Z => n158);
   U10 : CLKBUF_X1 port map( A => n433, Z => n159);
   U11 : CLKBUF_X1 port map( A => n434, Z => n166);
   U12 : CLKBUF_X1 port map( A => n432, Z => n153);
   U13 : CLKBUF_X1 port map( A => n432, Z => n154);
   U14 : CLKBUF_X1 port map( A => n431, Z => n147);
   U15 : CLKBUF_X1 port map( A => n431, Z => n148);
   U16 : CLKBUF_X1 port map( A => n139, Z => n142);
   U17 : CLKBUF_X1 port map( A => n433, Z => n160);
   U18 : CLKBUF_X1 port map( A => n434, Z => n167);
   U19 : CLKBUF_X1 port map( A => n432, Z => n155);
   U20 : CLKBUF_X1 port map( A => n431, Z => n149);
   U21 : CLKBUF_X1 port map( A => n139, Z => n143);
   U22 : CLKBUF_X1 port map( A => n433, Z => n161);
   U23 : CLKBUF_X1 port map( A => n434, Z => n168);
   U24 : CLKBUF_X1 port map( A => n432, Z => n156);
   U25 : CLKBUF_X1 port map( A => n431, Z => n150);
   U26 : CLKBUF_X1 port map( A => n139, Z => n144);
   U27 : CLKBUF_X1 port map( A => n433, Z => n162);
   U28 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U29 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U30 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U31 : CLKBUF_X1 port map( A => n139, Z => n145);
   U32 : CLKBUF_X1 port map( A => n431, Z => n151);
   U33 : CLKBUF_X1 port map( A => n432, Z => n157);
   U34 : CLKBUF_X1 port map( A => n433, Z => n163);
   U35 : CLKBUF_X1 port map( A => n434, Z => n169);
   U36 : INV_X1 port map( A => SEL(1), ZN => n172);
   U37 : INV_X1 port map( A => SEL(2), ZN => n170);
   U38 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U39 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U40 : INV_X1 port map( A => SEL(0), ZN => n174);
   U41 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U42 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U43 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U44 : INV_X1 port map( A => n175, ZN => n431);
   U45 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U46 : INV_X1 port map( A => n176, ZN => n432);
   U47 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U48 : INV_X1 port map( A => n177, ZN => n434);
   U49 : INV_X1 port map( A => n178, ZN => n433);
   U50 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U51 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U52 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U53 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U54 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U55 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U56 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U57 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U58 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U59 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U60 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U61 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U62 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U63 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U64 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U65 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U66 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U67 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U68 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U69 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U70 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U71 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U72 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U73 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U74 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U75 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U76 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U77 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U78 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U79 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U80 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U81 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U82 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U83 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U84 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U85 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U86 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U87 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U88 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U89 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U90 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U91 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U92 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U93 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U94 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U95 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U96 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U97 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U98 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U99 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U100 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(10));
   U101 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U102 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U103 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U104 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U105 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN
                           => Y(11));
   U106 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U107 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U108 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U109 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U110 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U111 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U112 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U113 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U114 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U115 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U116 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U117 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U118 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U119 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U120 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U121 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U122 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U123 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U124 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U125 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U126 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U127 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U128 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U129 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U130 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U131 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U132 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U133 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U134 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U135 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U136 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U138 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U139 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U140 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U141 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U142 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U143 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U144 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U145 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U146 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U147 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U148 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U149 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U150 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U151 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U152 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U153 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U154 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U155 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U156 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U157 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U158 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U159 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U160 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U161 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U162 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U163 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U164 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U165 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U166 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U167 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U168 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U169 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U170 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U171 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U172 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U173 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U174 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U175 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U176 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U177 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U178 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U179 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U180 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U181 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U182 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U183 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U184 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U185 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U186 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U187 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U188 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U189 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U190 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U191 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U192 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U193 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U194 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U195 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U196 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U197 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U198 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U199 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U200 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U201 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U202 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U203 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U204 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U205 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U206 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U207 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U208 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U209 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U210 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U211 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U212 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U213 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U214 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U215 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U216 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U217 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U218 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U219 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U220 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U221 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U222 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U223 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U224 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U225 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U226 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U227 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U228 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U229 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U230 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U231 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U232 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U233 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U234 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U235 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U236 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U237 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U238 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U239 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U240 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U241 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U242 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U243 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U244 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U245 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U246 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U247 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U248 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U249 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U250 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U251 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U252 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U253 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U254 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U255 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U256 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U257 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U258 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U259 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U260 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U261 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U262 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U263 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U264 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U265 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U266 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U267 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U268 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U269 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U270 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U271 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U272 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U273 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U274 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U275 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U276 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U277 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U278 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U279 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U280 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U281 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U282 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U283 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U284 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U285 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U286 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U287 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U288 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U289 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U290 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U291 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U292 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U293 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U294 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U295 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U296 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U297 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U298 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U299 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U300 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U301 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U302 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U303 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U304 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U305 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U306 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U307 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U308 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U309 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U310 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U311 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U312 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U313 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U314 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U315 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U316 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U317 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U318 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U319 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U320 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U321 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U322 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U323 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U324 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U325 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U326 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U327 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U328 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U329 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U330 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U331 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U332 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U333 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U334 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U335 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U336 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U337 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U338 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U339 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U340 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U341 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U342 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U343 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U344 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U345 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U346 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U347 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U348 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U349 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U350 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U351 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U352 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U353 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U354 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U355 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => Y(61));
   U356 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U357 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U358 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U359 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_6 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_6;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_6 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X2 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN 
                           => Y(11));
   U2 : NAND4_X2 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN 
                           => Y(61));
   U3 : NAND4_X2 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN 
                           => Y(62));
   U4 : BUF_X2 port map( A => n434, Z => n164);
   U5 : BUF_X2 port map( A => n432, Z => n152);
   U6 : BUF_X2 port map( A => n431, Z => n146);
   U7 : BUF_X2 port map( A => n139, Z => n140);
   U8 : BUF_X2 port map( A => n433, Z => n158);
   U9 : CLKBUF_X1 port map( A => n434, Z => n165);
   U10 : CLKBUF_X1 port map( A => n434, Z => n166);
   U11 : CLKBUF_X1 port map( A => n432, Z => n153);
   U12 : CLKBUF_X1 port map( A => n432, Z => n154);
   U13 : CLKBUF_X1 port map( A => n431, Z => n147);
   U14 : CLKBUF_X1 port map( A => n431, Z => n148);
   U15 : CLKBUF_X1 port map( A => n139, Z => n141);
   U16 : CLKBUF_X1 port map( A => n139, Z => n142);
   U17 : CLKBUF_X1 port map( A => n433, Z => n159);
   U18 : CLKBUF_X1 port map( A => n433, Z => n160);
   U19 : CLKBUF_X1 port map( A => n434, Z => n167);
   U20 : CLKBUF_X1 port map( A => n432, Z => n155);
   U21 : CLKBUF_X1 port map( A => n431, Z => n149);
   U22 : CLKBUF_X1 port map( A => n139, Z => n143);
   U23 : CLKBUF_X1 port map( A => n433, Z => n161);
   U24 : CLKBUF_X1 port map( A => n434, Z => n168);
   U25 : CLKBUF_X1 port map( A => n432, Z => n156);
   U26 : CLKBUF_X1 port map( A => n431, Z => n150);
   U27 : CLKBUF_X1 port map( A => n139, Z => n144);
   U28 : CLKBUF_X1 port map( A => n433, Z => n162);
   U29 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U30 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U31 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U32 : CLKBUF_X1 port map( A => n139, Z => n145);
   U33 : CLKBUF_X1 port map( A => n431, Z => n151);
   U34 : CLKBUF_X1 port map( A => n432, Z => n157);
   U35 : CLKBUF_X1 port map( A => n433, Z => n163);
   U36 : CLKBUF_X1 port map( A => n434, Z => n169);
   U37 : INV_X1 port map( A => SEL(1), ZN => n172);
   U38 : INV_X1 port map( A => SEL(2), ZN => n170);
   U39 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U40 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U41 : INV_X1 port map( A => SEL(0), ZN => n174);
   U42 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U43 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U44 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U45 : INV_X1 port map( A => n175, ZN => n431);
   U46 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U47 : INV_X1 port map( A => n176, ZN => n432);
   U48 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U49 : INV_X1 port map( A => n177, ZN => n434);
   U50 : INV_X1 port map( A => n178, ZN => n433);
   U51 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U52 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U53 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U54 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U55 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U56 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U57 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U58 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U59 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U60 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U61 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U62 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U63 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U64 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U65 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U66 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U67 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U68 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U69 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U70 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U71 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U72 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U73 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U74 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U75 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U76 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U77 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U78 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U79 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U80 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U81 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U82 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U83 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U84 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U85 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U86 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U87 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U88 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U89 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U90 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U91 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U92 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U93 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U94 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U95 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U96 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U97 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U98 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U99 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U100 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U101 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U102 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(10));
   U103 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U104 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U105 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U106 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U107 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U108 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U109 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U110 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U111 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U112 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U113 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U114 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U115 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U116 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U117 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U118 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U119 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U120 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U121 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U122 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U123 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U124 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U125 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U126 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U127 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U128 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U129 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U130 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U131 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U132 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U133 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U134 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U135 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U136 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U137 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U138 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U139 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U140 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U141 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U142 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U143 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U144 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U145 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U146 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U147 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U148 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U149 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U150 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U151 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U152 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U153 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U154 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U155 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U156 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U157 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U158 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U159 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U160 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U161 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U162 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U163 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U164 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U165 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U166 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U167 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U168 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U169 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U170 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U171 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U172 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U173 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U174 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U175 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U176 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U177 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U178 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U179 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U180 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U181 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U182 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U183 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U184 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U185 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U186 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U187 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U188 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U189 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U190 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U191 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U192 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U193 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U194 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U195 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U196 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U197 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U198 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U199 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U200 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U201 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U202 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U203 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U204 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U205 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U206 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U207 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U208 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U209 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U210 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U211 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U212 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U213 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U214 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U215 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U216 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U217 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U218 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U219 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U220 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U221 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U222 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U223 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U224 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U225 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U226 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U227 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U228 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U229 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U230 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U231 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U232 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U233 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U234 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U235 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U236 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U237 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U238 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U239 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U240 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U241 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U242 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U243 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U244 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U245 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U246 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U247 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U248 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U249 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U250 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U251 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U252 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U253 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U254 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U255 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U256 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U257 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U258 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U259 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U260 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U261 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U262 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U263 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U264 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U265 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U266 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U267 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U268 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U269 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U270 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U271 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U272 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U273 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U274 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U275 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U276 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U277 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U278 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U279 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U280 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U281 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U282 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U283 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U284 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U285 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U286 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U287 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U288 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U289 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U290 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U291 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U292 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U293 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U294 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U295 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U296 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U297 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U298 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U299 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U300 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U301 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U302 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U303 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U304 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U305 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U306 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U307 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U308 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U309 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U310 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U311 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U312 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U313 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U314 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U315 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U316 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U317 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U318 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U319 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U320 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U321 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U322 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U323 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U324 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U325 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U326 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U327 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U328 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U329 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U330 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U331 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U332 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U333 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U334 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U335 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U336 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U337 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U338 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U339 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U340 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U341 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U342 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U343 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U344 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U345 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U346 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U347 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U348 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U349 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U350 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U351 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U352 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U353 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U354 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U355 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U356 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U357 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U358 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U359 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_5 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_5;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_5 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X2 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN 
                           => Y(10));
   U2 : NAND4_X2 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U3 : BUF_X2 port map( A => n434, Z => n164);
   U4 : BUF_X2 port map( A => n432, Z => n152);
   U5 : BUF_X2 port map( A => n431, Z => n146);
   U6 : BUF_X2 port map( A => n139, Z => n140);
   U7 : BUF_X2 port map( A => n433, Z => n158);
   U8 : CLKBUF_X1 port map( A => n434, Z => n165);
   U9 : CLKBUF_X1 port map( A => n432, Z => n153);
   U10 : CLKBUF_X1 port map( A => n431, Z => n147);
   U11 : CLKBUF_X1 port map( A => n139, Z => n141);
   U12 : CLKBUF_X1 port map( A => n433, Z => n159);
   U13 : CLKBUF_X1 port map( A => n434, Z => n167);
   U14 : CLKBUF_X1 port map( A => n434, Z => n166);
   U15 : CLKBUF_X1 port map( A => n432, Z => n155);
   U16 : CLKBUF_X1 port map( A => n432, Z => n154);
   U17 : CLKBUF_X1 port map( A => n431, Z => n149);
   U18 : CLKBUF_X1 port map( A => n431, Z => n148);
   U19 : CLKBUF_X1 port map( A => n139, Z => n142);
   U20 : CLKBUF_X1 port map( A => n139, Z => n143);
   U21 : CLKBUF_X1 port map( A => n433, Z => n161);
   U22 : CLKBUF_X1 port map( A => n433, Z => n160);
   U23 : CLKBUF_X1 port map( A => n434, Z => n168);
   U24 : CLKBUF_X1 port map( A => n432, Z => n156);
   U25 : CLKBUF_X1 port map( A => n431, Z => n150);
   U26 : CLKBUF_X1 port map( A => n139, Z => n144);
   U27 : CLKBUF_X1 port map( A => n433, Z => n162);
   U28 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U29 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U30 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U31 : CLKBUF_X1 port map( A => n139, Z => n145);
   U32 : CLKBUF_X1 port map( A => n431, Z => n151);
   U33 : CLKBUF_X1 port map( A => n432, Z => n157);
   U34 : CLKBUF_X1 port map( A => n433, Z => n163);
   U35 : CLKBUF_X1 port map( A => n434, Z => n169);
   U36 : INV_X1 port map( A => SEL(1), ZN => n172);
   U37 : INV_X1 port map( A => SEL(2), ZN => n170);
   U38 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U39 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U40 : INV_X1 port map( A => SEL(0), ZN => n174);
   U41 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U42 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U43 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U44 : INV_X1 port map( A => n175, ZN => n431);
   U45 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U46 : INV_X1 port map( A => n176, ZN => n432);
   U47 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U48 : INV_X1 port map( A => n177, ZN => n434);
   U49 : INV_X1 port map( A => n178, ZN => n433);
   U50 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U51 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U52 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U53 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U54 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U55 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U56 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U57 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U58 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U59 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U60 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U61 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U62 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U63 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U64 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U65 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U66 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U67 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U68 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U69 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U70 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U71 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U72 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U73 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U74 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U75 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U76 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U77 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U78 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U79 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U80 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U81 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U82 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U83 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U84 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U85 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U86 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U87 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U88 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U89 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U90 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U91 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U92 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U93 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U94 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U95 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U96 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U97 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U98 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U99 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U100 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U101 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U102 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U103 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U104 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN
                           => Y(11));
   U105 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U106 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U107 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U108 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U109 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U110 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U111 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U112 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U113 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U114 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U115 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U116 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U117 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U118 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U119 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U120 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U121 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U122 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U123 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U124 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U125 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U126 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U127 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U128 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U129 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U130 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U131 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U132 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U133 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U134 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U135 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U136 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U137 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U138 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U139 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U140 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U141 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U142 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U143 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U144 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U145 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U146 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U147 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U148 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U149 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U150 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U151 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U152 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U153 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U154 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U155 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U156 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U157 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U158 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U159 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U160 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U161 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U162 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U163 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U164 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U165 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U166 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U167 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U168 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U169 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U170 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U171 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U172 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U173 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U174 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U175 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U176 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U177 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U178 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U179 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U180 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U181 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U182 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U183 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U184 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U185 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U186 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U187 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U188 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U189 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U190 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U191 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U192 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U193 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U194 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U195 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U196 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U197 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U198 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U199 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U200 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U201 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U202 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U203 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U204 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U205 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U206 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U207 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U208 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U209 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U210 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U211 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U212 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U213 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U214 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U215 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U216 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U217 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U218 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U219 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U220 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U221 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U222 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U223 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U224 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U225 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U226 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U227 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U228 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U229 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U230 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U231 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U232 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U233 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U234 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U235 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U236 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U237 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U238 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U239 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U240 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U241 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U242 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U243 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U244 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U245 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U246 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U247 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U248 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U249 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U250 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U251 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U252 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U253 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U254 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U255 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U256 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U257 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U258 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U259 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U260 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U261 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U262 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U263 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U264 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U265 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U266 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U267 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U268 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U269 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U270 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U271 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U272 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U273 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U274 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U275 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U276 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U277 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U278 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U279 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U280 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U281 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U282 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U283 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U284 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U285 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U286 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U287 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U288 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U289 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U290 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U291 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U292 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U293 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U294 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U295 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U296 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U297 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U298 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U299 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U300 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U301 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U302 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U303 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U304 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U305 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U306 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U307 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U308 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U309 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U310 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U311 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U312 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U313 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U314 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U315 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U316 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U317 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U318 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U319 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U320 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U321 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U322 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U323 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U324 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U325 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U326 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U327 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U328 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U329 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U330 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U331 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U332 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U333 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U334 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U335 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U336 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U337 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U338 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U339 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U340 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U341 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U342 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U343 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U344 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U345 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U346 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U347 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U348 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U349 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U350 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U351 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U352 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U353 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U354 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => Y(61));
   U355 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U356 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U357 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U358 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U359 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => Y(62));
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_4 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_4;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_4 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN 
                           => Y(61));
   U2 : NAND4_X2 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U3 : NAND4_X2 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN 
                           => Y(11));
   U4 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN =>
                           n139);
   U5 : BUF_X2 port map( A => n434, Z => n164);
   U6 : BUF_X2 port map( A => n432, Z => n152);
   U7 : BUF_X2 port map( A => n431, Z => n146);
   U8 : BUF_X2 port map( A => n139, Z => n140);
   U9 : BUF_X2 port map( A => n433, Z => n158);
   U10 : CLKBUF_X1 port map( A => n434, Z => n165);
   U11 : CLKBUF_X1 port map( A => n432, Z => n153);
   U12 : CLKBUF_X1 port map( A => n431, Z => n147);
   U13 : CLKBUF_X1 port map( A => n139, Z => n141);
   U14 : CLKBUF_X1 port map( A => n433, Z => n159);
   U15 : CLKBUF_X1 port map( A => n434, Z => n166);
   U16 : CLKBUF_X1 port map( A => n432, Z => n154);
   U17 : CLKBUF_X1 port map( A => n431, Z => n148);
   U18 : CLKBUF_X1 port map( A => n139, Z => n142);
   U19 : CLKBUF_X1 port map( A => n139, Z => n143);
   U20 : CLKBUF_X1 port map( A => n433, Z => n160);
   U21 : CLKBUF_X1 port map( A => n434, Z => n168);
   U22 : CLKBUF_X1 port map( A => n434, Z => n167);
   U23 : CLKBUF_X1 port map( A => n432, Z => n156);
   U24 : CLKBUF_X1 port map( A => n432, Z => n155);
   U25 : CLKBUF_X1 port map( A => n431, Z => n150);
   U26 : CLKBUF_X1 port map( A => n431, Z => n149);
   U27 : CLKBUF_X1 port map( A => n139, Z => n144);
   U28 : CLKBUF_X1 port map( A => n433, Z => n162);
   U29 : CLKBUF_X1 port map( A => n433, Z => n161);
   U30 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U31 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U32 : CLKBUF_X1 port map( A => n139, Z => n145);
   U33 : CLKBUF_X1 port map( A => n431, Z => n151);
   U34 : CLKBUF_X1 port map( A => n432, Z => n157);
   U35 : CLKBUF_X1 port map( A => n433, Z => n163);
   U36 : CLKBUF_X1 port map( A => n434, Z => n169);
   U37 : INV_X1 port map( A => SEL(1), ZN => n172);
   U38 : INV_X1 port map( A => SEL(2), ZN => n170);
   U39 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U40 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U41 : INV_X1 port map( A => SEL(0), ZN => n174);
   U42 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U43 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U44 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U45 : INV_X1 port map( A => n175, ZN => n431);
   U46 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U47 : INV_X1 port map( A => n176, ZN => n432);
   U48 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U49 : INV_X1 port map( A => n177, ZN => n434);
   U50 : INV_X1 port map( A => n178, ZN => n433);
   U51 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U52 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U53 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U54 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U55 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U56 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U57 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U58 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U59 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U60 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U61 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U62 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U63 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U64 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U65 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U66 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U67 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U68 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U69 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U70 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U71 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U72 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U73 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U74 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U75 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U76 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U77 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U78 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U79 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U80 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U81 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U82 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U83 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U84 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U85 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U86 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U87 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U88 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U89 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U90 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U91 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U92 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U93 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U94 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U95 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U96 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U97 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U98 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U99 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U100 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U101 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(10));
   U102 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U103 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U104 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U105 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U106 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U107 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U108 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U109 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U110 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U111 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U112 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U113 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U114 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U115 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U116 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U117 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U118 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U119 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U120 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U121 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U122 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U123 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U124 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U125 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U126 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U127 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U128 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U129 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U130 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U131 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U132 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U133 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U134 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U135 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U136 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U138 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U139 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U140 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U141 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U142 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U143 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U144 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U145 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U146 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U147 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U148 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U149 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U150 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U151 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U152 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U153 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U154 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U155 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U156 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U157 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U158 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U159 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U160 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U161 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U162 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U163 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U164 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U165 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U166 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U167 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U168 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U169 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U170 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U171 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U172 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U173 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U174 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U175 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U176 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U177 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U178 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U179 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U180 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U181 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U182 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U183 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U184 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U185 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U186 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U187 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U188 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U189 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U190 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U191 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U192 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U193 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U194 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U195 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U196 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U197 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U198 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U199 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U200 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U201 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U202 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U203 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U204 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U205 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U206 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U207 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U208 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U209 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U210 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U211 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U212 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U213 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U214 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U215 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U216 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U217 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U218 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U219 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U220 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U221 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U222 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U223 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U224 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U225 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U226 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U227 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U228 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U229 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U230 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U231 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U232 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U233 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U234 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U235 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U236 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U237 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U238 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U239 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U240 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U241 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U242 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U243 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U244 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U245 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U246 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U247 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U248 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U249 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U250 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U251 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U252 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U253 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U254 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U255 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U256 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U257 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U258 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U259 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U260 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U261 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U262 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U263 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U264 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U265 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U266 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U267 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U268 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U269 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U270 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U271 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U272 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U273 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U274 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U275 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U276 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U277 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U278 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U279 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U280 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U281 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U282 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U283 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U284 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U285 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U286 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U287 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U288 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U289 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U290 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U291 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U292 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U293 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U294 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U295 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U296 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U297 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U298 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U299 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U300 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U301 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U302 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U303 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U304 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U305 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U306 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U307 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U308 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U309 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U310 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U311 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U312 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U313 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U314 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U315 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U316 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U317 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U318 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U319 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U320 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U321 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U322 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U323 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U324 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U325 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U326 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U327 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U328 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U329 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U330 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U331 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U332 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U333 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U334 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U335 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U336 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U337 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U338 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U339 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U340 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U341 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U342 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U343 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U344 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U345 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U346 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U347 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U348 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U349 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U350 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U351 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U352 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U353 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U354 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U355 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U356 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U357 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U358 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U359 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => Y(62));
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_3 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_3;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_3 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN 
                           => Y(61));
   U2 : NAND4_X2 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN 
                           => Y(60));
   U3 : BUF_X1 port map( A => n434, Z => n164);
   U4 : BUF_X1 port map( A => n432, Z => n152);
   U5 : BUF_X1 port map( A => n431, Z => n146);
   U6 : BUF_X1 port map( A => n139, Z => n140);
   U7 : BUF_X1 port map( A => n433, Z => n158);
   U8 : CLKBUF_X1 port map( A => n434, Z => n165);
   U9 : CLKBUF_X1 port map( A => n432, Z => n153);
   U10 : CLKBUF_X1 port map( A => n431, Z => n147);
   U11 : CLKBUF_X1 port map( A => n139, Z => n141);
   U12 : CLKBUF_X1 port map( A => n433, Z => n159);
   U13 : CLKBUF_X1 port map( A => n434, Z => n166);
   U14 : CLKBUF_X1 port map( A => n432, Z => n154);
   U15 : CLKBUF_X1 port map( A => n431, Z => n148);
   U16 : CLKBUF_X1 port map( A => n139, Z => n142);
   U17 : CLKBUF_X1 port map( A => n433, Z => n160);
   U18 : CLKBUF_X1 port map( A => n434, Z => n168);
   U19 : CLKBUF_X1 port map( A => n434, Z => n167);
   U20 : CLKBUF_X1 port map( A => n432, Z => n156);
   U21 : CLKBUF_X1 port map( A => n432, Z => n155);
   U22 : CLKBUF_X1 port map( A => n431, Z => n150);
   U23 : CLKBUF_X1 port map( A => n431, Z => n149);
   U24 : CLKBUF_X1 port map( A => n139, Z => n144);
   U25 : CLKBUF_X1 port map( A => n139, Z => n143);
   U26 : CLKBUF_X1 port map( A => n433, Z => n162);
   U27 : CLKBUF_X1 port map( A => n433, Z => n161);
   U28 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U29 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U30 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U31 : CLKBUF_X1 port map( A => n139, Z => n145);
   U32 : CLKBUF_X1 port map( A => n431, Z => n151);
   U33 : CLKBUF_X1 port map( A => n432, Z => n157);
   U34 : CLKBUF_X1 port map( A => n433, Z => n163);
   U35 : CLKBUF_X1 port map( A => n434, Z => n169);
   U36 : INV_X1 port map( A => SEL(1), ZN => n172);
   U37 : INV_X1 port map( A => SEL(2), ZN => n170);
   U38 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U39 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U40 : INV_X1 port map( A => SEL(0), ZN => n174);
   U41 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U42 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U43 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U44 : INV_X1 port map( A => n175, ZN => n431);
   U45 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U46 : INV_X1 port map( A => n176, ZN => n432);
   U47 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U48 : INV_X1 port map( A => n177, ZN => n434);
   U49 : INV_X1 port map( A => n178, ZN => n433);
   U50 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U51 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U52 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U53 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U54 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U55 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U56 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U57 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U58 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U59 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U60 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U61 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U62 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U63 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U64 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U65 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U66 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U67 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U68 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U69 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U70 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U71 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U72 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U73 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U74 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U75 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U76 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U77 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U78 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U79 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U80 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U81 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U82 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U83 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U84 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U85 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U86 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U87 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U88 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U89 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U90 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U91 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U92 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U93 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U94 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U95 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U96 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U97 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U98 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U99 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U100 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U101 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(10));
   U102 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U103 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U104 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U105 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U106 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN
                           => Y(11));
   U107 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U108 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U109 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U110 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U111 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U112 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U113 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U114 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U115 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U116 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U117 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U118 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U119 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U120 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U121 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U122 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U123 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U124 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U125 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U126 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U127 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U128 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U129 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U130 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U131 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U132 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U133 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U134 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U135 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U136 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U137 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U138 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U139 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U140 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U141 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U142 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U143 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U144 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U145 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U146 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U147 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U148 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U149 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U150 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U151 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U152 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U153 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U154 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U155 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U156 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U157 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U158 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U159 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U160 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U161 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U162 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U163 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U164 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U165 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U166 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U167 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U168 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U169 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U170 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U171 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U172 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U173 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U174 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U175 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U176 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U177 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U178 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U179 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U180 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U181 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U182 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U183 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U184 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U185 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U186 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U187 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U188 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U189 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U190 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U191 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U192 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U193 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U194 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U195 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U196 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U197 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U198 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U199 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U200 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U201 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U202 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U203 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U204 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U205 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U206 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U207 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U208 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U209 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U210 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U211 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U212 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U213 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U214 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U215 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U216 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U217 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U218 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U219 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U220 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U221 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U222 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U223 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U224 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U225 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U226 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U227 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U228 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U229 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U230 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U231 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U232 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U233 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U234 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U235 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U236 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U237 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U238 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U239 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U240 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U241 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U242 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U243 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U244 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U245 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U246 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U247 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U248 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U249 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U250 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U251 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U252 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U253 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U254 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U255 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U256 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U257 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U258 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U259 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U260 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U261 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U262 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U263 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U264 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U265 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U266 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U267 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U268 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U269 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U270 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U271 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U272 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U273 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U274 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U275 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U276 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U277 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U278 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U279 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U280 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U281 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U282 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U283 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U284 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U285 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U286 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U287 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U288 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U289 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U290 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U291 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U292 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U293 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U294 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U295 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U296 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U297 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U298 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U299 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U300 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U301 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U302 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U303 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U304 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U305 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U306 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U307 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U308 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U309 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U310 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U311 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U312 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U313 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U314 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U315 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U316 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U317 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U318 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U319 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U320 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U321 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U322 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U323 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U324 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U325 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U326 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U327 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U328 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U329 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U330 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U331 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U332 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U333 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U334 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U335 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U336 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U337 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U338 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U339 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U340 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U341 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U342 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U343 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U344 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U345 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U346 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U347 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U348 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U349 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U350 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U351 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U352 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U353 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U354 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U355 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U356 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U357 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U358 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U359 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => Y(62));
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_2 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_2;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_2 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : NAND4_X2 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN 
                           => Y(61));
   U2 : CLKBUF_X1 port map( A => n434, Z => n165);
   U3 : CLKBUF_X1 port map( A => n431, Z => n147);
   U4 : CLKBUF_X1 port map( A => n432, Z => n153);
   U5 : CLKBUF_X1 port map( A => n433, Z => n159);
   U6 : BUF_X1 port map( A => n139, Z => n140);
   U7 : BUF_X1 port map( A => n434, Z => n164);
   U8 : BUF_X1 port map( A => n432, Z => n152);
   U9 : BUF_X1 port map( A => n431, Z => n146);
   U10 : CLKBUF_X1 port map( A => n139, Z => n141);
   U11 : BUF_X1 port map( A => n433, Z => n158);
   U12 : CLKBUF_X1 port map( A => n434, Z => n166);
   U13 : CLKBUF_X1 port map( A => n432, Z => n154);
   U14 : CLKBUF_X1 port map( A => n431, Z => n148);
   U15 : CLKBUF_X1 port map( A => n139, Z => n142);
   U16 : CLKBUF_X1 port map( A => n433, Z => n160);
   U17 : CLKBUF_X1 port map( A => n434, Z => n167);
   U18 : CLKBUF_X1 port map( A => n432, Z => n155);
   U19 : CLKBUF_X1 port map( A => n431, Z => n149);
   U20 : CLKBUF_X1 port map( A => n139, Z => n143);
   U21 : CLKBUF_X1 port map( A => n433, Z => n161);
   U22 : CLKBUF_X1 port map( A => n434, Z => n168);
   U23 : CLKBUF_X1 port map( A => n432, Z => n156);
   U24 : CLKBUF_X1 port map( A => n431, Z => n150);
   U25 : CLKBUF_X1 port map( A => n139, Z => n144);
   U26 : CLKBUF_X1 port map( A => n433, Z => n162);
   U27 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U28 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U29 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U30 : CLKBUF_X1 port map( A => n139, Z => n145);
   U31 : CLKBUF_X1 port map( A => n431, Z => n151);
   U32 : CLKBUF_X1 port map( A => n432, Z => n157);
   U33 : CLKBUF_X1 port map( A => n433, Z => n163);
   U34 : CLKBUF_X1 port map( A => n434, Z => n169);
   U35 : INV_X1 port map( A => SEL(1), ZN => n172);
   U36 : INV_X1 port map( A => SEL(2), ZN => n170);
   U37 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U38 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U39 : INV_X1 port map( A => SEL(0), ZN => n174);
   U40 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U41 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U42 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U43 : INV_X1 port map( A => n175, ZN => n431);
   U44 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U45 : INV_X1 port map( A => n176, ZN => n432);
   U46 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U47 : INV_X1 port map( A => n177, ZN => n434);
   U48 : INV_X1 port map( A => n178, ZN => n433);
   U49 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U50 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U51 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U52 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U53 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U54 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U55 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U56 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U57 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U58 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U59 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U60 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U61 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U62 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U63 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U64 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U65 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U66 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U67 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U68 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U69 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U70 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U71 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U72 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U73 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U74 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U75 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U76 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U77 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U78 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U79 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U80 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U81 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U82 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U83 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U84 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U85 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U86 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U87 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U88 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U89 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U90 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U91 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U92 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U93 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U94 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U95 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U96 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U97 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U98 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U99 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U100 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN
                           => Y(10));
   U101 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U102 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U103 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U104 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U105 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN
                           => Y(11));
   U106 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U107 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U108 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U109 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U110 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U111 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U112 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U113 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U114 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U115 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U116 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U117 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U118 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U119 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U120 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U121 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U122 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U123 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U124 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U125 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U126 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U127 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U128 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U129 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U130 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U131 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U132 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U133 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U134 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U135 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U136 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U137 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U138 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U139 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U140 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U141 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U142 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U143 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U144 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U145 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U146 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U147 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U148 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U149 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U150 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U151 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U152 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U153 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U154 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U155 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U156 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U157 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U158 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U159 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U160 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U161 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U162 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U163 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U164 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U165 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U166 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U167 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U168 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U169 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U170 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U171 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U172 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U173 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U174 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U175 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U176 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U177 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U178 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U179 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U180 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U181 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U182 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U183 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U184 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U185 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U186 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U187 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U188 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U189 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U190 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U191 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U192 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U193 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U194 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U195 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U196 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U197 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U198 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U199 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U200 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U201 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U202 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U203 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U204 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U205 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U206 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U207 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U208 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U209 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U210 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U211 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U212 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U213 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U214 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U215 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U216 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U217 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U218 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U219 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U220 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U221 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U222 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U223 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U224 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U225 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U226 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U227 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U228 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U229 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U230 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U231 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U232 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U233 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U234 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U235 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U236 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U237 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U238 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U239 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U240 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U241 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U242 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U243 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U244 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U245 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U246 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U247 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U248 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U249 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U250 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U251 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U252 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U253 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U254 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U255 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U256 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U257 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U258 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U259 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U260 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U261 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U262 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U263 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U264 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U265 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U266 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U267 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U268 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U269 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U270 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U271 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U272 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U273 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U274 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U275 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U276 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U277 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U278 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U279 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U280 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U281 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U282 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U283 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U284 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U285 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U286 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U287 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U288 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U289 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U290 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U291 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U292 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U293 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U294 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U295 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U296 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U297 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U298 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U299 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U300 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U301 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U302 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U303 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U304 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U305 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U306 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U307 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U308 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U309 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U310 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U311 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U312 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U313 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U314 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U315 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U316 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U317 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U318 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U319 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U320 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U321 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U322 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U323 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U324 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U325 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U326 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U327 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U328 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U329 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U330 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U331 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U332 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U333 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U334 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U335 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U336 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U337 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U338 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U339 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U340 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U341 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U342 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U343 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U344 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U345 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U346 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U347 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U348 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U349 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U350 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U351 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U352 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U353 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U354 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U355 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U356 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U357 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U358 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U359 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => Y(62));
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_1 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_1;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_1 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, 
      n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, 
      n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, 
      n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, 
      n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, 
      n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, 
      n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, 
      n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, 
      n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, 
      n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, 
      n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, 
      n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, 
      n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, 
      n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, 
      n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, 
      n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, 
      n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, 
      n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, 
      n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365, 
      n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, 
      n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389, 
      n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, 
      n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, 
      n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, 
      n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, 
      n438 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n434, Z => n164);
   U2 : BUF_X1 port map( A => n432, Z => n152);
   U3 : BUF_X1 port map( A => n431, Z => n146);
   U4 : BUF_X1 port map( A => n139, Z => n140);
   U5 : CLKBUF_X1 port map( A => n139, Z => n141);
   U6 : BUF_X1 port map( A => n433, Z => n158);
   U7 : CLKBUF_X1 port map( A => n434, Z => n165);
   U8 : CLKBUF_X1 port map( A => n434, Z => n166);
   U9 : CLKBUF_X1 port map( A => n432, Z => n153);
   U10 : CLKBUF_X1 port map( A => n432, Z => n154);
   U11 : CLKBUF_X1 port map( A => n431, Z => n147);
   U12 : CLKBUF_X1 port map( A => n431, Z => n148);
   U13 : CLKBUF_X1 port map( A => n139, Z => n142);
   U14 : CLKBUF_X1 port map( A => n433, Z => n159);
   U15 : CLKBUF_X1 port map( A => n433, Z => n160);
   U16 : CLKBUF_X1 port map( A => n434, Z => n167);
   U17 : CLKBUF_X1 port map( A => n432, Z => n155);
   U18 : CLKBUF_X1 port map( A => n431, Z => n149);
   U19 : CLKBUF_X1 port map( A => n139, Z => n143);
   U20 : CLKBUF_X1 port map( A => n433, Z => n161);
   U21 : CLKBUF_X1 port map( A => n434, Z => n168);
   U22 : CLKBUF_X1 port map( A => n432, Z => n156);
   U23 : CLKBUF_X1 port map( A => n431, Z => n150);
   U24 : CLKBUF_X1 port map( A => n139, Z => n144);
   U25 : CLKBUF_X1 port map( A => n433, Z => n162);
   U26 : AND4_X1 port map( A1 => n175, A2 => n176, A3 => n178, A4 => n177, ZN 
                           => n139);
   U27 : NAND2_X1 port map( A1 => n174, A2 => n173, ZN => n177);
   U28 : NAND2_X1 port map( A1 => n174, A2 => n171, ZN => n178);
   U29 : CLKBUF_X1 port map( A => n139, Z => n145);
   U30 : CLKBUF_X1 port map( A => n431, Z => n151);
   U31 : CLKBUF_X1 port map( A => n432, Z => n157);
   U32 : CLKBUF_X1 port map( A => n433, Z => n163);
   U33 : CLKBUF_X1 port map( A => n434, Z => n169);
   U34 : INV_X1 port map( A => SEL(1), ZN => n172);
   U35 : INV_X1 port map( A => SEL(2), ZN => n170);
   U36 : NAND3_X1 port map( A1 => SEL(0), A2 => n172, A3 => n170, ZN => n175);
   U37 : NAND3_X1 port map( A1 => SEL(0), A2 => SEL(1), A3 => n170, ZN => n176)
                           ;
   U38 : INV_X1 port map( A => SEL(0), ZN => n174);
   U39 : NOR2_X1 port map( A1 => SEL(1), A2 => SEL(2), ZN => n171);
   U40 : NOR2_X1 port map( A1 => n172, A2 => SEL(2), ZN => n173);
   U41 : NAND2_X1 port map( A1 => E(0), A2 => n140, ZN => n182);
   U42 : INV_X1 port map( A => n175, ZN => n431);
   U43 : NAND2_X1 port map( A1 => B(0), A2 => n146, ZN => n181);
   U44 : INV_X1 port map( A => n176, ZN => n432);
   U45 : NAND2_X1 port map( A1 => D(0), A2 => n152, ZN => n180);
   U46 : INV_X1 port map( A => n177, ZN => n434);
   U47 : INV_X1 port map( A => n178, ZN => n433);
   U48 : AOI22_X1 port map( A1 => C(0), A2 => n164, B1 => A(0), B2 => n158, ZN 
                           => n179);
   U49 : NAND4_X1 port map( A1 => n182, A2 => n181, A3 => n180, A4 => n179, ZN 
                           => Y(0));
   U50 : NAND2_X1 port map( A1 => E(1), A2 => n140, ZN => n186);
   U51 : NAND2_X1 port map( A1 => B(1), A2 => n146, ZN => n185);
   U52 : NAND2_X1 port map( A1 => D(1), A2 => n152, ZN => n184);
   U53 : AOI22_X1 port map( A1 => C(1), A2 => n164, B1 => A(1), B2 => n158, ZN 
                           => n183);
   U54 : NAND4_X1 port map( A1 => n186, A2 => n185, A3 => n184, A4 => n183, ZN 
                           => Y(1));
   U55 : NAND2_X1 port map( A1 => E(2), A2 => n140, ZN => n190);
   U56 : NAND2_X1 port map( A1 => B(2), A2 => n146, ZN => n189);
   U57 : NAND2_X1 port map( A1 => D(2), A2 => n152, ZN => n188);
   U58 : AOI22_X1 port map( A1 => C(2), A2 => n164, B1 => A(2), B2 => n158, ZN 
                           => n187);
   U59 : NAND4_X1 port map( A1 => n190, A2 => n189, A3 => n188, A4 => n187, ZN 
                           => Y(2));
   U60 : NAND2_X1 port map( A1 => E(3), A2 => n140, ZN => n194);
   U61 : NAND2_X1 port map( A1 => B(3), A2 => n146, ZN => n193);
   U62 : NAND2_X1 port map( A1 => D(3), A2 => n152, ZN => n192);
   U63 : AOI22_X1 port map( A1 => C(3), A2 => n164, B1 => A(3), B2 => n158, ZN 
                           => n191);
   U64 : NAND4_X1 port map( A1 => n194, A2 => n193, A3 => n192, A4 => n191, ZN 
                           => Y(3));
   U65 : NAND2_X1 port map( A1 => E(4), A2 => n140, ZN => n198);
   U66 : NAND2_X1 port map( A1 => B(4), A2 => n146, ZN => n197);
   U67 : NAND2_X1 port map( A1 => D(4), A2 => n152, ZN => n196);
   U68 : AOI22_X1 port map( A1 => C(4), A2 => n164, B1 => A(4), B2 => n158, ZN 
                           => n195);
   U69 : NAND4_X1 port map( A1 => n198, A2 => n197, A3 => n196, A4 => n195, ZN 
                           => Y(4));
   U70 : NAND2_X1 port map( A1 => E(5), A2 => n140, ZN => n202);
   U71 : NAND2_X1 port map( A1 => B(5), A2 => n146, ZN => n201);
   U72 : NAND2_X1 port map( A1 => D(5), A2 => n152, ZN => n200);
   U73 : AOI22_X1 port map( A1 => C(5), A2 => n164, B1 => A(5), B2 => n158, ZN 
                           => n199);
   U74 : NAND4_X1 port map( A1 => n202, A2 => n201, A3 => n200, A4 => n199, ZN 
                           => Y(5));
   U75 : NAND2_X1 port map( A1 => E(6), A2 => n140, ZN => n206);
   U76 : NAND2_X1 port map( A1 => B(6), A2 => n146, ZN => n205);
   U77 : NAND2_X1 port map( A1 => D(6), A2 => n152, ZN => n204);
   U78 : AOI22_X1 port map( A1 => C(6), A2 => n164, B1 => A(6), B2 => n158, ZN 
                           => n203);
   U79 : NAND4_X1 port map( A1 => n206, A2 => n205, A3 => n204, A4 => n203, ZN 
                           => Y(6));
   U80 : NAND2_X1 port map( A1 => E(7), A2 => n140, ZN => n210);
   U81 : NAND2_X1 port map( A1 => B(7), A2 => n146, ZN => n209);
   U82 : NAND2_X1 port map( A1 => D(7), A2 => n152, ZN => n208);
   U83 : AOI22_X1 port map( A1 => C(7), A2 => n164, B1 => A(7), B2 => n158, ZN 
                           => n207);
   U84 : NAND4_X1 port map( A1 => n210, A2 => n209, A3 => n208, A4 => n207, ZN 
                           => Y(7));
   U85 : NAND2_X1 port map( A1 => E(8), A2 => n140, ZN => n214);
   U86 : NAND2_X1 port map( A1 => B(8), A2 => n146, ZN => n213);
   U87 : NAND2_X1 port map( A1 => D(8), A2 => n152, ZN => n212);
   U88 : AOI22_X1 port map( A1 => C(8), A2 => n164, B1 => A(8), B2 => n158, ZN 
                           => n211);
   U89 : NAND4_X1 port map( A1 => n214, A2 => n213, A3 => n212, A4 => n211, ZN 
                           => Y(8));
   U90 : NAND2_X1 port map( A1 => E(9), A2 => n140, ZN => n218);
   U91 : NAND2_X1 port map( A1 => B(9), A2 => n146, ZN => n217);
   U92 : NAND2_X1 port map( A1 => D(9), A2 => n152, ZN => n216);
   U93 : AOI22_X1 port map( A1 => C(9), A2 => n164, B1 => A(9), B2 => n158, ZN 
                           => n215);
   U94 : NAND4_X1 port map( A1 => n218, A2 => n217, A3 => n216, A4 => n215, ZN 
                           => Y(9));
   U95 : NAND2_X1 port map( A1 => E(10), A2 => n140, ZN => n222);
   U96 : NAND2_X1 port map( A1 => B(10), A2 => n146, ZN => n221);
   U97 : NAND2_X1 port map( A1 => D(10), A2 => n152, ZN => n220);
   U98 : AOI22_X1 port map( A1 => C(10), A2 => n164, B1 => A(10), B2 => n158, 
                           ZN => n219);
   U99 : NAND4_X1 port map( A1 => n222, A2 => n221, A3 => n220, A4 => n219, ZN 
                           => Y(10));
   U100 : NAND2_X1 port map( A1 => E(11), A2 => n140, ZN => n226);
   U101 : NAND2_X1 port map( A1 => B(11), A2 => n146, ZN => n225);
   U102 : NAND2_X1 port map( A1 => D(11), A2 => n152, ZN => n224);
   U103 : AOI22_X1 port map( A1 => C(11), A2 => n164, B1 => A(11), B2 => n158, 
                           ZN => n223);
   U104 : NAND4_X1 port map( A1 => n226, A2 => n225, A3 => n224, A4 => n223, ZN
                           => Y(11));
   U105 : NAND2_X1 port map( A1 => E(12), A2 => n141, ZN => n230);
   U106 : NAND2_X1 port map( A1 => B(12), A2 => n147, ZN => n229);
   U107 : NAND2_X1 port map( A1 => D(12), A2 => n153, ZN => n228);
   U108 : AOI22_X1 port map( A1 => C(12), A2 => n165, B1 => A(12), B2 => n159, 
                           ZN => n227);
   U109 : NAND4_X1 port map( A1 => n230, A2 => n229, A3 => n228, A4 => n227, ZN
                           => Y(12));
   U110 : NAND2_X1 port map( A1 => E(13), A2 => n141, ZN => n234);
   U111 : NAND2_X1 port map( A1 => B(13), A2 => n147, ZN => n233);
   U112 : NAND2_X1 port map( A1 => D(13), A2 => n153, ZN => n232);
   U113 : AOI22_X1 port map( A1 => C(13), A2 => n165, B1 => A(13), B2 => n159, 
                           ZN => n231);
   U114 : NAND4_X1 port map( A1 => n234, A2 => n233, A3 => n232, A4 => n231, ZN
                           => Y(13));
   U115 : NAND2_X1 port map( A1 => E(14), A2 => n141, ZN => n238);
   U116 : NAND2_X1 port map( A1 => B(14), A2 => n147, ZN => n237);
   U117 : NAND2_X1 port map( A1 => D(14), A2 => n153, ZN => n236);
   U118 : AOI22_X1 port map( A1 => C(14), A2 => n165, B1 => A(14), B2 => n159, 
                           ZN => n235);
   U119 : NAND4_X1 port map( A1 => n238, A2 => n237, A3 => n236, A4 => n235, ZN
                           => Y(14));
   U120 : NAND2_X1 port map( A1 => E(15), A2 => n141, ZN => n242);
   U121 : NAND2_X1 port map( A1 => B(15), A2 => n147, ZN => n241);
   U122 : NAND2_X1 port map( A1 => D(15), A2 => n153, ZN => n240);
   U123 : AOI22_X1 port map( A1 => C(15), A2 => n165, B1 => A(15), B2 => n159, 
                           ZN => n239);
   U124 : NAND4_X1 port map( A1 => n242, A2 => n241, A3 => n240, A4 => n239, ZN
                           => Y(15));
   U125 : NAND2_X1 port map( A1 => E(16), A2 => n141, ZN => n246);
   U126 : NAND2_X1 port map( A1 => B(16), A2 => n147, ZN => n245);
   U127 : NAND2_X1 port map( A1 => D(16), A2 => n153, ZN => n244);
   U128 : AOI22_X1 port map( A1 => C(16), A2 => n165, B1 => A(16), B2 => n159, 
                           ZN => n243);
   U129 : NAND4_X1 port map( A1 => n246, A2 => n245, A3 => n244, A4 => n243, ZN
                           => Y(16));
   U130 : NAND2_X1 port map( A1 => E(17), A2 => n141, ZN => n250);
   U131 : NAND2_X1 port map( A1 => B(17), A2 => n147, ZN => n249);
   U132 : NAND2_X1 port map( A1 => D(17), A2 => n153, ZN => n248);
   U133 : AOI22_X1 port map( A1 => C(17), A2 => n165, B1 => A(17), B2 => n159, 
                           ZN => n247);
   U134 : NAND4_X1 port map( A1 => n250, A2 => n249, A3 => n248, A4 => n247, ZN
                           => Y(17));
   U135 : NAND2_X1 port map( A1 => E(18), A2 => n141, ZN => n254);
   U136 : NAND2_X1 port map( A1 => B(18), A2 => n147, ZN => n253);
   U137 : NAND2_X1 port map( A1 => D(18), A2 => n153, ZN => n252);
   U138 : AOI22_X1 port map( A1 => C(18), A2 => n165, B1 => A(18), B2 => n159, 
                           ZN => n251);
   U139 : NAND4_X1 port map( A1 => n254, A2 => n253, A3 => n252, A4 => n251, ZN
                           => Y(18));
   U140 : NAND2_X1 port map( A1 => E(19), A2 => n141, ZN => n258);
   U141 : NAND2_X1 port map( A1 => B(19), A2 => n147, ZN => n257);
   U142 : NAND2_X1 port map( A1 => D(19), A2 => n153, ZN => n256);
   U143 : AOI22_X1 port map( A1 => C(19), A2 => n165, B1 => A(19), B2 => n159, 
                           ZN => n255);
   U144 : NAND4_X1 port map( A1 => n258, A2 => n257, A3 => n256, A4 => n255, ZN
                           => Y(19));
   U145 : NAND2_X1 port map( A1 => E(20), A2 => n141, ZN => n262);
   U146 : NAND2_X1 port map( A1 => B(20), A2 => n147, ZN => n261);
   U147 : NAND2_X1 port map( A1 => D(20), A2 => n153, ZN => n260);
   U148 : AOI22_X1 port map( A1 => C(20), A2 => n165, B1 => A(20), B2 => n159, 
                           ZN => n259);
   U149 : NAND4_X1 port map( A1 => n262, A2 => n261, A3 => n260, A4 => n259, ZN
                           => Y(20));
   U150 : NAND2_X1 port map( A1 => E(21), A2 => n141, ZN => n266);
   U151 : NAND2_X1 port map( A1 => B(21), A2 => n147, ZN => n265);
   U152 : NAND2_X1 port map( A1 => D(21), A2 => n153, ZN => n264);
   U153 : AOI22_X1 port map( A1 => C(21), A2 => n165, B1 => A(21), B2 => n159, 
                           ZN => n263);
   U154 : NAND4_X1 port map( A1 => n266, A2 => n265, A3 => n264, A4 => n263, ZN
                           => Y(21));
   U155 : NAND2_X1 port map( A1 => E(22), A2 => n141, ZN => n270);
   U156 : NAND2_X1 port map( A1 => B(22), A2 => n147, ZN => n269);
   U157 : NAND2_X1 port map( A1 => D(22), A2 => n153, ZN => n268);
   U158 : AOI22_X1 port map( A1 => C(22), A2 => n165, B1 => A(22), B2 => n159, 
                           ZN => n267);
   U159 : NAND4_X1 port map( A1 => n270, A2 => n269, A3 => n268, A4 => n267, ZN
                           => Y(22));
   U160 : NAND2_X1 port map( A1 => E(23), A2 => n141, ZN => n274);
   U161 : NAND2_X1 port map( A1 => B(23), A2 => n147, ZN => n273);
   U162 : NAND2_X1 port map( A1 => D(23), A2 => n153, ZN => n272);
   U163 : AOI22_X1 port map( A1 => C(23), A2 => n165, B1 => A(23), B2 => n159, 
                           ZN => n271);
   U164 : NAND4_X1 port map( A1 => n274, A2 => n273, A3 => n272, A4 => n271, ZN
                           => Y(23));
   U165 : NAND2_X1 port map( A1 => E(24), A2 => n142, ZN => n278);
   U166 : NAND2_X1 port map( A1 => B(24), A2 => n148, ZN => n277);
   U167 : NAND2_X1 port map( A1 => D(24), A2 => n154, ZN => n276);
   U168 : AOI22_X1 port map( A1 => C(24), A2 => n166, B1 => A(24), B2 => n160, 
                           ZN => n275);
   U169 : NAND4_X1 port map( A1 => n278, A2 => n277, A3 => n276, A4 => n275, ZN
                           => Y(24));
   U170 : NAND2_X1 port map( A1 => E(25), A2 => n142, ZN => n282);
   U171 : NAND2_X1 port map( A1 => B(25), A2 => n148, ZN => n281);
   U172 : NAND2_X1 port map( A1 => D(25), A2 => n154, ZN => n280);
   U173 : AOI22_X1 port map( A1 => C(25), A2 => n166, B1 => A(25), B2 => n160, 
                           ZN => n279);
   U174 : NAND4_X1 port map( A1 => n282, A2 => n281, A3 => n280, A4 => n279, ZN
                           => Y(25));
   U175 : NAND2_X1 port map( A1 => E(26), A2 => n142, ZN => n286);
   U176 : NAND2_X1 port map( A1 => B(26), A2 => n148, ZN => n285);
   U177 : NAND2_X1 port map( A1 => D(26), A2 => n154, ZN => n284);
   U178 : AOI22_X1 port map( A1 => C(26), A2 => n166, B1 => A(26), B2 => n160, 
                           ZN => n283);
   U179 : NAND4_X1 port map( A1 => n286, A2 => n285, A3 => n284, A4 => n283, ZN
                           => Y(26));
   U180 : NAND2_X1 port map( A1 => E(27), A2 => n142, ZN => n290);
   U181 : NAND2_X1 port map( A1 => B(27), A2 => n148, ZN => n289);
   U182 : NAND2_X1 port map( A1 => D(27), A2 => n154, ZN => n288);
   U183 : AOI22_X1 port map( A1 => C(27), A2 => n166, B1 => A(27), B2 => n160, 
                           ZN => n287);
   U184 : NAND4_X1 port map( A1 => n290, A2 => n289, A3 => n288, A4 => n287, ZN
                           => Y(27));
   U185 : NAND2_X1 port map( A1 => E(28), A2 => n142, ZN => n294);
   U186 : NAND2_X1 port map( A1 => B(28), A2 => n148, ZN => n293);
   U187 : NAND2_X1 port map( A1 => D(28), A2 => n154, ZN => n292);
   U188 : AOI22_X1 port map( A1 => C(28), A2 => n166, B1 => A(28), B2 => n160, 
                           ZN => n291);
   U189 : NAND4_X1 port map( A1 => n294, A2 => n293, A3 => n292, A4 => n291, ZN
                           => Y(28));
   U190 : NAND2_X1 port map( A1 => E(29), A2 => n142, ZN => n298);
   U191 : NAND2_X1 port map( A1 => B(29), A2 => n148, ZN => n297);
   U192 : NAND2_X1 port map( A1 => D(29), A2 => n154, ZN => n296);
   U193 : AOI22_X1 port map( A1 => C(29), A2 => n166, B1 => A(29), B2 => n160, 
                           ZN => n295);
   U194 : NAND4_X1 port map( A1 => n298, A2 => n297, A3 => n296, A4 => n295, ZN
                           => Y(29));
   U195 : NAND2_X1 port map( A1 => E(30), A2 => n142, ZN => n302);
   U196 : NAND2_X1 port map( A1 => B(30), A2 => n148, ZN => n301);
   U197 : NAND2_X1 port map( A1 => D(30), A2 => n154, ZN => n300);
   U198 : AOI22_X1 port map( A1 => C(30), A2 => n166, B1 => A(30), B2 => n160, 
                           ZN => n299);
   U199 : NAND4_X1 port map( A1 => n302, A2 => n301, A3 => n300, A4 => n299, ZN
                           => Y(30));
   U200 : NAND2_X1 port map( A1 => E(31), A2 => n142, ZN => n306);
   U201 : NAND2_X1 port map( A1 => B(31), A2 => n148, ZN => n305);
   U202 : NAND2_X1 port map( A1 => D(31), A2 => n154, ZN => n304);
   U203 : AOI22_X1 port map( A1 => C(31), A2 => n166, B1 => A(31), B2 => n160, 
                           ZN => n303);
   U204 : NAND4_X1 port map( A1 => n306, A2 => n305, A3 => n304, A4 => n303, ZN
                           => Y(31));
   U205 : NAND2_X1 port map( A1 => E(32), A2 => n142, ZN => n310);
   U206 : NAND2_X1 port map( A1 => B(32), A2 => n148, ZN => n309);
   U207 : NAND2_X1 port map( A1 => D(32), A2 => n154, ZN => n308);
   U208 : AOI22_X1 port map( A1 => C(32), A2 => n166, B1 => A(32), B2 => n160, 
                           ZN => n307);
   U209 : NAND4_X1 port map( A1 => n310, A2 => n309, A3 => n308, A4 => n307, ZN
                           => Y(32));
   U210 : NAND2_X1 port map( A1 => E(33), A2 => n142, ZN => n314);
   U211 : NAND2_X1 port map( A1 => B(33), A2 => n148, ZN => n313);
   U212 : NAND2_X1 port map( A1 => D(33), A2 => n154, ZN => n312);
   U213 : AOI22_X1 port map( A1 => C(33), A2 => n166, B1 => A(33), B2 => n160, 
                           ZN => n311);
   U214 : NAND4_X1 port map( A1 => n314, A2 => n313, A3 => n312, A4 => n311, ZN
                           => Y(33));
   U215 : NAND2_X1 port map( A1 => E(34), A2 => n142, ZN => n318);
   U216 : NAND2_X1 port map( A1 => B(34), A2 => n148, ZN => n317);
   U217 : NAND2_X1 port map( A1 => D(34), A2 => n154, ZN => n316);
   U218 : AOI22_X1 port map( A1 => C(34), A2 => n166, B1 => A(34), B2 => n160, 
                           ZN => n315);
   U219 : NAND4_X1 port map( A1 => n318, A2 => n317, A3 => n316, A4 => n315, ZN
                           => Y(34));
   U220 : NAND2_X1 port map( A1 => E(35), A2 => n142, ZN => n322);
   U221 : NAND2_X1 port map( A1 => B(35), A2 => n148, ZN => n321);
   U222 : NAND2_X1 port map( A1 => D(35), A2 => n154, ZN => n320);
   U223 : AOI22_X1 port map( A1 => C(35), A2 => n166, B1 => A(35), B2 => n160, 
                           ZN => n319);
   U224 : NAND4_X1 port map( A1 => n322, A2 => n321, A3 => n320, A4 => n319, ZN
                           => Y(35));
   U225 : NAND2_X1 port map( A1 => E(36), A2 => n143, ZN => n326);
   U226 : NAND2_X1 port map( A1 => B(36), A2 => n149, ZN => n325);
   U227 : NAND2_X1 port map( A1 => D(36), A2 => n155, ZN => n324);
   U228 : AOI22_X1 port map( A1 => C(36), A2 => n167, B1 => A(36), B2 => n161, 
                           ZN => n323);
   U229 : NAND4_X1 port map( A1 => n326, A2 => n325, A3 => n324, A4 => n323, ZN
                           => Y(36));
   U230 : NAND2_X1 port map( A1 => E(37), A2 => n143, ZN => n330);
   U231 : NAND2_X1 port map( A1 => B(37), A2 => n149, ZN => n329);
   U232 : NAND2_X1 port map( A1 => D(37), A2 => n155, ZN => n328);
   U233 : AOI22_X1 port map( A1 => C(37), A2 => n167, B1 => A(37), B2 => n161, 
                           ZN => n327);
   U234 : NAND4_X1 port map( A1 => n330, A2 => n329, A3 => n328, A4 => n327, ZN
                           => Y(37));
   U235 : NAND2_X1 port map( A1 => E(38), A2 => n143, ZN => n334);
   U236 : NAND2_X1 port map( A1 => B(38), A2 => n149, ZN => n333);
   U237 : NAND2_X1 port map( A1 => D(38), A2 => n155, ZN => n332);
   U238 : AOI22_X1 port map( A1 => C(38), A2 => n167, B1 => A(38), B2 => n161, 
                           ZN => n331);
   U239 : NAND4_X1 port map( A1 => n334, A2 => n333, A3 => n332, A4 => n331, ZN
                           => Y(38));
   U240 : NAND2_X1 port map( A1 => E(39), A2 => n143, ZN => n338);
   U241 : NAND2_X1 port map( A1 => B(39), A2 => n149, ZN => n337);
   U242 : NAND2_X1 port map( A1 => D(39), A2 => n155, ZN => n336);
   U243 : AOI22_X1 port map( A1 => C(39), A2 => n167, B1 => A(39), B2 => n161, 
                           ZN => n335);
   U244 : NAND4_X1 port map( A1 => n338, A2 => n337, A3 => n336, A4 => n335, ZN
                           => Y(39));
   U245 : NAND2_X1 port map( A1 => E(40), A2 => n143, ZN => n342);
   U246 : NAND2_X1 port map( A1 => B(40), A2 => n149, ZN => n341);
   U247 : NAND2_X1 port map( A1 => D(40), A2 => n155, ZN => n340);
   U248 : AOI22_X1 port map( A1 => C(40), A2 => n167, B1 => A(40), B2 => n161, 
                           ZN => n339);
   U249 : NAND4_X1 port map( A1 => n342, A2 => n341, A3 => n340, A4 => n339, ZN
                           => Y(40));
   U250 : NAND2_X1 port map( A1 => E(41), A2 => n143, ZN => n346);
   U251 : NAND2_X1 port map( A1 => B(41), A2 => n149, ZN => n345);
   U252 : NAND2_X1 port map( A1 => D(41), A2 => n155, ZN => n344);
   U253 : AOI22_X1 port map( A1 => C(41), A2 => n167, B1 => A(41), B2 => n161, 
                           ZN => n343);
   U254 : NAND4_X1 port map( A1 => n346, A2 => n345, A3 => n344, A4 => n343, ZN
                           => Y(41));
   U255 : NAND2_X1 port map( A1 => E(42), A2 => n143, ZN => n350);
   U256 : NAND2_X1 port map( A1 => B(42), A2 => n149, ZN => n349);
   U257 : NAND2_X1 port map( A1 => D(42), A2 => n155, ZN => n348);
   U258 : AOI22_X1 port map( A1 => C(42), A2 => n167, B1 => A(42), B2 => n161, 
                           ZN => n347);
   U259 : NAND4_X1 port map( A1 => n350, A2 => n349, A3 => n348, A4 => n347, ZN
                           => Y(42));
   U260 : NAND2_X1 port map( A1 => E(43), A2 => n143, ZN => n354);
   U261 : NAND2_X1 port map( A1 => B(43), A2 => n149, ZN => n353);
   U262 : NAND2_X1 port map( A1 => D(43), A2 => n155, ZN => n352);
   U263 : AOI22_X1 port map( A1 => C(43), A2 => n167, B1 => A(43), B2 => n161, 
                           ZN => n351);
   U264 : NAND4_X1 port map( A1 => n354, A2 => n353, A3 => n352, A4 => n351, ZN
                           => Y(43));
   U265 : NAND2_X1 port map( A1 => E(44), A2 => n143, ZN => n358);
   U266 : NAND2_X1 port map( A1 => B(44), A2 => n149, ZN => n357);
   U267 : NAND2_X1 port map( A1 => D(44), A2 => n155, ZN => n356);
   U268 : AOI22_X1 port map( A1 => C(44), A2 => n167, B1 => A(44), B2 => n161, 
                           ZN => n355);
   U269 : NAND4_X1 port map( A1 => n358, A2 => n357, A3 => n356, A4 => n355, ZN
                           => Y(44));
   U270 : NAND2_X1 port map( A1 => E(45), A2 => n143, ZN => n362);
   U271 : NAND2_X1 port map( A1 => B(45), A2 => n149, ZN => n361);
   U272 : NAND2_X1 port map( A1 => D(45), A2 => n155, ZN => n360);
   U273 : AOI22_X1 port map( A1 => C(45), A2 => n167, B1 => A(45), B2 => n161, 
                           ZN => n359);
   U274 : NAND4_X1 port map( A1 => n362, A2 => n361, A3 => n360, A4 => n359, ZN
                           => Y(45));
   U275 : NAND2_X1 port map( A1 => E(46), A2 => n143, ZN => n366);
   U276 : NAND2_X1 port map( A1 => B(46), A2 => n149, ZN => n365);
   U277 : NAND2_X1 port map( A1 => D(46), A2 => n155, ZN => n364);
   U278 : AOI22_X1 port map( A1 => C(46), A2 => n167, B1 => A(46), B2 => n161, 
                           ZN => n363);
   U279 : NAND4_X1 port map( A1 => n366, A2 => n365, A3 => n364, A4 => n363, ZN
                           => Y(46));
   U280 : NAND2_X1 port map( A1 => E(47), A2 => n143, ZN => n370);
   U281 : NAND2_X1 port map( A1 => B(47), A2 => n149, ZN => n369);
   U282 : NAND2_X1 port map( A1 => D(47), A2 => n155, ZN => n368);
   U283 : AOI22_X1 port map( A1 => C(47), A2 => n167, B1 => A(47), B2 => n161, 
                           ZN => n367);
   U284 : NAND4_X1 port map( A1 => n370, A2 => n369, A3 => n368, A4 => n367, ZN
                           => Y(47));
   U285 : NAND2_X1 port map( A1 => E(48), A2 => n144, ZN => n374);
   U286 : NAND2_X1 port map( A1 => B(48), A2 => n150, ZN => n373);
   U287 : NAND2_X1 port map( A1 => D(48), A2 => n156, ZN => n372);
   U288 : AOI22_X1 port map( A1 => C(48), A2 => n168, B1 => A(48), B2 => n162, 
                           ZN => n371);
   U289 : NAND4_X1 port map( A1 => n374, A2 => n373, A3 => n372, A4 => n371, ZN
                           => Y(48));
   U290 : NAND2_X1 port map( A1 => E(49), A2 => n144, ZN => n378);
   U291 : NAND2_X1 port map( A1 => B(49), A2 => n150, ZN => n377);
   U292 : NAND2_X1 port map( A1 => D(49), A2 => n156, ZN => n376);
   U293 : AOI22_X1 port map( A1 => C(49), A2 => n168, B1 => A(49), B2 => n162, 
                           ZN => n375);
   U294 : NAND4_X1 port map( A1 => n378, A2 => n377, A3 => n376, A4 => n375, ZN
                           => Y(49));
   U295 : NAND2_X1 port map( A1 => E(50), A2 => n144, ZN => n382);
   U296 : NAND2_X1 port map( A1 => B(50), A2 => n150, ZN => n381);
   U297 : NAND2_X1 port map( A1 => D(50), A2 => n156, ZN => n380);
   U298 : AOI22_X1 port map( A1 => C(50), A2 => n168, B1 => A(50), B2 => n162, 
                           ZN => n379);
   U299 : NAND4_X1 port map( A1 => n382, A2 => n381, A3 => n380, A4 => n379, ZN
                           => Y(50));
   U300 : NAND2_X1 port map( A1 => E(51), A2 => n144, ZN => n386);
   U301 : NAND2_X1 port map( A1 => B(51), A2 => n150, ZN => n385);
   U302 : NAND2_X1 port map( A1 => D(51), A2 => n156, ZN => n384);
   U303 : AOI22_X1 port map( A1 => C(51), A2 => n168, B1 => A(51), B2 => n162, 
                           ZN => n383);
   U304 : NAND4_X1 port map( A1 => n386, A2 => n385, A3 => n384, A4 => n383, ZN
                           => Y(51));
   U305 : NAND2_X1 port map( A1 => E(52), A2 => n144, ZN => n390);
   U306 : NAND2_X1 port map( A1 => B(52), A2 => n150, ZN => n389);
   U307 : NAND2_X1 port map( A1 => D(52), A2 => n156, ZN => n388);
   U308 : AOI22_X1 port map( A1 => C(52), A2 => n168, B1 => A(52), B2 => n162, 
                           ZN => n387);
   U309 : NAND4_X1 port map( A1 => n390, A2 => n389, A3 => n388, A4 => n387, ZN
                           => Y(52));
   U310 : NAND2_X1 port map( A1 => E(53), A2 => n144, ZN => n394);
   U311 : NAND2_X1 port map( A1 => B(53), A2 => n150, ZN => n393);
   U312 : NAND2_X1 port map( A1 => D(53), A2 => n156, ZN => n392);
   U313 : AOI22_X1 port map( A1 => C(53), A2 => n168, B1 => A(53), B2 => n162, 
                           ZN => n391);
   U314 : NAND4_X1 port map( A1 => n394, A2 => n393, A3 => n392, A4 => n391, ZN
                           => Y(53));
   U315 : NAND2_X1 port map( A1 => E(54), A2 => n144, ZN => n398);
   U316 : NAND2_X1 port map( A1 => B(54), A2 => n150, ZN => n397);
   U317 : NAND2_X1 port map( A1 => D(54), A2 => n156, ZN => n396);
   U318 : AOI22_X1 port map( A1 => C(54), A2 => n168, B1 => A(54), B2 => n162, 
                           ZN => n395);
   U319 : NAND4_X1 port map( A1 => n398, A2 => n397, A3 => n396, A4 => n395, ZN
                           => Y(54));
   U320 : NAND2_X1 port map( A1 => E(55), A2 => n144, ZN => n402);
   U321 : NAND2_X1 port map( A1 => B(55), A2 => n150, ZN => n401);
   U322 : NAND2_X1 port map( A1 => D(55), A2 => n156, ZN => n400);
   U323 : AOI22_X1 port map( A1 => C(55), A2 => n168, B1 => A(55), B2 => n162, 
                           ZN => n399);
   U324 : NAND4_X1 port map( A1 => n402, A2 => n401, A3 => n400, A4 => n399, ZN
                           => Y(55));
   U325 : NAND2_X1 port map( A1 => E(56), A2 => n144, ZN => n406);
   U326 : NAND2_X1 port map( A1 => B(56), A2 => n150, ZN => n405);
   U327 : NAND2_X1 port map( A1 => D(56), A2 => n156, ZN => n404);
   U328 : AOI22_X1 port map( A1 => C(56), A2 => n168, B1 => A(56), B2 => n162, 
                           ZN => n403);
   U329 : NAND4_X1 port map( A1 => n406, A2 => n405, A3 => n404, A4 => n403, ZN
                           => Y(56));
   U330 : NAND2_X1 port map( A1 => E(57), A2 => n144, ZN => n410);
   U331 : NAND2_X1 port map( A1 => B(57), A2 => n150, ZN => n409);
   U332 : NAND2_X1 port map( A1 => D(57), A2 => n156, ZN => n408);
   U333 : AOI22_X1 port map( A1 => C(57), A2 => n168, B1 => A(57), B2 => n162, 
                           ZN => n407);
   U334 : NAND4_X1 port map( A1 => n410, A2 => n409, A3 => n408, A4 => n407, ZN
                           => Y(57));
   U335 : NAND2_X1 port map( A1 => E(58), A2 => n144, ZN => n414);
   U336 : NAND2_X1 port map( A1 => B(58), A2 => n150, ZN => n413);
   U337 : NAND2_X1 port map( A1 => D(58), A2 => n156, ZN => n412);
   U338 : AOI22_X1 port map( A1 => C(58), A2 => n168, B1 => A(58), B2 => n162, 
                           ZN => n411);
   U339 : NAND4_X1 port map( A1 => n414, A2 => n413, A3 => n412, A4 => n411, ZN
                           => Y(58));
   U340 : NAND2_X1 port map( A1 => E(59), A2 => n144, ZN => n418);
   U341 : NAND2_X1 port map( A1 => B(59), A2 => n150, ZN => n417);
   U342 : NAND2_X1 port map( A1 => D(59), A2 => n156, ZN => n416);
   U343 : AOI22_X1 port map( A1 => C(59), A2 => n168, B1 => A(59), B2 => n162, 
                           ZN => n415);
   U344 : NAND4_X1 port map( A1 => n418, A2 => n417, A3 => n416, A4 => n415, ZN
                           => Y(59));
   U345 : NAND2_X1 port map( A1 => E(60), A2 => n145, ZN => n422);
   U346 : NAND2_X1 port map( A1 => B(60), A2 => n151, ZN => n421);
   U347 : NAND2_X1 port map( A1 => D(60), A2 => n157, ZN => n420);
   U348 : AOI22_X1 port map( A1 => C(60), A2 => n169, B1 => A(60), B2 => n163, 
                           ZN => n419);
   U349 : NAND4_X1 port map( A1 => n422, A2 => n421, A3 => n420, A4 => n419, ZN
                           => Y(60));
   U350 : NAND2_X1 port map( A1 => E(61), A2 => n145, ZN => n426);
   U351 : NAND2_X1 port map( A1 => B(61), A2 => n151, ZN => n425);
   U352 : NAND2_X1 port map( A1 => D(61), A2 => n157, ZN => n424);
   U353 : AOI22_X1 port map( A1 => C(61), A2 => n169, B1 => A(61), B2 => n163, 
                           ZN => n423);
   U354 : NAND4_X1 port map( A1 => n426, A2 => n425, A3 => n424, A4 => n423, ZN
                           => Y(61));
   U355 : NAND2_X1 port map( A1 => E(62), A2 => n145, ZN => n430);
   U356 : NAND2_X1 port map( A1 => B(62), A2 => n151, ZN => n429);
   U357 : NAND2_X1 port map( A1 => D(62), A2 => n157, ZN => n428);
   U358 : AOI22_X1 port map( A1 => C(62), A2 => n169, B1 => A(62), B2 => n163, 
                           ZN => n427);
   U359 : NAND4_X1 port map( A1 => n430, A2 => n429, A3 => n428, A4 => n427, ZN
                           => Y(62));
   U360 : NAND2_X1 port map( A1 => E(63), A2 => n145, ZN => n438);
   U361 : NAND2_X1 port map( A1 => B(63), A2 => n151, ZN => n437);
   U362 : NAND2_X1 port map( A1 => D(63), A2 => n157, ZN => n436);
   U363 : AOI22_X1 port map( A1 => C(63), A2 => n169, B1 => A(63), B2 => n163, 
                           ZN => n435);
   U364 : NAND4_X1 port map( A1 => n438, A2 => n437, A3 => n436, A4 => n435, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_19 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_19;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7, n8, n9, n10, n11, n12, n14 : std_logic;

begin
   
   U1 : OR2_X1 port map( A1 => I(1), A2 => I(0), ZN => n9);
   U2 : MUX2_X2 port map( A => n5, B => n6, S => I(2), Z => O(1));
   U3 : AND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n5);
   U4 : AND2_X1 port map( A1 => n12, A2 => n14, ZN => n6);
   U5 : AOI21_X1 port map( B1 => n10, B2 => n14, A => I(2), ZN => O(0));
   U6 : INV_X1 port map( A => I(1), ZN => n7);
   U7 : INV_X1 port map( A => I(0), ZN => n8);
   U8 : AND3_X2 port map( A1 => n10, A2 => I(2), A3 => n11, ZN => O(2));
   U9 : NAND2_X1 port map( A1 => n9, A2 => n14, ZN => n10);
   U10 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n11);
   U11 : NAND2_X1 port map( A1 => n7, A2 => n8, ZN => n12);
   U12 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n14);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_18 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_18;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n4, n5, n6, n7, n9, n10, n11 : std_logic;

begin
   
   U1 : BUF_X1 port map( A => n11, Z => n4);
   U2 : NAND2_X1 port map( A1 => n5, A2 => n6, ZN => n7);
   U3 : NAND2_X1 port map( A1 => n7, A2 => n11, ZN => n10);
   U4 : INV_X1 port map( A => I(0), ZN => n5);
   U5 : INV_X1 port map( A => I(1), ZN => n6);
   U6 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n11);
   U7 : AND3_X1 port map( A1 => n4, A2 => I(2), A3 => n10, ZN => O(2));
   U8 : AOI21_X1 port map( B1 => n10, B2 => n4, A => I(2), ZN => O(0));
   U9 : MUX2_X1 port map( A => n4, B => n10, S => I(2), Z => n9);
   U10 : INV_X1 port map( A => n9, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_17 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_17;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_16 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_16;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_15 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_15;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_14 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_14;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_13 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_13;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_12 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_12;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_11 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_11;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_10 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_10;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_9 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_9;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_8 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_8;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_7 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_7;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_6 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_6;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_5 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_5;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n5, n6, n7 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => I(0), B2 => I(1), A => n7, ZN => n6);
   U2 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n7);
   U3 : AND3_X1 port map( A1 => n7, A2 => I(2), A3 => n6, ZN => O(2));
   U4 : AOI21_X1 port map( B1 => n7, B2 => n6, A => I(2), ZN => O(0));
   U5 : MUX2_X1 port map( A => n7, B => n6, S => I(2), Z => n5);
   U6 : INV_X1 port map( A => n5, ZN => O(1));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net148457, net148418, net138085, net138084, n3 : std_logic;

begin
   
   U1 : OAI21_X1 port map( B1 => n3, B2 => net138084, A => net138085, ZN => Co)
                           ;
   U2 : NAND2_X1 port map( A1 => net148418, A2 => net148457, ZN => net138085);
   U3 : CLKBUF_X1 port map( A => B, Z => net148457);
   U4 : CLKBUF_X1 port map( A => A, Z => net148418);
   U5 : INV_X1 port map( A => Ci, ZN => net138084);
   U6 : XNOR2_X1 port map( A => A, B => B, ZN => n3);
   U7 : XNOR2_X1 port map( A => n3, B => Ci, ZN => S);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTHMUL_N32_DW01_add_0 is

   port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (63 downto 0);  CO : out std_logic);

end BOOTHMUL_N32_DW01_add_0;

architecture SYN_rpl of BOOTHMUL_N32_DW01_add_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal carry_61_port, carry_60_port, carry_59_port, carry_58_port, 
      carry_57_port, carry_56_port, carry_55_port, carry_54_port, carry_53_port
      , carry_52_port, carry_51_port, carry_50_port, carry_49_port, 
      carry_48_port, carry_47_port, carry_46_port, carry_45_port, carry_44_port
      , carry_43_port, carry_42_port, carry_41_port, carry_40_port, 
      carry_39_port, carry_38_port, carry_37_port, carry_36_port, carry_35_port
      , carry_34_port, carry_33_port, carry_32_port, carry_31_port, 
      carry_30_port, carry_29_port, carry_28_port, carry_27_port, carry_26_port
      , carry_25_port, carry_24_port, carry_23_port, carry_22_port, 
      carry_21_port, carry_20_port, carry_19_port, carry_18_port, carry_17_port
      , carry_16_port, carry_15_port, carry_14_port, carry_13_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port, carry_3_port, 
      carry_2_port, carry_1_port, carry_62_port, n1 : std_logic;

begin
   
   U7 : XOR2_X1 port map( A => A(60), B => carry_60_port, Z => SUM(60));
   U9 : XOR2_X1 port map( A => A(59), B => carry_59_port, Z => SUM(59));
   U11 : XOR2_X1 port map( A => A(58), B => carry_58_port, Z => SUM(58));
   U13 : XOR2_X1 port map( A => A(57), B => carry_57_port, Z => SUM(57));
   U15 : XOR2_X1 port map( A => A(56), B => carry_56_port, Z => SUM(56));
   U17 : XOR2_X1 port map( A => A(55), B => carry_55_port, Z => SUM(55));
   U19 : XOR2_X1 port map( A => A(54), B => carry_54_port, Z => SUM(54));
   U21 : XOR2_X1 port map( A => A(53), B => carry_53_port, Z => SUM(53));
   U23 : XOR2_X1 port map( A => A(52), B => carry_52_port, Z => SUM(52));
   U25 : XOR2_X1 port map( A => A(51), B => carry_51_port, Z => SUM(51));
   U27 : XOR2_X1 port map( A => A(50), B => carry_50_port, Z => SUM(50));
   U29 : XOR2_X1 port map( A => A(49), B => carry_49_port, Z => SUM(49));
   U31 : XOR2_X1 port map( A => A(48), B => carry_48_port, Z => SUM(48));
   U33 : XOR2_X1 port map( A => A(47), B => carry_47_port, Z => SUM(47));
   U35 : XOR2_X1 port map( A => A(46), B => carry_46_port, Z => SUM(46));
   U37 : XOR2_X1 port map( A => A(45), B => carry_45_port, Z => SUM(45));
   U39 : XOR2_X1 port map( A => A(44), B => carry_44_port, Z => SUM(44));
   U41 : XOR2_X1 port map( A => A(43), B => carry_43_port, Z => SUM(43));
   U43 : XOR2_X1 port map( A => A(42), B => carry_42_port, Z => SUM(42));
   U45 : XOR2_X1 port map( A => A(41), B => carry_41_port, Z => SUM(41));
   U47 : XOR2_X1 port map( A => A(40), B => carry_40_port, Z => SUM(40));
   U49 : XOR2_X1 port map( A => A(39), B => carry_39_port, Z => SUM(39));
   U51 : XOR2_X1 port map( A => A(38), B => carry_38_port, Z => SUM(38));
   U53 : XOR2_X1 port map( A => A(37), B => carry_37_port, Z => SUM(37));
   U55 : XOR2_X1 port map( A => A(36), B => carry_36_port, Z => SUM(36));
   U57 : XOR2_X1 port map( A => A(35), B => carry_35_port, Z => SUM(35));
   U59 : XOR2_X1 port map( A => A(34), B => carry_34_port, Z => SUM(34));
   U61 : XOR2_X1 port map( A => A(33), B => carry_33_port, Z => SUM(33));
   U63 : XOR2_X1 port map( A => A(32), B => carry_32_port, Z => SUM(32));
   U65 : XOR2_X1 port map( A => A(31), B => carry_31_port, Z => SUM(31));
   U67 : XOR2_X1 port map( A => A(30), B => carry_30_port, Z => SUM(30));
   U69 : XOR2_X1 port map( A => A(29), B => carry_29_port, Z => SUM(29));
   U71 : XOR2_X1 port map( A => A(28), B => carry_28_port, Z => SUM(28));
   U73 : XOR2_X1 port map( A => A(27), B => carry_27_port, Z => SUM(27));
   U75 : XOR2_X1 port map( A => A(26), B => carry_26_port, Z => SUM(26));
   U77 : XOR2_X1 port map( A => A(25), B => carry_25_port, Z => SUM(25));
   U79 : XOR2_X1 port map( A => A(24), B => carry_24_port, Z => SUM(24));
   U81 : XOR2_X1 port map( A => A(23), B => carry_23_port, Z => SUM(23));
   U83 : XOR2_X1 port map( A => A(22), B => carry_22_port, Z => SUM(22));
   U85 : XOR2_X1 port map( A => A(21), B => carry_21_port, Z => SUM(21));
   U87 : XOR2_X1 port map( A => A(20), B => carry_20_port, Z => SUM(20));
   U89 : XOR2_X1 port map( A => A(19), B => carry_19_port, Z => SUM(19));
   U91 : XOR2_X1 port map( A => A(18), B => carry_18_port, Z => SUM(18));
   U93 : XOR2_X1 port map( A => A(17), B => carry_17_port, Z => SUM(17));
   U95 : XOR2_X1 port map( A => A(16), B => carry_16_port, Z => SUM(16));
   U97 : XOR2_X1 port map( A => A(15), B => carry_15_port, Z => SUM(15));
   U99 : XOR2_X1 port map( A => A(14), B => carry_14_port, Z => SUM(14));
   U101 : XOR2_X1 port map( A => A(13), B => carry_13_port, Z => SUM(13));
   U103 : XOR2_X1 port map( A => A(12), B => carry_12_port, Z => SUM(12));
   U105 : XOR2_X1 port map( A => A(11), B => carry_11_port, Z => SUM(11));
   U107 : XOR2_X1 port map( A => A(10), B => carry_10_port, Z => SUM(10));
   U109 : XOR2_X1 port map( A => A(9), B => carry_9_port, Z => SUM(9));
   U111 : XOR2_X1 port map( A => A(8), B => carry_8_port, Z => SUM(8));
   U113 : XOR2_X1 port map( A => A(7), B => carry_7_port, Z => SUM(7));
   U115 : XOR2_X1 port map( A => A(6), B => carry_6_port, Z => SUM(6));
   U117 : XOR2_X1 port map( A => A(5), B => carry_5_port, Z => SUM(5));
   U119 : XOR2_X1 port map( A => A(4), B => carry_4_port, Z => SUM(4));
   U121 : XOR2_X1 port map( A => A(3), B => carry_3_port, Z => SUM(3));
   U123 : XOR2_X1 port map( A => A(2), B => carry_2_port, Z => SUM(2));
   U125 : XOR2_X1 port map( A => A(1), B => carry_1_port, Z => SUM(1));
   U127 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));
   U5 : XOR2_X1 port map( A => A(61), B => carry_61_port, Z => SUM(61));
   U3 : XOR2_X1 port map( A => carry_62_port, B => A(62), Z => SUM(62));
   U1 : AND2_X1 port map( A1 => A(61), A2 => carry_61_port, ZN => carry_62_port
                           );
   U2 : XNOR2_X1 port map( A => A(63), B => n1, ZN => SUM(63));
   U4 : NAND2_X1 port map( A1 => carry_62_port, A2 => A(62), ZN => n1);
   U6 : AND2_X1 port map( A1 => carry_57_port, A2 => A(57), ZN => carry_58_port
                           );
   U8 : AND2_X1 port map( A1 => A(56), A2 => carry_56_port, ZN => carry_57_port
                           );
   U10 : AND2_X1 port map( A1 => A(54), A2 => carry_54_port, ZN => 
                           carry_55_port);
   U12 : AND2_X1 port map( A1 => A(55), A2 => carry_55_port, ZN => 
                           carry_56_port);
   U14 : AND2_X1 port map( A1 => carry_53_port, A2 => A(53), ZN => 
                           carry_54_port);
   U16 : AND2_X1 port map( A1 => carry_52_port, A2 => A(52), ZN => 
                           carry_53_port);
   U18 : AND2_X1 port map( A1 => carry_51_port, A2 => A(51), ZN => 
                           carry_52_port);
   U20 : AND2_X1 port map( A1 => A(50), A2 => carry_50_port, ZN => 
                           carry_51_port);
   U22 : AND2_X1 port map( A1 => carry_49_port, A2 => A(49), ZN => 
                           carry_50_port);
   U24 : AND2_X1 port map( A1 => carry_46_port, A2 => A(46), ZN => 
                           carry_47_port);
   U26 : AND2_X1 port map( A1 => carry_41_port, A2 => A(41), ZN => 
                           carry_42_port);
   U28 : AND2_X1 port map( A1 => carry_40_port, A2 => A(40), ZN => 
                           carry_41_port);
   U30 : AND2_X1 port map( A1 => carry_39_port, A2 => A(39), ZN => 
                           carry_40_port);
   U32 : AND2_X1 port map( A1 => carry_37_port, A2 => A(37), ZN => 
                           carry_38_port);
   U34 : AND2_X1 port map( A1 => carry_35_port, A2 => A(35), ZN => 
                           carry_36_port);
   U36 : AND2_X1 port map( A1 => carry_25_port, A2 => A(25), ZN => 
                           carry_26_port);
   U38 : AND2_X1 port map( A1 => carry_24_port, A2 => A(24), ZN => 
                           carry_25_port);
   U40 : AND2_X1 port map( A1 => carry_60_port, A2 => A(60), ZN => 
                           carry_61_port);
   U42 : AND2_X1 port map( A1 => A(58), A2 => carry_58_port, ZN => 
                           carry_59_port);
   U44 : AND2_X1 port map( A1 => carry_59_port, A2 => A(59), ZN => 
                           carry_60_port);
   U46 : AND2_X1 port map( A1 => carry_48_port, A2 => A(48), ZN => 
                           carry_49_port);
   U48 : AND2_X1 port map( A1 => A(47), A2 => carry_47_port, ZN => 
                           carry_48_port);
   U50 : AND2_X1 port map( A1 => carry_45_port, A2 => A(45), ZN => 
                           carry_46_port);
   U52 : AND2_X1 port map( A1 => carry_44_port, A2 => A(44), ZN => 
                           carry_45_port);
   U54 : AND2_X1 port map( A1 => carry_43_port, A2 => A(43), ZN => 
                           carry_44_port);
   U56 : AND2_X1 port map( A1 => carry_42_port, A2 => A(42), ZN => 
                           carry_43_port);
   U58 : AND2_X1 port map( A1 => carry_38_port, A2 => A(38), ZN => 
                           carry_39_port);
   U60 : AND2_X1 port map( A1 => carry_36_port, A2 => A(36), ZN => 
                           carry_37_port);
   U62 : AND2_X1 port map( A1 => carry_34_port, A2 => A(34), ZN => 
                           carry_35_port);
   U64 : AND2_X1 port map( A1 => carry_33_port, A2 => A(33), ZN => 
                           carry_34_port);
   U66 : AND2_X1 port map( A1 => carry_32_port, A2 => A(32), ZN => 
                           carry_33_port);
   U68 : AND2_X1 port map( A1 => carry_31_port, A2 => A(31), ZN => 
                           carry_32_port);
   U70 : AND2_X1 port map( A1 => carry_29_port, A2 => A(29), ZN => 
                           carry_30_port);
   U72 : AND2_X1 port map( A1 => carry_30_port, A2 => A(30), ZN => 
                           carry_31_port);
   U74 : AND2_X1 port map( A1 => carry_28_port, A2 => A(28), ZN => 
                           carry_29_port);
   U76 : AND2_X1 port map( A1 => carry_27_port, A2 => A(27), ZN => 
                           carry_28_port);
   U78 : AND2_X1 port map( A1 => carry_26_port, A2 => A(26), ZN => 
                           carry_27_port);
   U80 : AND2_X1 port map( A1 => carry_23_port, A2 => A(23), ZN => 
                           carry_24_port);
   U82 : AND2_X1 port map( A1 => carry_22_port, A2 => A(22), ZN => 
                           carry_23_port);
   U84 : AND2_X1 port map( A1 => carry_21_port, A2 => A(21), ZN => 
                           carry_22_port);
   U86 : AND2_X1 port map( A1 => carry_20_port, A2 => A(20), ZN => 
                           carry_21_port);
   U88 : AND2_X1 port map( A1 => carry_19_port, A2 => A(19), ZN => 
                           carry_20_port);
   U90 : AND2_X1 port map( A1 => carry_18_port, A2 => A(18), ZN => 
                           carry_19_port);
   U92 : AND2_X1 port map( A1 => carry_17_port, A2 => A(17), ZN => 
                           carry_18_port);
   U94 : AND2_X1 port map( A1 => carry_16_port, A2 => A(16), ZN => 
                           carry_17_port);
   U96 : AND2_X1 port map( A1 => carry_15_port, A2 => A(15), ZN => 
                           carry_16_port);
   U98 : AND2_X1 port map( A1 => carry_14_port, A2 => A(14), ZN => 
                           carry_15_port);
   U100 : AND2_X1 port map( A1 => carry_13_port, A2 => A(13), ZN => 
                           carry_14_port);
   U102 : AND2_X1 port map( A1 => carry_12_port, A2 => A(12), ZN => 
                           carry_13_port);
   U104 : AND2_X1 port map( A1 => carry_11_port, A2 => A(11), ZN => 
                           carry_12_port);
   U106 : AND2_X1 port map( A1 => carry_10_port, A2 => A(10), ZN => 
                           carry_11_port);
   U108 : AND2_X1 port map( A1 => carry_9_port, A2 => A(9), ZN => carry_10_port
                           );
   U110 : AND2_X1 port map( A1 => carry_8_port, A2 => A(8), ZN => carry_9_port)
                           ;
   U112 : AND2_X1 port map( A1 => carry_7_port, A2 => A(7), ZN => carry_8_port)
                           ;
   U114 : AND2_X1 port map( A1 => carry_6_port, A2 => A(6), ZN => carry_7_port)
                           ;
   U116 : AND2_X1 port map( A1 => carry_5_port, A2 => A(5), ZN => carry_6_port)
                           ;
   U118 : AND2_X1 port map( A1 => carry_4_port, A2 => A(4), ZN => carry_5_port)
                           ;
   U120 : AND2_X1 port map( A1 => carry_3_port, A2 => A(3), ZN => carry_4_port)
                           ;
   U122 : AND2_X1 port map( A1 => carry_2_port, A2 => A(2), ZN => carry_3_port)
                           ;
   U124 : AND2_X1 port map( A1 => carry_1_port, A2 => A(1), ZN => carry_2_port)
                           ;
   U126 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => carry_1_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity RCA_generic_N64_0 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_generic_N64_0;

architecture SYN_STRUCTURAL of RCA_generic_N64_0 is

   component FA_945
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_946
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_947
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_948
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_949
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_950
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_951
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_952
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_953
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_954
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_955
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_956
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_957
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_958
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_959
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_960
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_961
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_962
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_963
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_964
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_965
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_966
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_967
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_968
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_969
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_970
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_971
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_972
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_973
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_974
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_975
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_976
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_977
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_978
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_979
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_980
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_981
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_982
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_983
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_984
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_985
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_986
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_987
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_988
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_989
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_990
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_991
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_992
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_993
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_994
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_995
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_996
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_997
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_998
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_999
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1000
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1001
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1002
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1003
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1004
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1005
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1006
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_1007
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_63_port, CTMP_62_port, CTMP_61_port, CTMP_60_port, CTMP_59_port,
      CTMP_58_port, CTMP_57_port, CTMP_56_port, CTMP_55_port, CTMP_54_port, 
      CTMP_53_port, CTMP_52_port, CTMP_51_port, CTMP_50_port, CTMP_49_port, 
      CTMP_48_port, CTMP_47_port, CTMP_46_port, CTMP_45_port, CTMP_44_port, 
      CTMP_43_port, CTMP_42_port, CTMP_41_port, CTMP_40_port, CTMP_39_port, 
      CTMP_38_port, CTMP_37_port, CTMP_36_port, CTMP_35_port, CTMP_34_port, 
      CTMP_33_port, CTMP_32_port, CTMP_31_port, CTMP_30_port, CTMP_29_port, 
      CTMP_28_port, CTMP_27_port, CTMP_26_port, CTMP_25_port, CTMP_24_port, 
      CTMP_23_port, CTMP_22_port, CTMP_21_port, CTMP_20_port, CTMP_19_port, 
      CTMP_18_port, CTMP_17_port, CTMP_16_port, CTMP_15_port, CTMP_14_port, 
      CTMP_13_port, CTMP_12_port, CTMP_11_port, CTMP_10_port, CTMP_9_port, 
      CTMP_8_port, CTMP_7_port, CTMP_6_port, CTMP_5_port, CTMP_4_port, 
      CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   FAI_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   FAI_2 : FA_1007 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1)
                           , Co => CTMP_2_port);
   FAI_3 : FA_1006 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2)
                           , Co => CTMP_3_port);
   FAI_4 : FA_1005 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3)
                           , Co => CTMP_4_port);
   FAI_5 : FA_1004 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4)
                           , Co => CTMP_5_port);
   FAI_6 : FA_1003 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5)
                           , Co => CTMP_6_port);
   FAI_7 : FA_1002 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6)
                           , Co => CTMP_7_port);
   FAI_8 : FA_1001 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7)
                           , Co => CTMP_8_port);
   FAI_9 : FA_1000 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8)
                           , Co => CTMP_9_port);
   FAI_10 : FA_999 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9)
                           , Co => CTMP_10_port);
   FAI_11 : FA_998 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   FAI_12 : FA_997 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   FAI_13 : FA_996 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   FAI_14 : FA_995 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   FAI_15 : FA_994 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   FAI_16 : FA_993 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   FAI_17 : FA_992 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   FAI_18 : FA_991 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   FAI_19 : FA_990 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   FAI_20 : FA_989 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   FAI_21 : FA_988 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   FAI_22 : FA_987 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   FAI_23 : FA_986 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   FAI_24 : FA_985 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   FAI_25 : FA_984 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   FAI_26 : FA_983 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   FAI_27 : FA_982 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   FAI_28 : FA_981 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   FAI_29 : FA_980 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   FAI_30 : FA_979 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   FAI_31 : FA_978 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   FAI_32 : FA_977 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => CTMP_32_port);
   FAI_33 : FA_976 port map( A => A(32), B => B(32), Ci => CTMP_32_port, S => 
                           S(32), Co => CTMP_33_port);
   FAI_34 : FA_975 port map( A => A(33), B => B(33), Ci => CTMP_33_port, S => 
                           S(33), Co => CTMP_34_port);
   FAI_35 : FA_974 port map( A => A(34), B => B(34), Ci => CTMP_34_port, S => 
                           S(34), Co => CTMP_35_port);
   FAI_36 : FA_973 port map( A => A(35), B => B(35), Ci => CTMP_35_port, S => 
                           S(35), Co => CTMP_36_port);
   FAI_37 : FA_972 port map( A => A(36), B => B(36), Ci => CTMP_36_port, S => 
                           S(36), Co => CTMP_37_port);
   FAI_38 : FA_971 port map( A => A(37), B => B(37), Ci => CTMP_37_port, S => 
                           S(37), Co => CTMP_38_port);
   FAI_39 : FA_970 port map( A => A(38), B => B(38), Ci => CTMP_38_port, S => 
                           S(38), Co => CTMP_39_port);
   FAI_40 : FA_969 port map( A => A(39), B => B(39), Ci => CTMP_39_port, S => 
                           S(39), Co => CTMP_40_port);
   FAI_41 : FA_968 port map( A => A(40), B => B(40), Ci => CTMP_40_port, S => 
                           S(40), Co => CTMP_41_port);
   FAI_42 : FA_967 port map( A => A(41), B => B(41), Ci => CTMP_41_port, S => 
                           S(41), Co => CTMP_42_port);
   FAI_43 : FA_966 port map( A => A(42), B => B(42), Ci => CTMP_42_port, S => 
                           S(42), Co => CTMP_43_port);
   FAI_44 : FA_965 port map( A => A(43), B => B(43), Ci => CTMP_43_port, S => 
                           S(43), Co => CTMP_44_port);
   FAI_45 : FA_964 port map( A => A(44), B => B(44), Ci => CTMP_44_port, S => 
                           S(44), Co => CTMP_45_port);
   FAI_46 : FA_963 port map( A => A(45), B => B(45), Ci => CTMP_45_port, S => 
                           S(45), Co => CTMP_46_port);
   FAI_47 : FA_962 port map( A => A(46), B => B(46), Ci => CTMP_46_port, S => 
                           S(46), Co => CTMP_47_port);
   FAI_48 : FA_961 port map( A => A(47), B => B(47), Ci => CTMP_47_port, S => 
                           S(47), Co => CTMP_48_port);
   FAI_49 : FA_960 port map( A => A(48), B => B(48), Ci => CTMP_48_port, S => 
                           S(48), Co => CTMP_49_port);
   FAI_50 : FA_959 port map( A => A(49), B => B(49), Ci => CTMP_49_port, S => 
                           S(49), Co => CTMP_50_port);
   FAI_51 : FA_958 port map( A => A(50), B => B(50), Ci => CTMP_50_port, S => 
                           S(50), Co => CTMP_51_port);
   FAI_52 : FA_957 port map( A => A(51), B => B(51), Ci => CTMP_51_port, S => 
                           S(51), Co => CTMP_52_port);
   FAI_53 : FA_956 port map( A => A(52), B => B(52), Ci => CTMP_52_port, S => 
                           S(52), Co => CTMP_53_port);
   FAI_54 : FA_955 port map( A => A(53), B => B(53), Ci => CTMP_53_port, S => 
                           S(53), Co => CTMP_54_port);
   FAI_55 : FA_954 port map( A => A(54), B => B(54), Ci => CTMP_54_port, S => 
                           S(54), Co => CTMP_55_port);
   FAI_56 : FA_953 port map( A => A(55), B => B(55), Ci => CTMP_55_port, S => 
                           S(55), Co => CTMP_56_port);
   FAI_57 : FA_952 port map( A => A(56), B => B(56), Ci => CTMP_56_port, S => 
                           S(56), Co => CTMP_57_port);
   FAI_58 : FA_951 port map( A => A(57), B => B(57), Ci => CTMP_57_port, S => 
                           S(57), Co => CTMP_58_port);
   FAI_59 : FA_950 port map( A => A(58), B => B(58), Ci => CTMP_58_port, S => 
                           S(58), Co => CTMP_59_port);
   FAI_60 : FA_949 port map( A => A(59), B => B(59), Ci => CTMP_59_port, S => 
                           S(59), Co => CTMP_60_port);
   FAI_61 : FA_948 port map( A => A(60), B => B(60), Ci => CTMP_60_port, S => 
                           S(60), Co => CTMP_61_port);
   FAI_62 : FA_947 port map( A => A(61), B => B(61), Ci => CTMP_61_port, S => 
                           S(61), Co => CTMP_62_port);
   FAI_63 : FA_946 port map( A => A(62), B => B(62), Ci => CTMP_62_port, S => 
                           S(62), Co => CTMP_63_port);
   FAI_64 : FA_945 port map( A => A(63), B => B(63), Ci => CTMP_63_port, S => 
                           S(63), Co => Co);

end SYN_STRUCTURAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity MUX51_GENERIC_N64_0 is

   port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto 0)
         );

end MUX51_GENERIC_N64_0;

architecture SYN_BEHAVIORAL of MUX51_GENERIC_N64_0 is

   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X4
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal net142158, net142406, net145869, net145867, net145865, net145863, 
      net145879, net145875, net145893, net145891, net145889, net145887, 
      net145885, net145903, net145901, net145899, net145897, net145917, 
      net145915, net145909, net148517, net148599, net158795, net157198, 
      net148598, net145883, net142411, net142410, net142409, net149357, 
      net148545, net148525, net148524, net142421, net142420, net142417, 
      net142415, net142414, net142412, net142408, net149341, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, 
      n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, 
      n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, 
      n202, n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, 
      n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, 
      n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, 
      n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, 
      n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, 
      n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, 
      n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, 
      n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, 
      n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, 
      n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, 
      n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, 
      n334, n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345, 
      n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, 
      n358, n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, 
      n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, 
      n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393, 
      n394, n395 : std_logic;

begin
   
   U1 : BUF_X2 port map( A => n142, Z => net145903);
   U2 : INV_X1 port map( A => net142412, ZN => n139);
   U3 : CLKBUF_X1 port map( A => SEL(0), Z => net149357);
   U4 : BUF_X1 port map( A => n140, Z => net145875);
   U5 : AND2_X1 port map( A1 => net142420, A2 => net142417, ZN => n140);
   U6 : OR2_X1 port map( A1 => net148525, A2 => n143, ZN => n144);
   U7 : CLKBUF_X1 port map( A => SEL(1), Z => n141);
   U8 : INV_X1 port map( A => net142415, ZN => n142);
   U9 : CLKBUF_X1 port map( A => net142158, Z => net145897);
   U10 : AND2_X1 port map( A1 => net157198, A2 => E(0), ZN => net149341);
   U11 : NAND2_X1 port map( A1 => net148545, A2 => net149341, ZN => net142408);
   U12 : AND4_X1 port map( A1 => net157198, A2 => net142415, A3 => net142412, 
                           A4 => net142414, ZN => net148517);
   U13 : INV_X1 port map( A => n144, ZN => net148599);
   U14 : INV_X1 port map( A => SEL(1), ZN => n143);
   U15 : OR2_X1 port map( A1 => n143, A2 => net148525, ZN => net157198);
   U16 : NAND3_X1 port map( A1 => n143, A2 => net149357, A3 => net142421, ZN =>
                           net142415);
   U17 : AND3_X1 port map( A1 => SEL(1), A2 => net149357, A3 => net142421, ZN 
                           => net158795);
   U18 : NAND3_X1 port map( A1 => n141, A2 => net149357, A3 => net142421, ZN =>
                           net142414);
   U19 : NOR2_X1 port map( A1 => SEL(2), A2 => SEL(1), ZN => net142420);
   U20 : NAND4_X1 port map( A1 => net142408, A2 => net142411, A3 => net142410, 
                           A4 => net142409, ZN => Y(0));
   U21 : AND3_X1 port map( A1 => net142415, A2 => net142412, A3 => net142414, 
                           ZN => net148545);
   U22 : INV_X1 port map( A => SEL(2), ZN => net142421);
   U23 : INV_X1 port map( A => net142415, ZN => net142158);
   U24 : NAND2_X1 port map( A1 => net142420, A2 => net142417, ZN => net142412);
   U25 : INV_X1 port map( A => SEL(0), ZN => net142417);
   U26 : NAND2_X1 port map( A1 => net142417, A2 => net148524, ZN => net148525);
   U27 : INV_X1 port map( A => SEL(2), ZN => net148524);
   U28 : NAND2_X1 port map( A1 => B(0), A2 => net142158, ZN => net142409);
   U29 : NAND2_X1 port map( A1 => D(0), A2 => net145883, ZN => net142410);
   U30 : BUF_X1 port map( A => net158795, Z => net145883);
   U31 : NAND2_X1 port map( A1 => D(1), A2 => net145883, ZN => net142406);
   U32 : AOI22_X1 port map( A1 => net148598, A2 => C(0), B1 => n139, B2 => A(0)
                           , ZN => net142411);
   U33 : INV_X1 port map( A => n144, ZN => net148598);
   U34 : CLKBUF_X1 port map( A => net148599, Z => net145867);
   U35 : BUF_X4 port map( A => net148599, Z => net145865);
   U36 : CLKBUF_X3 port map( A => net148517, Z => net145909);
   U37 : BUF_X4 port map( A => n140, Z => net145879);
   U38 : BUF_X1 port map( A => net158795, Z => net145885);
   U39 : BUF_X1 port map( A => net158795, Z => net145887);
   U40 : CLKBUF_X2 port map( A => net148517, Z => net145915);
   U41 : CLKBUF_X1 port map( A => n142, Z => net145901);
   U42 : CLKBUF_X1 port map( A => net158795, Z => net145889);
   U43 : CLKBUF_X1 port map( A => net158795, Z => net145891);
   U44 : CLKBUF_X1 port map( A => n142, Z => net145899);
   U45 : CLKBUF_X1 port map( A => net148599, Z => net145863);
   U46 : CLKBUF_X1 port map( A => net148517, Z => net145917);
   U47 : CLKBUF_X1 port map( A => net158795, Z => net145893);
   U48 : CLKBUF_X1 port map( A => net148599, Z => net145869);
   U49 : NAND2_X1 port map( A1 => E(1), A2 => net148517, ZN => n147);
   U50 : NAND2_X1 port map( A1 => B(1), A2 => net142158, ZN => n146);
   U51 : AOI22_X1 port map( A1 => C(1), A2 => net148599, B1 => A(1), B2 => n140
                           , ZN => n145);
   U52 : NAND4_X1 port map( A1 => n147, A2 => n146, A3 => net142406, A4 => n145
                           , ZN => Y(1));
   U53 : NAND2_X1 port map( A1 => E(2), A2 => net145917, ZN => n151);
   U54 : NAND2_X1 port map( A1 => B(2), A2 => n142, ZN => n150);
   U55 : NAND2_X1 port map( A1 => D(2), A2 => net145887, ZN => n149);
   U56 : AOI22_X1 port map( A1 => C(2), A2 => net145867, B1 => A(2), B2 => n140
                           , ZN => n148);
   U57 : NAND4_X1 port map( A1 => n151, A2 => n150, A3 => n149, A4 => n148, ZN 
                           => Y(2));
   U58 : NAND2_X1 port map( A1 => E(3), A2 => net145909, ZN => n155);
   U59 : NAND2_X1 port map( A1 => B(3), A2 => net145897, ZN => n154);
   U60 : NAND2_X1 port map( A1 => D(3), A2 => net145885, ZN => n153);
   U61 : AOI22_X1 port map( A1 => C(3), A2 => net145863, B1 => A(3), B2 => 
                           net145875, ZN => n152);
   U62 : NAND4_X1 port map( A1 => n155, A2 => n154, A3 => n153, A4 => n152, ZN 
                           => Y(3));
   U63 : NAND2_X1 port map( A1 => E(4), A2 => net145909, ZN => n159);
   U64 : NAND2_X1 port map( A1 => B(4), A2 => net145899, ZN => n158);
   U65 : NAND2_X1 port map( A1 => D(4), A2 => net145893, ZN => n157);
   U66 : AOI22_X1 port map( A1 => C(4), A2 => net145863, B1 => A(4), B2 => 
                           net145875, ZN => n156);
   U67 : NAND4_X1 port map( A1 => n159, A2 => n158, A3 => n157, A4 => n156, ZN 
                           => Y(4));
   U68 : NAND2_X1 port map( A1 => E(5), A2 => net145909, ZN => n163);
   U69 : NAND2_X1 port map( A1 => B(5), A2 => net145901, ZN => n162);
   U70 : NAND2_X1 port map( A1 => D(5), A2 => net145891, ZN => n161);
   U71 : AOI22_X1 port map( A1 => C(5), A2 => net145865, B1 => A(5), B2 => 
                           net145875, ZN => n160);
   U72 : NAND4_X1 port map( A1 => n163, A2 => n162, A3 => n161, A4 => n160, ZN 
                           => Y(5));
   U73 : NAND2_X1 port map( A1 => E(6), A2 => net145915, ZN => n167);
   U74 : NAND2_X1 port map( A1 => B(6), A2 => net145903, ZN => n166);
   U75 : NAND2_X1 port map( A1 => D(6), A2 => net145889, ZN => n165);
   U76 : AOI22_X1 port map( A1 => C(6), A2 => net145869, B1 => A(6), B2 => 
                           net145875, ZN => n164);
   U77 : NAND4_X1 port map( A1 => n167, A2 => n166, A3 => n165, A4 => n164, ZN 
                           => Y(6));
   U78 : NAND2_X1 port map( A1 => E(7), A2 => net145915, ZN => n171);
   U79 : NAND2_X1 port map( A1 => B(7), A2 => net145903, ZN => n170);
   U80 : NAND2_X1 port map( A1 => D(7), A2 => net145887, ZN => n169);
   U81 : AOI22_X1 port map( A1 => C(7), A2 => net145865, B1 => A(7), B2 => 
                           net145875, ZN => n168);
   U82 : NAND4_X1 port map( A1 => n171, A2 => n170, A3 => n169, A4 => n168, ZN 
                           => Y(7));
   U83 : NAND2_X1 port map( A1 => E(8), A2 => net145915, ZN => n175);
   U84 : NAND2_X1 port map( A1 => B(8), A2 => net145903, ZN => n174);
   U85 : NAND2_X1 port map( A1 => D(8), A2 => net145885, ZN => n173);
   U86 : AOI22_X1 port map( A1 => C(8), A2 => net145865, B1 => A(8), B2 => 
                           net145879, ZN => n172);
   U87 : NAND4_X1 port map( A1 => n175, A2 => n174, A3 => n173, A4 => n172, ZN 
                           => Y(8));
   U88 : NAND2_X1 port map( A1 => E(9), A2 => net145915, ZN => n179);
   U89 : NAND2_X1 port map( A1 => B(9), A2 => net145903, ZN => n178);
   U90 : NAND2_X1 port map( A1 => D(9), A2 => net145893, ZN => n177);
   U91 : AOI22_X1 port map( A1 => C(9), A2 => net145865, B1 => A(9), B2 => 
                           net145879, ZN => n176);
   U92 : NAND4_X1 port map( A1 => n179, A2 => n178, A3 => n177, A4 => n176, ZN 
                           => Y(9));
   U93 : NAND2_X1 port map( A1 => E(10), A2 => net145915, ZN => n183);
   U94 : NAND2_X1 port map( A1 => B(10), A2 => net145903, ZN => n182);
   U95 : NAND2_X1 port map( A1 => D(10), A2 => net145891, ZN => n181);
   U96 : AOI22_X1 port map( A1 => C(10), A2 => net145865, B1 => A(10), B2 => 
                           net145879, ZN => n180);
   U97 : NAND4_X1 port map( A1 => n183, A2 => n182, A3 => n181, A4 => n180, ZN 
                           => Y(10));
   U98 : NAND2_X1 port map( A1 => E(11), A2 => net145915, ZN => n187);
   U99 : NAND2_X1 port map( A1 => B(11), A2 => net145903, ZN => n186);
   U100 : NAND2_X1 port map( A1 => D(11), A2 => net145889, ZN => n185);
   U101 : AOI22_X1 port map( A1 => C(11), A2 => net145865, B1 => A(11), B2 => 
                           net145879, ZN => n184);
   U102 : NAND4_X1 port map( A1 => n187, A2 => n186, A3 => n185, A4 => n184, ZN
                           => Y(11));
   U103 : NAND2_X1 port map( A1 => E(12), A2 => net145915, ZN => n191);
   U104 : NAND2_X1 port map( A1 => B(12), A2 => net145897, ZN => n190);
   U105 : NAND2_X1 port map( A1 => D(12), A2 => net145887, ZN => n189);
   U106 : AOI22_X1 port map( A1 => C(12), A2 => net145865, B1 => A(12), B2 => 
                           net145879, ZN => n188);
   U107 : NAND4_X1 port map( A1 => n191, A2 => n190, A3 => n189, A4 => n188, ZN
                           => Y(12));
   U108 : NAND2_X1 port map( A1 => E(13), A2 => net145915, ZN => n195);
   U109 : NAND2_X1 port map( A1 => B(13), A2 => net145897, ZN => n194);
   U110 : NAND2_X1 port map( A1 => D(13), A2 => net145885, ZN => n193);
   U111 : AOI22_X1 port map( A1 => C(13), A2 => net145865, B1 => A(13), B2 => 
                           net145879, ZN => n192);
   U112 : NAND4_X1 port map( A1 => n195, A2 => n194, A3 => n193, A4 => n192, ZN
                           => Y(13));
   U113 : NAND2_X1 port map( A1 => E(14), A2 => net145915, ZN => n199);
   U114 : NAND2_X1 port map( A1 => B(14), A2 => net145897, ZN => n198);
   U115 : NAND2_X1 port map( A1 => D(14), A2 => net145893, ZN => n197);
   U116 : AOI22_X1 port map( A1 => C(14), A2 => net145865, B1 => A(14), B2 => 
                           net145879, ZN => n196);
   U117 : NAND4_X1 port map( A1 => n199, A2 => n198, A3 => n197, A4 => n196, ZN
                           => Y(14));
   U118 : NAND2_X1 port map( A1 => E(15), A2 => net145915, ZN => n203);
   U119 : NAND2_X1 port map( A1 => B(15), A2 => net145897, ZN => n202);
   U120 : NAND2_X1 port map( A1 => D(15), A2 => net145891, ZN => n201);
   U121 : AOI22_X1 port map( A1 => C(15), A2 => net145865, B1 => A(15), B2 => 
                           net145879, ZN => n200);
   U122 : NAND4_X1 port map( A1 => n203, A2 => n202, A3 => n201, A4 => n200, ZN
                           => Y(15));
   U123 : NAND2_X1 port map( A1 => E(16), A2 => net145915, ZN => n207);
   U124 : NAND2_X1 port map( A1 => B(16), A2 => net145897, ZN => n206);
   U125 : NAND2_X1 port map( A1 => D(16), A2 => net145889, ZN => n205);
   U126 : AOI22_X1 port map( A1 => C(16), A2 => net145865, B1 => A(16), B2 => 
                           net145879, ZN => n204);
   U127 : NAND4_X1 port map( A1 => n207, A2 => n206, A3 => n205, A4 => n204, ZN
                           => Y(16));
   U128 : NAND2_X1 port map( A1 => E(17), A2 => net145915, ZN => n211);
   U129 : NAND2_X1 port map( A1 => B(17), A2 => net145897, ZN => n210);
   U130 : NAND2_X1 port map( A1 => D(17), A2 => net145887, ZN => n209);
   U131 : AOI22_X1 port map( A1 => C(17), A2 => net145865, B1 => A(17), B2 => 
                           net145879, ZN => n208);
   U132 : NAND4_X1 port map( A1 => n211, A2 => n210, A3 => n209, A4 => n208, ZN
                           => Y(17));
   U133 : NAND2_X1 port map( A1 => E(18), A2 => net145915, ZN => n215);
   U134 : NAND2_X1 port map( A1 => B(18), A2 => net145897, ZN => n214);
   U135 : NAND2_X1 port map( A1 => D(18), A2 => net145885, ZN => n213);
   U136 : AOI22_X1 port map( A1 => C(18), A2 => net145869, B1 => A(18), B2 => 
                           net145879, ZN => n212);
   U137 : NAND4_X1 port map( A1 => n215, A2 => n214, A3 => n213, A4 => n212, ZN
                           => Y(18));
   U138 : NAND2_X1 port map( A1 => E(19), A2 => net145915, ZN => n219);
   U139 : NAND2_X1 port map( A1 => B(19), A2 => net145897, ZN => n218);
   U140 : NAND2_X1 port map( A1 => D(19), A2 => net145893, ZN => n217);
   U141 : AOI22_X1 port map( A1 => C(19), A2 => net145869, B1 => A(19), B2 => 
                           net145879, ZN => n216);
   U142 : NAND4_X1 port map( A1 => n219, A2 => n218, A3 => n217, A4 => n216, ZN
                           => Y(19));
   U143 : NAND2_X1 port map( A1 => E(20), A2 => net145915, ZN => n223);
   U144 : NAND2_X1 port map( A1 => B(20), A2 => net145897, ZN => n222);
   U145 : NAND2_X1 port map( A1 => D(20), A2 => net145891, ZN => n221);
   U146 : AOI22_X1 port map( A1 => C(20), A2 => net145865, B1 => A(20), B2 => 
                           net145879, ZN => n220);
   U147 : NAND4_X1 port map( A1 => n223, A2 => n222, A3 => n221, A4 => n220, ZN
                           => Y(20));
   U148 : NAND2_X1 port map( A1 => E(21), A2 => net145915, ZN => n227);
   U149 : NAND2_X1 port map( A1 => B(21), A2 => net145897, ZN => n226);
   U150 : NAND2_X1 port map( A1 => D(21), A2 => net145889, ZN => n225);
   U151 : AOI22_X1 port map( A1 => C(21), A2 => net145869, B1 => A(21), B2 => 
                           net145879, ZN => n224);
   U152 : NAND4_X1 port map( A1 => n227, A2 => n226, A3 => n225, A4 => n224, ZN
                           => Y(21));
   U153 : NAND2_X1 port map( A1 => E(22), A2 => net145915, ZN => n231);
   U154 : NAND2_X1 port map( A1 => B(22), A2 => net145897, ZN => n230);
   U155 : NAND2_X1 port map( A1 => D(22), A2 => net145887, ZN => n229);
   U156 : AOI22_X1 port map( A1 => C(22), A2 => net145865, B1 => A(22), B2 => 
                           net145879, ZN => n228);
   U157 : NAND4_X1 port map( A1 => n231, A2 => n230, A3 => n229, A4 => n228, ZN
                           => Y(22));
   U158 : NAND2_X1 port map( A1 => E(23), A2 => net145915, ZN => n235);
   U159 : NAND2_X1 port map( A1 => B(23), A2 => net145897, ZN => n234);
   U160 : NAND2_X1 port map( A1 => D(23), A2 => net145885, ZN => n233);
   U161 : AOI22_X1 port map( A1 => C(23), A2 => net145869, B1 => A(23), B2 => 
                           net145879, ZN => n232);
   U162 : NAND4_X1 port map( A1 => n235, A2 => n234, A3 => n233, A4 => n232, ZN
                           => Y(23));
   U163 : NAND2_X1 port map( A1 => E(24), A2 => net145915, ZN => n239);
   U164 : NAND2_X1 port map( A1 => B(24), A2 => net145899, ZN => n238);
   U165 : NAND2_X1 port map( A1 => D(24), A2 => net145893, ZN => n237);
   U166 : AOI22_X1 port map( A1 => C(24), A2 => net145865, B1 => A(24), B2 => 
                           net145879, ZN => n236);
   U167 : NAND4_X1 port map( A1 => n239, A2 => n238, A3 => n237, A4 => n236, ZN
                           => Y(24));
   U168 : NAND2_X1 port map( A1 => E(25), A2 => net145915, ZN => n243);
   U169 : NAND2_X1 port map( A1 => B(25), A2 => net145899, ZN => n242);
   U170 : NAND2_X1 port map( A1 => D(25), A2 => net145891, ZN => n241);
   U171 : AOI22_X1 port map( A1 => C(25), A2 => net145869, B1 => A(25), B2 => 
                           net145879, ZN => n240);
   U172 : NAND4_X1 port map( A1 => n243, A2 => n242, A3 => n241, A4 => n240, ZN
                           => Y(25));
   U173 : NAND2_X1 port map( A1 => E(26), A2 => net145915, ZN => n247);
   U174 : NAND2_X1 port map( A1 => B(26), A2 => net145899, ZN => n246);
   U175 : NAND2_X1 port map( A1 => D(26), A2 => net145889, ZN => n245);
   U176 : AOI22_X1 port map( A1 => C(26), A2 => net145865, B1 => A(26), B2 => 
                           net145879, ZN => n244);
   U177 : NAND4_X1 port map( A1 => n247, A2 => n246, A3 => n245, A4 => n244, ZN
                           => Y(26));
   U178 : NAND2_X1 port map( A1 => E(27), A2 => net145915, ZN => n251);
   U179 : NAND2_X1 port map( A1 => B(27), A2 => net145899, ZN => n250);
   U180 : NAND2_X1 port map( A1 => D(27), A2 => net145887, ZN => n249);
   U181 : AOI22_X1 port map( A1 => C(27), A2 => net145869, B1 => A(27), B2 => 
                           net145879, ZN => n248);
   U182 : NAND4_X1 port map( A1 => n251, A2 => n250, A3 => n249, A4 => n248, ZN
                           => Y(27));
   U183 : NAND2_X1 port map( A1 => E(28), A2 => net145915, ZN => n255);
   U184 : NAND2_X1 port map( A1 => B(28), A2 => net145899, ZN => n254);
   U185 : NAND2_X1 port map( A1 => D(28), A2 => net145885, ZN => n253);
   U186 : AOI22_X1 port map( A1 => C(28), A2 => net145865, B1 => A(28), B2 => 
                           net145879, ZN => n252);
   U187 : NAND4_X1 port map( A1 => n255, A2 => n254, A3 => n253, A4 => n252, ZN
                           => Y(28));
   U188 : NAND2_X1 port map( A1 => E(29), A2 => net145915, ZN => n259);
   U189 : NAND2_X1 port map( A1 => B(29), A2 => net145899, ZN => n258);
   U190 : NAND2_X1 port map( A1 => D(29), A2 => net145893, ZN => n257);
   U191 : AOI22_X1 port map( A1 => C(29), A2 => net145869, B1 => A(29), B2 => 
                           net145879, ZN => n256);
   U192 : NAND4_X1 port map( A1 => n259, A2 => n258, A3 => n257, A4 => n256, ZN
                           => Y(29));
   U193 : NAND2_X1 port map( A1 => E(30), A2 => net145915, ZN => n263);
   U194 : NAND2_X1 port map( A1 => B(30), A2 => net145899, ZN => n262);
   U195 : NAND2_X1 port map( A1 => D(30), A2 => net145891, ZN => n261);
   U196 : AOI22_X1 port map( A1 => C(30), A2 => net145865, B1 => A(30), B2 => 
                           net145879, ZN => n260);
   U197 : NAND4_X1 port map( A1 => n263, A2 => n262, A3 => n261, A4 => n260, ZN
                           => Y(30));
   U198 : NAND2_X1 port map( A1 => E(31), A2 => net145915, ZN => n267);
   U199 : NAND2_X1 port map( A1 => B(31), A2 => net145899, ZN => n266);
   U200 : NAND2_X1 port map( A1 => D(31), A2 => net145889, ZN => n265);
   U201 : AOI22_X1 port map( A1 => C(31), A2 => net145869, B1 => A(31), B2 => 
                           net145879, ZN => n264);
   U202 : NAND4_X1 port map( A1 => n267, A2 => n266, A3 => n265, A4 => n264, ZN
                           => Y(31));
   U203 : NAND2_X1 port map( A1 => E(32), A2 => net145915, ZN => n271);
   U204 : NAND2_X1 port map( A1 => B(32), A2 => net145899, ZN => n270);
   U205 : NAND2_X1 port map( A1 => D(32), A2 => net145887, ZN => n269);
   U206 : AOI22_X1 port map( A1 => C(32), A2 => net145865, B1 => A(32), B2 => 
                           net145879, ZN => n268);
   U207 : NAND4_X1 port map( A1 => n271, A2 => n270, A3 => n269, A4 => n268, ZN
                           => Y(32));
   U208 : NAND2_X1 port map( A1 => E(33), A2 => net145909, ZN => n275);
   U209 : NAND2_X1 port map( A1 => B(33), A2 => net145899, ZN => n274);
   U210 : NAND2_X1 port map( A1 => D(33), A2 => net145885, ZN => n273);
   U211 : AOI22_X1 port map( A1 => C(33), A2 => net145869, B1 => A(33), B2 => 
                           net145879, ZN => n272);
   U212 : NAND4_X1 port map( A1 => n275, A2 => n274, A3 => n273, A4 => n272, ZN
                           => Y(33));
   U213 : NAND2_X1 port map( A1 => E(34), A2 => net145915, ZN => n279);
   U214 : NAND2_X1 port map( A1 => B(34), A2 => net145899, ZN => n278);
   U215 : NAND2_X1 port map( A1 => D(34), A2 => net145893, ZN => n277);
   U216 : AOI22_X1 port map( A1 => C(34), A2 => net145869, B1 => A(34), B2 => 
                           net145879, ZN => n276);
   U217 : NAND4_X1 port map( A1 => n279, A2 => n278, A3 => n277, A4 => n276, ZN
                           => Y(34));
   U218 : NAND2_X1 port map( A1 => E(35), A2 => net145909, ZN => n283);
   U219 : NAND2_X1 port map( A1 => B(35), A2 => net145899, ZN => n282);
   U220 : NAND2_X1 port map( A1 => D(35), A2 => net145891, ZN => n281);
   U221 : AOI22_X1 port map( A1 => C(35), A2 => net145865, B1 => A(35), B2 => 
                           net145879, ZN => n280);
   U222 : NAND4_X1 port map( A1 => n283, A2 => n282, A3 => n281, A4 => n280, ZN
                           => Y(35));
   U223 : NAND2_X1 port map( A1 => E(36), A2 => net145915, ZN => n287);
   U224 : NAND2_X1 port map( A1 => B(36), A2 => net145901, ZN => n286);
   U225 : NAND2_X1 port map( A1 => D(36), A2 => net145889, ZN => n285);
   U226 : AOI22_X1 port map( A1 => C(36), A2 => net145865, B1 => A(36), B2 => 
                           net145879, ZN => n284);
   U227 : NAND4_X1 port map( A1 => n287, A2 => n286, A3 => n285, A4 => n284, ZN
                           => Y(36));
   U228 : NAND2_X1 port map( A1 => E(37), A2 => net145909, ZN => n291);
   U229 : NAND2_X1 port map( A1 => B(37), A2 => net145901, ZN => n290);
   U230 : NAND2_X1 port map( A1 => D(37), A2 => net145887, ZN => n289);
   U231 : AOI22_X1 port map( A1 => C(37), A2 => net145865, B1 => A(37), B2 => 
                           net145879, ZN => n288);
   U232 : NAND4_X1 port map( A1 => n291, A2 => n290, A3 => n289, A4 => n288, ZN
                           => Y(37));
   U233 : NAND2_X1 port map( A1 => E(38), A2 => net145915, ZN => n295);
   U234 : NAND2_X1 port map( A1 => B(38), A2 => net145901, ZN => n294);
   U235 : NAND2_X1 port map( A1 => D(38), A2 => net145885, ZN => n293);
   U236 : AOI22_X1 port map( A1 => C(38), A2 => net145869, B1 => A(38), B2 => 
                           net145879, ZN => n292);
   U237 : NAND4_X1 port map( A1 => n295, A2 => n294, A3 => n293, A4 => n292, ZN
                           => Y(38));
   U238 : NAND2_X1 port map( A1 => E(39), A2 => net145909, ZN => n299);
   U239 : NAND2_X1 port map( A1 => B(39), A2 => net145901, ZN => n298);
   U240 : NAND2_X1 port map( A1 => D(39), A2 => net145893, ZN => n297);
   U241 : AOI22_X1 port map( A1 => C(39), A2 => net145865, B1 => A(39), B2 => 
                           net145879, ZN => n296);
   U242 : NAND4_X1 port map( A1 => n299, A2 => n298, A3 => n297, A4 => n296, ZN
                           => Y(39));
   U243 : NAND2_X1 port map( A1 => E(40), A2 => net145915, ZN => n303);
   U244 : NAND2_X1 port map( A1 => B(40), A2 => net145901, ZN => n302);
   U245 : NAND2_X1 port map( A1 => D(40), A2 => net145891, ZN => n301);
   U246 : AOI22_X1 port map( A1 => C(40), A2 => net145865, B1 => A(40), B2 => 
                           net145879, ZN => n300);
   U247 : NAND4_X1 port map( A1 => n303, A2 => n302, A3 => n301, A4 => n300, ZN
                           => Y(40));
   U248 : NAND2_X1 port map( A1 => E(41), A2 => net145909, ZN => n307);
   U249 : NAND2_X1 port map( A1 => B(41), A2 => net145901, ZN => n306);
   U250 : NAND2_X1 port map( A1 => D(41), A2 => net145889, ZN => n305);
   U251 : AOI22_X1 port map( A1 => C(41), A2 => net145865, B1 => A(41), B2 => 
                           net145879, ZN => n304);
   U252 : NAND4_X1 port map( A1 => n307, A2 => n306, A3 => n305, A4 => n304, ZN
                           => Y(41));
   U253 : NAND2_X1 port map( A1 => E(42), A2 => net145915, ZN => n311);
   U254 : NAND2_X1 port map( A1 => B(42), A2 => net145901, ZN => n310);
   U255 : NAND2_X1 port map( A1 => D(42), A2 => net145887, ZN => n309);
   U256 : AOI22_X1 port map( A1 => C(42), A2 => net145869, B1 => A(42), B2 => 
                           net145879, ZN => n308);
   U257 : NAND4_X1 port map( A1 => n311, A2 => n310, A3 => n309, A4 => n308, ZN
                           => Y(42));
   U258 : NAND2_X1 port map( A1 => E(43), A2 => net145909, ZN => n315);
   U259 : NAND2_X1 port map( A1 => B(43), A2 => net145901, ZN => n314);
   U260 : NAND2_X1 port map( A1 => D(43), A2 => net145885, ZN => n313);
   U261 : AOI22_X1 port map( A1 => C(43), A2 => net145865, B1 => A(43), B2 => 
                           net145879, ZN => n312);
   U262 : NAND4_X1 port map( A1 => n315, A2 => n314, A3 => n313, A4 => n312, ZN
                           => Y(43));
   U263 : NAND2_X1 port map( A1 => E(44), A2 => net145915, ZN => n319);
   U264 : NAND2_X1 port map( A1 => B(44), A2 => net145901, ZN => n318);
   U265 : NAND2_X1 port map( A1 => D(44), A2 => net145893, ZN => n317);
   U266 : AOI22_X1 port map( A1 => C(44), A2 => net145865, B1 => A(44), B2 => 
                           net145879, ZN => n316);
   U267 : NAND4_X1 port map( A1 => n319, A2 => n318, A3 => n317, A4 => n316, ZN
                           => Y(44));
   U268 : NAND2_X1 port map( A1 => E(45), A2 => net145915, ZN => n323);
   U269 : NAND2_X1 port map( A1 => B(45), A2 => net145901, ZN => n322);
   U270 : NAND2_X1 port map( A1 => D(45), A2 => net145891, ZN => n321);
   U271 : AOI22_X1 port map( A1 => C(45), A2 => net145869, B1 => A(45), B2 => 
                           net145879, ZN => n320);
   U272 : NAND4_X1 port map( A1 => n323, A2 => n322, A3 => n321, A4 => n320, ZN
                           => Y(45));
   U273 : NAND2_X1 port map( A1 => E(46), A2 => net145909, ZN => n327);
   U274 : NAND2_X1 port map( A1 => B(46), A2 => net145901, ZN => n326);
   U275 : NAND2_X1 port map( A1 => D(46), A2 => net145889, ZN => n325);
   U276 : AOI22_X1 port map( A1 => C(46), A2 => net145865, B1 => A(46), B2 => 
                           net145879, ZN => n324);
   U277 : NAND4_X1 port map( A1 => n327, A2 => n326, A3 => n325, A4 => n324, ZN
                           => Y(46));
   U278 : NAND2_X1 port map( A1 => E(47), A2 => net145909, ZN => n331);
   U279 : NAND2_X1 port map( A1 => B(47), A2 => net145901, ZN => n330);
   U280 : NAND2_X1 port map( A1 => D(47), A2 => net145887, ZN => n329);
   U281 : AOI22_X1 port map( A1 => C(47), A2 => net145865, B1 => A(47), B2 => 
                           net145875, ZN => n328);
   U282 : NAND4_X1 port map( A1 => n331, A2 => n330, A3 => n329, A4 => n328, ZN
                           => Y(47));
   U283 : NAND2_X1 port map( A1 => E(48), A2 => net145909, ZN => n335);
   U284 : NAND2_X1 port map( A1 => B(48), A2 => net145903, ZN => n334);
   U285 : NAND2_X1 port map( A1 => D(48), A2 => net145885, ZN => n333);
   U286 : AOI22_X1 port map( A1 => C(48), A2 => net145869, B1 => A(48), B2 => 
                           net145879, ZN => n332);
   U287 : NAND4_X1 port map( A1 => n335, A2 => n334, A3 => n333, A4 => n332, ZN
                           => Y(48));
   U288 : NAND2_X1 port map( A1 => E(49), A2 => net145909, ZN => n339);
   U289 : NAND2_X1 port map( A1 => B(49), A2 => net145903, ZN => n338);
   U290 : NAND2_X1 port map( A1 => D(49), A2 => net145893, ZN => n337);
   U291 : AOI22_X1 port map( A1 => C(49), A2 => net145865, B1 => A(49), B2 => 
                           net145879, ZN => n336);
   U292 : NAND4_X1 port map( A1 => n339, A2 => n338, A3 => n337, A4 => n336, ZN
                           => Y(49));
   U293 : NAND2_X1 port map( A1 => E(50), A2 => net145915, ZN => n343);
   U294 : NAND2_X1 port map( A1 => B(50), A2 => net145903, ZN => n342);
   U295 : NAND2_X1 port map( A1 => D(50), A2 => net145891, ZN => n341);
   U296 : AOI22_X1 port map( A1 => C(50), A2 => net145865, B1 => A(50), B2 => 
                           net145879, ZN => n340);
   U297 : NAND4_X1 port map( A1 => n343, A2 => n342, A3 => n341, A4 => n340, ZN
                           => Y(50));
   U298 : NAND2_X1 port map( A1 => E(51), A2 => net145909, ZN => n347);
   U299 : NAND2_X1 port map( A1 => B(51), A2 => net145903, ZN => n346);
   U300 : NAND2_X1 port map( A1 => D(51), A2 => net145889, ZN => n345);
   U301 : AOI22_X1 port map( A1 => C(51), A2 => net145869, B1 => A(51), B2 => 
                           net145879, ZN => n344);
   U302 : NAND4_X1 port map( A1 => n347, A2 => n346, A3 => n345, A4 => n344, ZN
                           => Y(51));
   U303 : NAND2_X1 port map( A1 => E(52), A2 => net145915, ZN => n351);
   U304 : NAND2_X1 port map( A1 => B(52), A2 => net145903, ZN => n350);
   U305 : NAND2_X1 port map( A1 => D(52), A2 => net145887, ZN => n349);
   U306 : AOI22_X1 port map( A1 => C(52), A2 => net145865, B1 => A(52), B2 => 
                           net145875, ZN => n348);
   U307 : NAND4_X1 port map( A1 => n351, A2 => n350, A3 => n349, A4 => n348, ZN
                           => Y(52));
   U308 : NAND2_X1 port map( A1 => E(53), A2 => net145915, ZN => n355);
   U309 : NAND2_X1 port map( A1 => B(53), A2 => net145903, ZN => n354);
   U310 : NAND2_X1 port map( A1 => D(53), A2 => net145885, ZN => n353);
   U311 : AOI22_X1 port map( A1 => C(53), A2 => net145865, B1 => A(53), B2 => 
                           net145879, ZN => n352);
   U312 : NAND4_X1 port map( A1 => n355, A2 => n354, A3 => n353, A4 => n352, ZN
                           => Y(53));
   U313 : NAND2_X1 port map( A1 => E(54), A2 => net145909, ZN => n359);
   U314 : NAND2_X1 port map( A1 => B(54), A2 => net145903, ZN => n358);
   U315 : NAND2_X1 port map( A1 => D(54), A2 => net145893, ZN => n357);
   U316 : AOI22_X1 port map( A1 => C(54), A2 => net145863, B1 => A(54), B2 => 
                           net145879, ZN => n356);
   U317 : NAND4_X1 port map( A1 => n359, A2 => n358, A3 => n357, A4 => n356, ZN
                           => Y(54));
   U318 : NAND2_X1 port map( A1 => E(55), A2 => net145915, ZN => n363);
   U319 : NAND2_X1 port map( A1 => B(55), A2 => net145903, ZN => n362);
   U320 : NAND2_X1 port map( A1 => D(55), A2 => net145891, ZN => n361);
   U321 : AOI22_X1 port map( A1 => C(55), A2 => net145865, B1 => A(55), B2 => 
                           net145879, ZN => n360);
   U322 : NAND4_X1 port map( A1 => n363, A2 => n362, A3 => n361, A4 => n360, ZN
                           => Y(55));
   U323 : NAND2_X1 port map( A1 => E(56), A2 => net145909, ZN => n367);
   U324 : NAND2_X1 port map( A1 => B(56), A2 => net145903, ZN => n366);
   U325 : NAND2_X1 port map( A1 => D(56), A2 => net145889, ZN => n365);
   U326 : AOI22_X1 port map( A1 => C(56), A2 => net145869, B1 => A(56), B2 => 
                           net145879, ZN => n364);
   U327 : NAND4_X1 port map( A1 => n367, A2 => n366, A3 => n365, A4 => n364, ZN
                           => Y(56));
   U328 : NAND2_X1 port map( A1 => E(57), A2 => net145915, ZN => n371);
   U329 : NAND2_X1 port map( A1 => B(57), A2 => net145903, ZN => n370);
   U330 : NAND2_X1 port map( A1 => D(57), A2 => net145887, ZN => n369);
   U331 : AOI22_X1 port map( A1 => C(57), A2 => net145865, B1 => A(57), B2 => 
                           net145879, ZN => n368);
   U332 : NAND4_X1 port map( A1 => n371, A2 => n370, A3 => n369, A4 => n368, ZN
                           => Y(57));
   U333 : NAND2_X1 port map( A1 => E(58), A2 => net145909, ZN => n375);
   U334 : NAND2_X1 port map( A1 => B(58), A2 => net145903, ZN => n374);
   U335 : NAND2_X1 port map( A1 => D(58), A2 => net145885, ZN => n373);
   U336 : AOI22_X1 port map( A1 => C(58), A2 => net145865, B1 => A(58), B2 => 
                           net145879, ZN => n372);
   U337 : NAND4_X1 port map( A1 => n375, A2 => n374, A3 => n373, A4 => n372, ZN
                           => Y(58));
   U338 : NAND2_X1 port map( A1 => E(59), A2 => net145915, ZN => n379);
   U339 : NAND2_X1 port map( A1 => B(59), A2 => net145903, ZN => n378);
   U340 : NAND2_X1 port map( A1 => D(59), A2 => net145893, ZN => n377);
   U341 : AOI22_X1 port map( A1 => C(59), A2 => net145863, B1 => A(59), B2 => 
                           net145875, ZN => n376);
   U342 : NAND4_X1 port map( A1 => n379, A2 => n378, A3 => n377, A4 => n376, ZN
                           => Y(59));
   U343 : NAND2_X1 port map( A1 => E(60), A2 => net145909, ZN => n383);
   U344 : NAND2_X1 port map( A1 => B(60), A2 => net145903, ZN => n382);
   U345 : NAND2_X1 port map( A1 => D(60), A2 => net145891, ZN => n381);
   U346 : AOI22_X1 port map( A1 => C(60), A2 => net145869, B1 => A(60), B2 => 
                           net145879, ZN => n380);
   U347 : NAND4_X1 port map( A1 => n383, A2 => n382, A3 => n381, A4 => n380, ZN
                           => Y(60));
   U348 : NAND2_X1 port map( A1 => E(61), A2 => net145915, ZN => n387);
   U349 : NAND2_X1 port map( A1 => B(61), A2 => net145903, ZN => n386);
   U350 : NAND2_X1 port map( A1 => D(61), A2 => net145889, ZN => n385);
   U351 : AOI22_X1 port map( A1 => C(61), A2 => net145863, B1 => A(61), B2 => 
                           net145879, ZN => n384);
   U352 : NAND4_X1 port map( A1 => n387, A2 => n386, A3 => n385, A4 => n384, ZN
                           => Y(61));
   U353 : NAND2_X1 port map( A1 => E(62), A2 => net145909, ZN => n391);
   U354 : NAND2_X1 port map( A1 => B(62), A2 => net145903, ZN => n390);
   U355 : NAND2_X1 port map( A1 => D(62), A2 => net145887, ZN => n389);
   U356 : AOI22_X1 port map( A1 => C(62), A2 => net145865, B1 => A(62), B2 => 
                           net145879, ZN => n388);
   U357 : NAND4_X1 port map( A1 => n391, A2 => n390, A3 => n389, A4 => n388, ZN
                           => Y(62));
   U358 : NAND2_X1 port map( A1 => E(63), A2 => net145915, ZN => n395);
   U359 : NAND2_X1 port map( A1 => B(63), A2 => net145901, ZN => n394);
   U360 : NAND2_X1 port map( A1 => D(63), A2 => net145885, ZN => n393);
   U361 : AOI22_X1 port map( A1 => C(63), A2 => net145865, B1 => A(63), B2 => 
                           net145879, ZN => n392);
   U362 : NAND4_X1 port map( A1 => n395, A2 => n394, A3 => n393, A4 => n392, ZN
                           => Y(63));

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTH_ENCODER_4 is

   port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
         downto 0));

end BOOTH_ENCODER_4;

architecture SYN_BEHAVIORAL of BOOTH_ENCODER_4 is

   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal net142483, net156612, net158600, net158612, net158610, net158606, 
      net158605, n4 : std_logic;

begin
   
   U1 : NAND2_X1 port map( A1 => net158610, A2 => net158612, ZN => net158606);
   U2 : INV_X1 port map( A => I(0), ZN => net158612);
   U3 : NAND2_X1 port map( A1 => I(1), A2 => I(0), ZN => n4);
   U4 : XNOR2_X1 port map( A => n4, B => I(2), ZN => net158605);
   U5 : AND2_X2 port map( A1 => net158605, A2 => net158606, ZN => O(1));
   U6 : INV_X1 port map( A => I(1), ZN => net158610);
   U7 : AOI21_X1 port map( B1 => net156612, B2 => net142483, A => I(2), ZN => 
                           O(0));
   U8 : AND3_X2 port map( A1 => net158600, A2 => I(2), A3 => net142483, ZN => 
                           O(2));
   U9 : NAND2_X1 port map( A1 => I(0), A2 => I(1), ZN => net142483);
   U10 : XNOR2_X1 port map( A => I(1), B => I(0), ZN => net158600);
   U11 : XNOR2_X1 port map( A => I(1), B => I(0), ZN => net156612);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_BOOTHMUL_N32.all;

entity BOOTHMUL_N32 is

   port( A, B : in std_logic_vector (31 downto 0);  P : out std_logic_vector 
         (63 downto 0));

end BOOTHMUL_N32;

architecture SYN_STRUCTURAL of BOOTHMUL_N32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component BOOTHMUL_N32_DW01_add_0
      port( A, B : in std_logic_vector (63 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (63 downto 0);  CO : out std_logic);
   end component;
   
   component RCA_generic_N64_1
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_2
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_3
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_4
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_5
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_6
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_7
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_8
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_9
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_10
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_11
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_12
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_13
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_14
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_generic_N64_0
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX51_GENERIC_N64_1
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_2
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_3
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_4
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_5
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_6
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_7
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_8
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_9
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_10
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_11
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_12
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_13
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_14
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_15
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component MUX51_GENERIC_N64_0
      port( A, B, C, D, E : in std_logic_vector (63 downto 0);  SEL : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (63 downto
            0));
   end component;
   
   component BOOTH_ENCODER_5
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_6
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_7
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_8
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_9
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_10
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_11
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_12
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_13
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_14
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_15
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_16
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_17
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_18
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_19
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   component BOOTH_ENCODER_4
      port( I : in std_logic_vector (2 downto 0);  O : out std_logic_vector (2 
            downto 0));
   end component;
   
   signal X_Logic1_port, X_Logic0_port, encoder_out_47_port, 
      encoder_out_46_port, encoder_out_45_port, encoder_out_44_port, 
      encoder_out_43_port, encoder_out_42_port, encoder_out_41_port, 
      encoder_out_40_port, encoder_out_39_port, encoder_out_38_port, 
      encoder_out_37_port, encoder_out_36_port, encoder_out_35_port, 
      encoder_out_34_port, encoder_out_33_port, encoder_out_32_port, 
      encoder_out_31_port, encoder_out_30_port, encoder_out_29_port, 
      encoder_out_28_port, encoder_out_27_port, encoder_out_26_port, 
      encoder_out_25_port, encoder_out_24_port, encoder_out_23_port, 
      encoder_out_22_port, encoder_out_21_port, encoder_out_20_port, 
      encoder_out_19_port, encoder_out_18_port, encoder_out_17_port, 
      encoder_out_16_port, encoder_out_15_port, encoder_out_14_port, 
      encoder_out_13_port, encoder_out_12_port, encoder_out_11_port, 
      encoder_out_10_port, encoder_out_9_port, encoder_out_8_port, 
      encoder_out_7_port, encoder_out_6_port, encoder_out_5_port, 
      encoder_out_4_port, encoder_out_3_port, encoder_out_2_port, 
      encoder_out_1_port, encoder_out_0_port, mode_15_port, mode_14_port, 
      mode_13_port, mode_12_port, mode_11_port, mode_10_port, mode_9_port, 
      mode_8_port, mode_7_port, mode_6_port, mode_5_port, mode_4_port, 
      mode_3_port, mode_2_port, mode_1_port, mux_out_7_63_port, 
      mux_out_7_62_port, mux_out_7_61_port, mux_out_7_60_port, 
      mux_out_7_59_port, mux_out_7_58_port, mux_out_7_57_port, 
      mux_out_7_56_port, mux_out_7_55_port, mux_out_7_54_port, 
      mux_out_7_53_port, mux_out_7_52_port, mux_out_7_51_port, 
      mux_out_7_50_port, mux_out_7_49_port, mux_out_7_48_port, 
      mux_out_7_47_port, mux_out_7_46_port, mux_out_7_45_port, 
      mux_out_7_44_port, mux_out_7_43_port, mux_out_7_42_port, 
      mux_out_7_41_port, mux_out_7_40_port, mux_out_7_39_port, 
      mux_out_7_38_port, mux_out_7_37_port, mux_out_7_36_port, 
      mux_out_7_35_port, mux_out_7_34_port, mux_out_7_33_port, 
      mux_out_7_32_port, mux_out_7_31_port, mux_out_7_30_port, 
      mux_out_7_29_port, mux_out_7_28_port, mux_out_7_27_port, 
      mux_out_7_26_port, mux_out_7_25_port, mux_out_7_24_port, 
      mux_out_7_23_port, mux_out_7_22_port, mux_out_7_21_port, 
      mux_out_7_20_port, mux_out_7_19_port, mux_out_7_18_port, 
      mux_out_7_17_port, mux_out_7_16_port, mux_out_7_15_port, 
      mux_out_7_14_port, mux_out_7_13_port, mux_out_7_12_port, 
      mux_out_7_11_port, mux_out_7_10_port, mux_out_7_9_port, mux_out_7_8_port,
      mux_out_7_7_port, mux_out_7_6_port, mux_out_7_5_port, mux_out_7_4_port, 
      mux_out_7_3_port, mux_out_7_2_port, mux_out_7_1_port, mux_out_7_0_port, 
      mux_out_6_63_port, mux_out_6_62_port, mux_out_6_61_port, 
      mux_out_6_60_port, mux_out_6_59_port, mux_out_6_58_port, 
      mux_out_6_57_port, mux_out_6_56_port, mux_out_6_55_port, 
      mux_out_6_54_port, mux_out_6_53_port, mux_out_6_52_port, 
      mux_out_6_51_port, mux_out_6_50_port, mux_out_6_49_port, 
      mux_out_6_48_port, mux_out_6_47_port, mux_out_6_46_port, 
      mux_out_6_45_port, mux_out_6_44_port, mux_out_6_43_port, 
      mux_out_6_42_port, mux_out_6_41_port, mux_out_6_40_port, 
      mux_out_6_39_port, mux_out_6_38_port, mux_out_6_37_port, 
      mux_out_6_36_port, mux_out_6_35_port, mux_out_6_34_port, 
      mux_out_6_33_port, mux_out_6_32_port, mux_out_6_31_port, 
      mux_out_6_30_port, mux_out_6_29_port, mux_out_6_28_port, 
      mux_out_6_27_port, mux_out_6_26_port, mux_out_6_25_port, 
      mux_out_6_24_port, mux_out_6_23_port, mux_out_6_22_port, 
      mux_out_6_21_port, mux_out_6_20_port, mux_out_6_19_port, 
      mux_out_6_18_port, mux_out_6_17_port, mux_out_6_16_port, 
      mux_out_6_15_port, mux_out_6_14_port, mux_out_6_13_port, 
      mux_out_6_12_port, mux_out_6_11_port, mux_out_6_10_port, mux_out_6_9_port
      , mux_out_6_8_port, mux_out_6_7_port, mux_out_6_6_port, mux_out_6_5_port,
      mux_out_6_4_port, mux_out_6_3_port, mux_out_6_2_port, mux_out_6_1_port, 
      mux_out_6_0_port, mux_out_5_63_port, mux_out_5_62_port, mux_out_5_61_port
      , mux_out_5_60_port, mux_out_5_59_port, mux_out_5_58_port, 
      mux_out_5_57_port, mux_out_5_56_port, mux_out_5_55_port, 
      mux_out_5_54_port, mux_out_5_53_port, mux_out_5_52_port, 
      mux_out_5_51_port, mux_out_5_50_port, mux_out_5_49_port, 
      mux_out_5_48_port, mux_out_5_47_port, mux_out_5_46_port, 
      mux_out_5_45_port, mux_out_5_44_port, mux_out_5_43_port, 
      mux_out_5_42_port, mux_out_5_41_port, mux_out_5_40_port, 
      mux_out_5_39_port, mux_out_5_38_port, mux_out_5_37_port, 
      mux_out_5_36_port, mux_out_5_35_port, mux_out_5_34_port, 
      mux_out_5_33_port, mux_out_5_32_port, mux_out_5_31_port, 
      mux_out_5_30_port, mux_out_5_29_port, mux_out_5_28_port, 
      mux_out_5_27_port, mux_out_5_26_port, mux_out_5_25_port, 
      mux_out_5_24_port, mux_out_5_23_port, mux_out_5_22_port, 
      mux_out_5_21_port, mux_out_5_20_port, mux_out_5_19_port, 
      mux_out_5_18_port, mux_out_5_17_port, mux_out_5_16_port, 
      mux_out_5_15_port, mux_out_5_14_port, mux_out_5_13_port, 
      mux_out_5_12_port, mux_out_5_11_port, mux_out_5_10_port, mux_out_5_9_port
      , mux_out_5_8_port, mux_out_5_7_port, mux_out_5_6_port, mux_out_5_5_port,
      mux_out_5_4_port, mux_out_5_3_port, mux_out_5_2_port, mux_out_5_1_port, 
      mux_out_5_0_port, mux_out_4_63_port, mux_out_4_62_port, mux_out_4_61_port
      , mux_out_4_60_port, mux_out_4_59_port, mux_out_4_58_port, 
      mux_out_4_57_port, mux_out_4_56_port, mux_out_4_55_port, 
      mux_out_4_54_port, mux_out_4_53_port, mux_out_4_52_port, 
      mux_out_4_51_port, mux_out_4_50_port, mux_out_4_49_port, 
      mux_out_4_48_port, mux_out_4_47_port, mux_out_4_46_port, 
      mux_out_4_45_port, mux_out_4_44_port, mux_out_4_43_port, 
      mux_out_4_42_port, mux_out_4_41_port, mux_out_4_40_port, 
      mux_out_4_39_port, mux_out_4_38_port, mux_out_4_37_port, 
      mux_out_4_36_port, mux_out_4_35_port, mux_out_4_34_port, 
      mux_out_4_33_port, mux_out_4_32_port, mux_out_4_31_port, 
      mux_out_4_30_port, mux_out_4_29_port, mux_out_4_28_port, 
      mux_out_4_27_port, mux_out_4_26_port, mux_out_4_25_port, 
      mux_out_4_24_port, mux_out_4_23_port, mux_out_4_22_port, 
      mux_out_4_21_port, mux_out_4_20_port, mux_out_4_19_port, 
      mux_out_4_18_port, mux_out_4_17_port, mux_out_4_16_port, 
      mux_out_4_15_port, mux_out_4_14_port, mux_out_4_13_port, 
      mux_out_4_12_port, mux_out_4_11_port, mux_out_4_10_port, mux_out_4_9_port
      , mux_out_4_8_port, mux_out_4_7_port, mux_out_4_6_port, mux_out_4_5_port,
      mux_out_4_4_port, mux_out_4_3_port, mux_out_4_2_port, mux_out_4_1_port, 
      mux_out_4_0_port, mux_out_3_63_port, mux_out_3_62_port, mux_out_3_61_port
      , mux_out_3_60_port, mux_out_3_59_port, mux_out_3_58_port, 
      mux_out_3_57_port, mux_out_3_56_port, mux_out_3_55_port, 
      mux_out_3_54_port, mux_out_3_53_port, mux_out_3_52_port, 
      mux_out_3_51_port, mux_out_3_50_port, mux_out_3_49_port, 
      mux_out_3_48_port, mux_out_3_47_port, mux_out_3_46_port, 
      mux_out_3_45_port, mux_out_3_44_port, mux_out_3_43_port, 
      mux_out_3_42_port, mux_out_3_41_port, mux_out_3_40_port, 
      mux_out_3_39_port, mux_out_3_38_port, mux_out_3_37_port, 
      mux_out_3_36_port, mux_out_3_35_port, mux_out_3_34_port, 
      mux_out_3_33_port, mux_out_3_32_port, mux_out_3_31_port, 
      mux_out_3_30_port, mux_out_3_29_port, mux_out_3_28_port, 
      mux_out_3_27_port, mux_out_3_26_port, mux_out_3_25_port, 
      mux_out_3_24_port, mux_out_3_23_port, mux_out_3_22_port, 
      mux_out_3_21_port, mux_out_3_20_port, mux_out_3_19_port, 
      mux_out_3_18_port, mux_out_3_17_port, mux_out_3_16_port, 
      mux_out_3_15_port, mux_out_3_14_port, mux_out_3_13_port, 
      mux_out_3_12_port, mux_out_3_11_port, mux_out_3_10_port, mux_out_3_9_port
      , mux_out_3_8_port, mux_out_3_7_port, mux_out_3_6_port, mux_out_3_5_port,
      mux_out_3_4_port, mux_out_3_3_port, mux_out_3_2_port, mux_out_3_1_port, 
      mux_out_3_0_port, mux_out_2_63_port, mux_out_2_62_port, mux_out_2_61_port
      , mux_out_2_60_port, mux_out_2_59_port, mux_out_2_58_port, 
      mux_out_2_57_port, mux_out_2_56_port, mux_out_2_55_port, 
      mux_out_2_54_port, mux_out_2_53_port, mux_out_2_52_port, 
      mux_out_2_51_port, mux_out_2_50_port, mux_out_2_49_port, 
      mux_out_2_48_port, mux_out_2_47_port, mux_out_2_46_port, 
      mux_out_2_45_port, mux_out_2_44_port, mux_out_2_43_port, 
      mux_out_2_42_port, mux_out_2_41_port, mux_out_2_40_port, 
      mux_out_2_39_port, mux_out_2_38_port, mux_out_2_37_port, 
      mux_out_2_36_port, mux_out_2_35_port, mux_out_2_34_port, 
      mux_out_2_33_port, mux_out_2_32_port, mux_out_2_31_port, 
      mux_out_2_30_port, mux_out_2_29_port, mux_out_2_28_port, 
      mux_out_2_27_port, mux_out_2_26_port, mux_out_2_25_port, 
      mux_out_2_24_port, mux_out_2_23_port, mux_out_2_22_port, 
      mux_out_2_21_port, mux_out_2_20_port, mux_out_2_19_port, 
      mux_out_2_18_port, mux_out_2_17_port, mux_out_2_16_port, 
      mux_out_2_15_port, mux_out_2_14_port, mux_out_2_13_port, 
      mux_out_2_12_port, mux_out_2_11_port, mux_out_2_10_port, mux_out_2_9_port
      , mux_out_2_8_port, mux_out_2_7_port, mux_out_2_6_port, mux_out_2_5_port,
      mux_out_2_4_port, mux_out_2_3_port, mux_out_2_2_port, mux_out_2_1_port, 
      mux_out_2_0_port, mux_out_1_63_port, mux_out_1_62_port, mux_out_1_61_port
      , mux_out_1_60_port, mux_out_1_59_port, mux_out_1_58_port, 
      mux_out_1_57_port, mux_out_1_56_port, mux_out_1_55_port, 
      mux_out_1_54_port, mux_out_1_53_port, mux_out_1_52_port, 
      mux_out_1_51_port, mux_out_1_50_port, mux_out_1_49_port, 
      mux_out_1_48_port, mux_out_1_47_port, mux_out_1_46_port, 
      mux_out_1_45_port, mux_out_1_44_port, mux_out_1_43_port, 
      mux_out_1_42_port, mux_out_1_41_port, mux_out_1_40_port, 
      mux_out_1_39_port, mux_out_1_38_port, mux_out_1_37_port, 
      mux_out_1_36_port, mux_out_1_35_port, mux_out_1_34_port, 
      mux_out_1_33_port, mux_out_1_32_port, mux_out_1_31_port, 
      mux_out_1_30_port, mux_out_1_29_port, mux_out_1_28_port, 
      mux_out_1_27_port, mux_out_1_26_port, mux_out_1_25_port, 
      mux_out_1_24_port, mux_out_1_23_port, mux_out_1_22_port, 
      mux_out_1_21_port, mux_out_1_20_port, mux_out_1_19_port, 
      mux_out_1_18_port, mux_out_1_17_port, mux_out_1_16_port, 
      mux_out_1_15_port, mux_out_1_14_port, mux_out_1_13_port, 
      mux_out_1_12_port, mux_out_1_11_port, mux_out_1_10_port, mux_out_1_9_port
      , mux_out_1_8_port, mux_out_1_7_port, mux_out_1_6_port, mux_out_1_5_port,
      mux_out_1_4_port, mux_out_1_3_port, mux_out_1_2_port, mux_out_1_1_port, 
      mux_out_1_0_port, mux_out_15_63_port, mux_out_15_62_port, 
      mux_out_15_61_port, mux_out_15_60_port, mux_out_15_59_port, 
      mux_out_15_58_port, mux_out_15_57_port, mux_out_15_56_port, 
      mux_out_15_55_port, mux_out_15_54_port, mux_out_15_53_port, 
      mux_out_15_52_port, mux_out_15_51_port, mux_out_15_50_port, 
      mux_out_15_49_port, mux_out_15_48_port, mux_out_15_47_port, 
      mux_out_15_46_port, mux_out_15_45_port, mux_out_15_44_port, 
      mux_out_15_43_port, mux_out_15_42_port, mux_out_15_41_port, 
      mux_out_15_40_port, mux_out_15_39_port, mux_out_15_38_port, 
      mux_out_15_37_port, mux_out_15_36_port, mux_out_15_35_port, 
      mux_out_15_34_port, mux_out_15_33_port, mux_out_15_32_port, 
      mux_out_15_31_port, mux_out_15_30_port, mux_out_15_29_port, 
      mux_out_15_28_port, mux_out_15_27_port, mux_out_15_26_port, 
      mux_out_15_25_port, mux_out_15_24_port, mux_out_15_23_port, 
      mux_out_15_22_port, mux_out_15_21_port, mux_out_15_20_port, 
      mux_out_15_19_port, mux_out_15_18_port, mux_out_15_17_port, 
      mux_out_15_16_port, mux_out_15_15_port, mux_out_15_14_port, 
      mux_out_15_13_port, mux_out_15_12_port, mux_out_15_11_port, 
      mux_out_15_10_port, mux_out_15_9_port, mux_out_15_8_port, 
      mux_out_15_7_port, mux_out_15_6_port, mux_out_15_5_port, 
      mux_out_15_4_port, mux_out_15_3_port, mux_out_15_2_port, 
      mux_out_15_1_port, mux_out_15_0_port, mux_out_14_63_port, 
      mux_out_14_62_port, mux_out_14_61_port, mux_out_14_60_port, 
      mux_out_14_59_port, mux_out_14_58_port, mux_out_14_57_port, 
      mux_out_14_56_port, mux_out_14_55_port, mux_out_14_54_port, 
      mux_out_14_53_port, mux_out_14_52_port, mux_out_14_51_port, 
      mux_out_14_50_port, mux_out_14_49_port, mux_out_14_48_port, 
      mux_out_14_47_port, mux_out_14_46_port, mux_out_14_45_port, 
      mux_out_14_44_port, mux_out_14_43_port, mux_out_14_42_port, 
      mux_out_14_41_port, mux_out_14_40_port, mux_out_14_39_port, 
      mux_out_14_38_port, mux_out_14_37_port, mux_out_14_36_port, 
      mux_out_14_35_port, mux_out_14_34_port, mux_out_14_33_port, 
      mux_out_14_32_port, mux_out_14_31_port, mux_out_14_30_port, 
      mux_out_14_29_port, mux_out_14_28_port, mux_out_14_27_port, 
      mux_out_14_26_port, mux_out_14_25_port, mux_out_14_24_port, 
      mux_out_14_23_port, mux_out_14_22_port, mux_out_14_21_port, 
      mux_out_14_20_port, mux_out_14_19_port, mux_out_14_18_port, 
      mux_out_14_17_port, mux_out_14_16_port, mux_out_14_15_port, 
      mux_out_14_14_port, mux_out_14_13_port, mux_out_14_12_port, 
      mux_out_14_11_port, mux_out_14_10_port, mux_out_14_9_port, 
      mux_out_14_8_port, mux_out_14_7_port, mux_out_14_6_port, 
      mux_out_14_5_port, mux_out_14_4_port, mux_out_14_3_port, 
      mux_out_14_2_port, mux_out_14_1_port, mux_out_14_0_port, 
      mux_out_13_63_port, mux_out_13_62_port, mux_out_13_61_port, 
      mux_out_13_60_port, mux_out_13_59_port, mux_out_13_58_port, 
      mux_out_13_57_port, mux_out_13_56_port, mux_out_13_55_port, 
      mux_out_13_54_port, mux_out_13_53_port, mux_out_13_52_port, 
      mux_out_13_51_port, mux_out_13_50_port, mux_out_13_49_port, 
      mux_out_13_48_port, mux_out_13_47_port, mux_out_13_46_port, 
      mux_out_13_45_port, mux_out_13_44_port, mux_out_13_43_port, 
      mux_out_13_42_port, mux_out_13_41_port, mux_out_13_40_port, 
      mux_out_13_39_port, mux_out_13_38_port, mux_out_13_37_port, 
      mux_out_13_36_port, mux_out_13_35_port, mux_out_13_34_port, 
      mux_out_13_33_port, mux_out_13_32_port, mux_out_13_31_port, 
      mux_out_13_30_port, mux_out_13_29_port, mux_out_13_28_port, 
      mux_out_13_27_port, mux_out_13_26_port, mux_out_13_25_port, 
      mux_out_13_24_port, mux_out_13_23_port, mux_out_13_22_port, 
      mux_out_13_21_port, mux_out_13_20_port, mux_out_13_19_port, 
      mux_out_13_18_port, mux_out_13_17_port, mux_out_13_16_port, 
      mux_out_13_15_port, mux_out_13_14_port, mux_out_13_13_port, 
      mux_out_13_12_port, mux_out_13_11_port, mux_out_13_10_port, 
      mux_out_13_9_port, mux_out_13_8_port, mux_out_13_7_port, 
      mux_out_13_6_port, mux_out_13_5_port, mux_out_13_4_port, 
      mux_out_13_3_port, mux_out_13_2_port, mux_out_13_1_port, 
      mux_out_13_0_port, mux_out_12_63_port, mux_out_12_62_port, 
      mux_out_12_61_port, mux_out_12_60_port, mux_out_12_59_port, 
      mux_out_12_58_port, mux_out_12_57_port, mux_out_12_56_port, 
      mux_out_12_55_port, mux_out_12_54_port, mux_out_12_53_port, 
      mux_out_12_52_port, mux_out_12_51_port, mux_out_12_50_port, 
      mux_out_12_49_port, mux_out_12_48_port, mux_out_12_47_port, 
      mux_out_12_46_port, mux_out_12_45_port, mux_out_12_44_port, 
      mux_out_12_43_port, mux_out_12_42_port, mux_out_12_41_port, 
      mux_out_12_40_port, mux_out_12_39_port, mux_out_12_38_port, 
      mux_out_12_37_port, mux_out_12_36_port, mux_out_12_35_port, 
      mux_out_12_34_port, mux_out_12_33_port, mux_out_12_32_port, 
      mux_out_12_31_port, mux_out_12_30_port, mux_out_12_29_port, 
      mux_out_12_28_port, mux_out_12_27_port, mux_out_12_26_port, 
      mux_out_12_25_port, mux_out_12_24_port, mux_out_12_23_port, 
      mux_out_12_22_port, mux_out_12_21_port, mux_out_12_20_port, 
      mux_out_12_19_port, mux_out_12_18_port, mux_out_12_17_port, 
      mux_out_12_16_port, mux_out_12_15_port, mux_out_12_14_port, 
      mux_out_12_13_port, mux_out_12_12_port, mux_out_12_11_port, 
      mux_out_12_10_port, mux_out_12_9_port, mux_out_12_8_port, 
      mux_out_12_7_port, mux_out_12_6_port, mux_out_12_5_port, 
      mux_out_12_4_port, mux_out_12_3_port, mux_out_12_2_port, 
      mux_out_12_1_port, mux_out_12_0_port, mux_out_11_63_port, 
      mux_out_11_62_port, mux_out_11_61_port, mux_out_11_60_port, 
      mux_out_11_59_port, mux_out_11_58_port, mux_out_11_57_port, 
      mux_out_11_56_port, mux_out_11_55_port, mux_out_11_54_port, 
      mux_out_11_53_port, mux_out_11_52_port, mux_out_11_51_port, 
      mux_out_11_50_port, mux_out_11_49_port, mux_out_11_48_port, 
      mux_out_11_47_port, mux_out_11_46_port, mux_out_11_45_port, 
      mux_out_11_44_port, mux_out_11_43_port, mux_out_11_42_port, 
      mux_out_11_41_port, mux_out_11_40_port, mux_out_11_39_port, 
      mux_out_11_38_port, mux_out_11_37_port, mux_out_11_36_port, 
      mux_out_11_35_port, mux_out_11_34_port, mux_out_11_33_port, 
      mux_out_11_32_port, mux_out_11_31_port, mux_out_11_30_port, 
      mux_out_11_29_port, mux_out_11_28_port, mux_out_11_27_port, 
      mux_out_11_26_port, mux_out_11_25_port, mux_out_11_24_port, 
      mux_out_11_23_port, mux_out_11_22_port, mux_out_11_21_port, 
      mux_out_11_20_port, mux_out_11_19_port, mux_out_11_18_port, 
      mux_out_11_17_port, mux_out_11_16_port, mux_out_11_15_port, 
      mux_out_11_14_port, mux_out_11_13_port, mux_out_11_12_port, 
      mux_out_11_11_port, mux_out_11_10_port, mux_out_11_9_port, 
      mux_out_11_8_port, mux_out_11_7_port, mux_out_11_6_port, 
      mux_out_11_5_port, mux_out_11_4_port, mux_out_11_3_port, 
      mux_out_11_2_port, mux_out_11_1_port, mux_out_11_0_port, 
      mux_out_10_63_port, mux_out_10_62_port, mux_out_10_61_port, 
      mux_out_10_60_port, mux_out_10_59_port, mux_out_10_58_port, 
      mux_out_10_57_port, mux_out_10_56_port, mux_out_10_55_port, 
      mux_out_10_54_port, mux_out_10_53_port, mux_out_10_52_port, 
      mux_out_10_51_port, mux_out_10_50_port, mux_out_10_49_port, 
      mux_out_10_48_port, mux_out_10_47_port, mux_out_10_46_port, 
      mux_out_10_45_port, mux_out_10_44_port, mux_out_10_43_port, 
      mux_out_10_42_port, mux_out_10_41_port, mux_out_10_40_port, 
      mux_out_10_39_port, mux_out_10_38_port, mux_out_10_37_port, 
      mux_out_10_36_port, mux_out_10_35_port, mux_out_10_34_port, 
      mux_out_10_33_port, mux_out_10_32_port, mux_out_10_31_port, 
      mux_out_10_30_port, mux_out_10_29_port, mux_out_10_28_port, 
      mux_out_10_27_port, mux_out_10_26_port, mux_out_10_25_port, 
      mux_out_10_24_port, mux_out_10_23_port, mux_out_10_22_port, 
      mux_out_10_21_port, mux_out_10_20_port, mux_out_10_19_port, 
      mux_out_10_18_port, mux_out_10_17_port, mux_out_10_16_port, 
      mux_out_10_15_port, mux_out_10_14_port, mux_out_10_13_port, 
      mux_out_10_12_port, mux_out_10_11_port, mux_out_10_10_port, 
      mux_out_10_9_port, mux_out_10_8_port, mux_out_10_7_port, 
      mux_out_10_6_port, mux_out_10_5_port, mux_out_10_4_port, 
      mux_out_10_3_port, mux_out_10_2_port, mux_out_10_1_port, 
      mux_out_10_0_port, mux_out_9_63_port, mux_out_9_62_port, 
      mux_out_9_61_port, mux_out_9_60_port, mux_out_9_59_port, 
      mux_out_9_58_port, mux_out_9_57_port, mux_out_9_56_port, 
      mux_out_9_55_port, mux_out_9_54_port, mux_out_9_53_port, 
      mux_out_9_52_port, mux_out_9_51_port, mux_out_9_50_port, 
      mux_out_9_49_port, mux_out_9_48_port, mux_out_9_47_port, 
      mux_out_9_46_port, mux_out_9_45_port, mux_out_9_44_port, 
      mux_out_9_43_port, mux_out_9_42_port, mux_out_9_41_port, 
      mux_out_9_40_port, mux_out_9_39_port, mux_out_9_38_port, 
      mux_out_9_37_port, mux_out_9_36_port, mux_out_9_35_port, 
      mux_out_9_34_port, mux_out_9_33_port, mux_out_9_32_port, 
      mux_out_9_31_port, mux_out_9_30_port, mux_out_9_29_port, 
      mux_out_9_28_port, mux_out_9_27_port, mux_out_9_26_port, 
      mux_out_9_25_port, mux_out_9_24_port, mux_out_9_23_port, 
      mux_out_9_22_port, mux_out_9_21_port, mux_out_9_20_port, 
      mux_out_9_19_port, mux_out_9_18_port, mux_out_9_17_port, 
      mux_out_9_16_port, mux_out_9_15_port, mux_out_9_14_port, 
      mux_out_9_13_port, mux_out_9_12_port, mux_out_9_11_port, 
      mux_out_9_10_port, mux_out_9_9_port, mux_out_9_8_port, mux_out_9_7_port, 
      mux_out_9_6_port, mux_out_9_5_port, mux_out_9_4_port, mux_out_9_3_port, 
      mux_out_9_2_port, mux_out_9_1_port, mux_out_9_0_port, mux_out_8_63_port, 
      mux_out_8_62_port, mux_out_8_61_port, mux_out_8_60_port, 
      mux_out_8_59_port, mux_out_8_58_port, mux_out_8_57_port, 
      mux_out_8_56_port, mux_out_8_55_port, mux_out_8_54_port, 
      mux_out_8_53_port, mux_out_8_52_port, mux_out_8_51_port, 
      mux_out_8_50_port, mux_out_8_49_port, mux_out_8_48_port, 
      mux_out_8_47_port, mux_out_8_46_port, mux_out_8_45_port, 
      mux_out_8_44_port, mux_out_8_43_port, mux_out_8_42_port, 
      mux_out_8_41_port, mux_out_8_40_port, mux_out_8_39_port, 
      mux_out_8_38_port, mux_out_8_37_port, mux_out_8_36_port, 
      mux_out_8_35_port, mux_out_8_34_port, mux_out_8_33_port, 
      mux_out_8_32_port, mux_out_8_31_port, mux_out_8_30_port, 
      mux_out_8_29_port, mux_out_8_28_port, mux_out_8_27_port, 
      mux_out_8_26_port, mux_out_8_25_port, mux_out_8_24_port, 
      mux_out_8_23_port, mux_out_8_22_port, mux_out_8_21_port, 
      mux_out_8_20_port, mux_out_8_19_port, mux_out_8_18_port, 
      mux_out_8_17_port, mux_out_8_16_port, mux_out_8_15_port, 
      mux_out_8_14_port, mux_out_8_13_port, mux_out_8_12_port, 
      mux_out_8_11_port, mux_out_8_10_port, mux_out_8_9_port, mux_out_8_8_port,
      mux_out_8_7_port, mux_out_8_6_port, mux_out_8_5_port, mux_out_8_4_port, 
      mux_out_8_3_port, mux_out_8_2_port, mux_out_8_1_port, mux_out_8_0_port, 
      add_in_7_63_port, add_in_7_62_port, add_in_7_61_port, add_in_7_60_port, 
      add_in_7_59_port, add_in_7_58_port, add_in_7_57_port, add_in_7_56_port, 
      add_in_7_55_port, add_in_7_54_port, add_in_7_53_port, add_in_7_52_port, 
      add_in_7_51_port, add_in_7_50_port, add_in_7_49_port, add_in_7_48_port, 
      add_in_7_47_port, add_in_7_46_port, add_in_7_45_port, add_in_7_44_port, 
      add_in_7_43_port, add_in_7_42_port, add_in_7_41_port, add_in_7_40_port, 
      add_in_7_39_port, add_in_7_38_port, add_in_7_37_port, add_in_7_36_port, 
      add_in_7_35_port, add_in_7_34_port, add_in_7_33_port, add_in_7_32_port, 
      add_in_7_31_port, add_in_7_30_port, add_in_7_29_port, add_in_7_28_port, 
      add_in_7_27_port, add_in_7_26_port, add_in_7_25_port, add_in_7_24_port, 
      add_in_7_23_port, add_in_7_22_port, add_in_7_21_port, add_in_7_20_port, 
      add_in_7_19_port, add_in_7_18_port, add_in_7_17_port, add_in_7_16_port, 
      add_in_7_15_port, add_in_7_14_port, add_in_7_13_port, add_in_7_12_port, 
      add_in_7_11_port, add_in_7_10_port, add_in_7_9_port, add_in_7_8_port, 
      add_in_7_7_port, add_in_7_6_port, add_in_7_5_port, add_in_7_4_port, 
      add_in_7_3_port, add_in_7_2_port, add_in_7_1_port, add_in_7_0_port, 
      add_in_6_63_port, add_in_6_62_port, add_in_6_61_port, add_in_6_60_port, 
      add_in_6_59_port, add_in_6_58_port, add_in_6_57_port, add_in_6_56_port, 
      add_in_6_55_port, add_in_6_54_port, add_in_6_53_port, add_in_6_52_port, 
      add_in_6_51_port, add_in_6_50_port, add_in_6_49_port, add_in_6_48_port, 
      add_in_6_47_port, add_in_6_46_port, add_in_6_45_port, add_in_6_44_port, 
      add_in_6_43_port, add_in_6_42_port, add_in_6_41_port, add_in_6_40_port, 
      add_in_6_39_port, add_in_6_38_port, add_in_6_37_port, add_in_6_36_port, 
      add_in_6_35_port, add_in_6_34_port, add_in_6_33_port, add_in_6_32_port, 
      add_in_6_31_port, add_in_6_30_port, add_in_6_29_port, add_in_6_28_port, 
      add_in_6_27_port, add_in_6_26_port, add_in_6_25_port, add_in_6_24_port, 
      add_in_6_23_port, add_in_6_22_port, add_in_6_21_port, add_in_6_20_port, 
      add_in_6_19_port, add_in_6_18_port, add_in_6_17_port, add_in_6_16_port, 
      add_in_6_15_port, add_in_6_14_port, add_in_6_13_port, add_in_6_12_port, 
      add_in_6_11_port, add_in_6_10_port, add_in_6_9_port, add_in_6_8_port, 
      add_in_6_7_port, add_in_6_6_port, add_in_6_5_port, add_in_6_4_port, 
      add_in_6_3_port, add_in_6_2_port, add_in_6_1_port, add_in_6_0_port, 
      add_in_5_63_port, add_in_5_62_port, add_in_5_61_port, add_in_5_60_port, 
      add_in_5_59_port, add_in_5_58_port, add_in_5_57_port, add_in_5_56_port, 
      add_in_5_55_port, add_in_5_54_port, add_in_5_53_port, add_in_5_52_port, 
      add_in_5_51_port, add_in_5_50_port, add_in_5_49_port, add_in_5_48_port, 
      add_in_5_47_port, add_in_5_46_port, add_in_5_45_port, add_in_5_44_port, 
      add_in_5_43_port, add_in_5_42_port, add_in_5_41_port, add_in_5_40_port, 
      add_in_5_39_port, add_in_5_38_port, add_in_5_37_port, add_in_5_36_port, 
      add_in_5_35_port, add_in_5_34_port, add_in_5_33_port, add_in_5_32_port, 
      add_in_5_31_port, add_in_5_30_port, add_in_5_29_port, add_in_5_28_port, 
      add_in_5_27_port, add_in_5_26_port, add_in_5_25_port, add_in_5_24_port, 
      add_in_5_23_port, add_in_5_22_port, add_in_5_21_port, add_in_5_20_port, 
      add_in_5_19_port, add_in_5_18_port, add_in_5_17_port, add_in_5_16_port, 
      add_in_5_15_port, add_in_5_14_port, add_in_5_13_port, add_in_5_12_port, 
      add_in_5_11_port, add_in_5_10_port, add_in_5_9_port, add_in_5_8_port, 
      add_in_5_7_port, add_in_5_6_port, add_in_5_5_port, add_in_5_4_port, 
      add_in_5_3_port, add_in_5_2_port, add_in_5_1_port, add_in_5_0_port, 
      add_in_4_63_port, add_in_4_62_port, add_in_4_61_port, add_in_4_60_port, 
      add_in_4_59_port, add_in_4_58_port, add_in_4_57_port, add_in_4_56_port, 
      add_in_4_55_port, add_in_4_54_port, add_in_4_53_port, add_in_4_52_port, 
      add_in_4_51_port, add_in_4_50_port, add_in_4_49_port, add_in_4_48_port, 
      add_in_4_47_port, add_in_4_46_port, add_in_4_45_port, add_in_4_44_port, 
      add_in_4_43_port, add_in_4_42_port, add_in_4_41_port, add_in_4_40_port, 
      add_in_4_39_port, add_in_4_38_port, add_in_4_37_port, add_in_4_36_port, 
      add_in_4_35_port, add_in_4_34_port, add_in_4_33_port, add_in_4_32_port, 
      add_in_4_31_port, add_in_4_30_port, add_in_4_29_port, add_in_4_28_port, 
      add_in_4_27_port, add_in_4_26_port, add_in_4_25_port, add_in_4_24_port, 
      add_in_4_23_port, add_in_4_22_port, add_in_4_21_port, add_in_4_20_port, 
      add_in_4_19_port, add_in_4_18_port, add_in_4_17_port, add_in_4_16_port, 
      add_in_4_15_port, add_in_4_14_port, add_in_4_13_port, add_in_4_12_port, 
      add_in_4_11_port, add_in_4_10_port, add_in_4_9_port, add_in_4_8_port, 
      add_in_4_7_port, add_in_4_6_port, add_in_4_5_port, add_in_4_4_port, 
      add_in_4_3_port, add_in_4_2_port, add_in_4_1_port, add_in_4_0_port, 
      add_in_3_63_port, add_in_3_62_port, add_in_3_61_port, add_in_3_60_port, 
      add_in_3_59_port, add_in_3_58_port, add_in_3_57_port, add_in_3_56_port, 
      add_in_3_55_port, add_in_3_54_port, add_in_3_53_port, add_in_3_52_port, 
      add_in_3_51_port, add_in_3_50_port, add_in_3_49_port, add_in_3_48_port, 
      add_in_3_47_port, add_in_3_46_port, add_in_3_45_port, add_in_3_44_port, 
      add_in_3_43_port, add_in_3_42_port, add_in_3_41_port, add_in_3_40_port, 
      add_in_3_39_port, add_in_3_38_port, add_in_3_37_port, add_in_3_36_port, 
      add_in_3_35_port, add_in_3_34_port, add_in_3_33_port, add_in_3_32_port, 
      add_in_3_31_port, add_in_3_30_port, add_in_3_29_port, add_in_3_28_port, 
      add_in_3_27_port, add_in_3_26_port, add_in_3_25_port, add_in_3_24_port, 
      add_in_3_23_port, add_in_3_22_port, add_in_3_21_port, add_in_3_20_port, 
      add_in_3_19_port, add_in_3_18_port, add_in_3_17_port, add_in_3_16_port, 
      add_in_3_15_port, add_in_3_14_port, add_in_3_13_port, add_in_3_12_port, 
      add_in_3_11_port, add_in_3_10_port, add_in_3_9_port, add_in_3_8_port, 
      add_in_3_7_port, add_in_3_6_port, add_in_3_5_port, add_in_3_4_port, 
      add_in_3_3_port, add_in_3_2_port, add_in_3_1_port, add_in_3_0_port, 
      add_in_2_63_port, add_in_2_62_port, add_in_2_61_port, add_in_2_60_port, 
      add_in_2_59_port, add_in_2_58_port, add_in_2_57_port, add_in_2_56_port, 
      add_in_2_55_port, add_in_2_54_port, add_in_2_53_port, add_in_2_52_port, 
      add_in_2_51_port, add_in_2_50_port, add_in_2_49_port, add_in_2_48_port, 
      add_in_2_47_port, add_in_2_46_port, add_in_2_45_port, add_in_2_44_port, 
      add_in_2_43_port, add_in_2_42_port, add_in_2_41_port, add_in_2_40_port, 
      add_in_2_39_port, add_in_2_38_port, add_in_2_37_port, add_in_2_36_port, 
      add_in_2_35_port, add_in_2_34_port, add_in_2_33_port, add_in_2_32_port, 
      add_in_2_31_port, add_in_2_30_port, add_in_2_29_port, add_in_2_28_port, 
      add_in_2_27_port, add_in_2_26_port, add_in_2_25_port, add_in_2_24_port, 
      add_in_2_23_port, add_in_2_22_port, add_in_2_21_port, add_in_2_20_port, 
      add_in_2_19_port, add_in_2_18_port, add_in_2_17_port, add_in_2_16_port, 
      add_in_2_15_port, add_in_2_14_port, add_in_2_13_port, add_in_2_12_port, 
      add_in_2_11_port, add_in_2_10_port, add_in_2_9_port, add_in_2_8_port, 
      add_in_2_7_port, add_in_2_6_port, add_in_2_5_port, add_in_2_4_port, 
      add_in_2_3_port, add_in_2_2_port, add_in_2_1_port, add_in_2_0_port, 
      add_in_1_63_port, add_in_1_62_port, add_in_1_61_port, add_in_1_60_port, 
      add_in_1_59_port, add_in_1_58_port, add_in_1_57_port, add_in_1_56_port, 
      add_in_1_55_port, add_in_1_54_port, add_in_1_53_port, add_in_1_52_port, 
      add_in_1_51_port, add_in_1_50_port, add_in_1_49_port, add_in_1_48_port, 
      add_in_1_47_port, add_in_1_46_port, add_in_1_45_port, add_in_1_44_port, 
      add_in_1_43_port, add_in_1_42_port, add_in_1_41_port, add_in_1_40_port, 
      add_in_1_39_port, add_in_1_38_port, add_in_1_37_port, add_in_1_36_port, 
      add_in_1_35_port, add_in_1_34_port, add_in_1_33_port, add_in_1_32_port, 
      add_in_1_31_port, add_in_1_30_port, add_in_1_29_port, add_in_1_28_port, 
      add_in_1_27_port, add_in_1_26_port, add_in_1_25_port, add_in_1_24_port, 
      add_in_1_23_port, add_in_1_22_port, add_in_1_21_port, add_in_1_20_port, 
      add_in_1_19_port, add_in_1_18_port, add_in_1_17_port, add_in_1_16_port, 
      add_in_1_15_port, add_in_1_14_port, add_in_1_13_port, add_in_1_12_port, 
      add_in_1_11_port, add_in_1_10_port, add_in_1_9_port, add_in_1_8_port, 
      add_in_1_7_port, add_in_1_6_port, add_in_1_5_port, add_in_1_4_port, 
      add_in_1_3_port, add_in_1_2_port, add_in_1_1_port, add_in_1_0_port, 
      add_in_0_63_port, add_in_0_62_port, add_in_0_61_port, add_in_0_60_port, 
      add_in_0_59_port, add_in_0_58_port, add_in_0_57_port, add_in_0_56_port, 
      add_in_0_55_port, add_in_0_54_port, add_in_0_53_port, add_in_0_52_port, 
      add_in_0_51_port, add_in_0_50_port, add_in_0_49_port, add_in_0_48_port, 
      add_in_0_47_port, add_in_0_46_port, add_in_0_45_port, add_in_0_44_port, 
      add_in_0_43_port, add_in_0_42_port, add_in_0_41_port, add_in_0_40_port, 
      add_in_0_39_port, add_in_0_38_port, add_in_0_37_port, add_in_0_36_port, 
      add_in_0_35_port, add_in_0_34_port, add_in_0_33_port, add_in_0_32_port, 
      add_in_0_31_port, add_in_0_30_port, add_in_0_29_port, add_in_0_28_port, 
      add_in_0_27_port, add_in_0_26_port, add_in_0_25_port, add_in_0_24_port, 
      add_in_0_23_port, add_in_0_22_port, add_in_0_21_port, add_in_0_20_port, 
      add_in_0_19_port, add_in_0_18_port, add_in_0_17_port, add_in_0_16_port, 
      add_in_0_15_port, add_in_0_14_port, add_in_0_13_port, add_in_0_12_port, 
      add_in_0_11_port, add_in_0_10_port, add_in_0_9_port, add_in_0_8_port, 
      add_in_0_7_port, add_in_0_6_port, add_in_0_5_port, add_in_0_4_port, 
      add_in_0_3_port, add_in_0_2_port, add_in_0_1_port, add_in_0_0_port, 
      add_in_15_63_port, add_in_15_62_port, add_in_15_61_port, 
      add_in_15_60_port, add_in_15_59_port, add_in_15_58_port, 
      add_in_15_57_port, add_in_15_56_port, add_in_15_55_port, 
      add_in_15_54_port, add_in_15_53_port, add_in_15_52_port, 
      add_in_15_51_port, add_in_15_50_port, add_in_15_49_port, 
      add_in_15_48_port, add_in_15_47_port, add_in_15_46_port, 
      add_in_15_45_port, add_in_15_44_port, add_in_15_43_port, 
      add_in_15_42_port, add_in_15_41_port, add_in_15_40_port, 
      add_in_15_39_port, add_in_15_38_port, add_in_15_37_port, 
      add_in_15_36_port, add_in_15_35_port, add_in_15_34_port, 
      add_in_15_33_port, add_in_15_32_port, add_in_15_31_port, 
      add_in_15_30_port, add_in_15_29_port, add_in_15_28_port, 
      add_in_15_27_port, add_in_15_26_port, add_in_15_25_port, 
      add_in_15_24_port, add_in_15_23_port, add_in_15_22_port, 
      add_in_15_21_port, add_in_15_20_port, add_in_15_19_port, 
      add_in_15_18_port, add_in_15_17_port, add_in_15_16_port, 
      add_in_15_15_port, add_in_15_14_port, add_in_15_13_port, 
      add_in_15_12_port, add_in_15_11_port, add_in_15_10_port, add_in_15_9_port
      , add_in_15_8_port, add_in_15_7_port, add_in_15_6_port, add_in_15_5_port,
      add_in_15_4_port, add_in_15_3_port, add_in_15_2_port, add_in_15_1_port, 
      add_in_15_0_port, add_in_14_63_port, add_in_14_62_port, add_in_14_61_port
      , add_in_14_60_port, add_in_14_59_port, add_in_14_58_port, 
      add_in_14_57_port, add_in_14_56_port, add_in_14_55_port, 
      add_in_14_54_port, add_in_14_53_port, add_in_14_52_port, 
      add_in_14_51_port, add_in_14_50_port, add_in_14_49_port, 
      add_in_14_48_port, add_in_14_47_port, add_in_14_46_port, 
      add_in_14_45_port, add_in_14_44_port, add_in_14_43_port, 
      add_in_14_42_port, add_in_14_41_port, add_in_14_40_port, 
      add_in_14_39_port, add_in_14_38_port, add_in_14_37_port, 
      add_in_14_36_port, add_in_14_35_port, add_in_14_34_port, 
      add_in_14_33_port, add_in_14_32_port, add_in_14_31_port, 
      add_in_14_30_port, add_in_14_29_port, add_in_14_28_port, 
      add_in_14_27_port, add_in_14_26_port, add_in_14_25_port, 
      add_in_14_24_port, add_in_14_23_port, add_in_14_22_port, 
      add_in_14_21_port, add_in_14_20_port, add_in_14_19_port, 
      add_in_14_18_port, add_in_14_17_port, add_in_14_16_port, 
      add_in_14_15_port, add_in_14_14_port, add_in_14_13_port, 
      add_in_14_12_port, add_in_14_11_port, add_in_14_10_port, add_in_14_9_port
      , add_in_14_8_port, add_in_14_7_port, add_in_14_6_port, add_in_14_5_port,
      add_in_14_4_port, add_in_14_3_port, add_in_14_2_port, add_in_14_1_port, 
      add_in_14_0_port, add_in_13_63_port, add_in_13_62_port, add_in_13_61_port
      , add_in_13_60_port, add_in_13_59_port, add_in_13_58_port, 
      add_in_13_57_port, add_in_13_56_port, add_in_13_55_port, 
      add_in_13_54_port, add_in_13_53_port, add_in_13_52_port, 
      add_in_13_51_port, add_in_13_50_port, add_in_13_49_port, 
      add_in_13_48_port, add_in_13_47_port, add_in_13_46_port, 
      add_in_13_45_port, add_in_13_44_port, add_in_13_43_port, 
      add_in_13_42_port, add_in_13_41_port, add_in_13_40_port, 
      add_in_13_39_port, add_in_13_38_port, add_in_13_37_port, 
      add_in_13_36_port, add_in_13_35_port, add_in_13_34_port, 
      add_in_13_33_port, add_in_13_32_port, add_in_13_31_port, 
      add_in_13_30_port, add_in_13_29_port, add_in_13_28_port, 
      add_in_13_27_port, add_in_13_26_port, add_in_13_25_port, 
      add_in_13_24_port, add_in_13_23_port, add_in_13_22_port, 
      add_in_13_21_port, add_in_13_20_port, add_in_13_19_port, 
      add_in_13_18_port, add_in_13_17_port, add_in_13_16_port, 
      add_in_13_15_port, add_in_13_14_port, add_in_13_13_port, 
      add_in_13_12_port, add_in_13_11_port, add_in_13_10_port, add_in_13_9_port
      , add_in_13_8_port, add_in_13_7_port, add_in_13_6_port, add_in_13_5_port,
      add_in_13_4_port, add_in_13_3_port, add_in_13_2_port, add_in_13_1_port, 
      add_in_13_0_port, add_in_12_63_port, add_in_12_62_port, add_in_12_61_port
      , add_in_12_60_port, add_in_12_59_port, add_in_12_58_port, 
      add_in_12_57_port, add_in_12_56_port, add_in_12_55_port, 
      add_in_12_54_port, add_in_12_53_port, add_in_12_52_port, 
      add_in_12_51_port, add_in_12_50_port, add_in_12_49_port, 
      add_in_12_48_port, add_in_12_47_port, add_in_12_46_port, 
      add_in_12_45_port, add_in_12_44_port, add_in_12_43_port, 
      add_in_12_42_port, add_in_12_41_port, add_in_12_40_port, 
      add_in_12_39_port, add_in_12_38_port, add_in_12_37_port, 
      add_in_12_36_port, add_in_12_35_port, add_in_12_34_port, 
      add_in_12_33_port, add_in_12_32_port, add_in_12_31_port, 
      add_in_12_30_port, add_in_12_29_port, add_in_12_28_port, 
      add_in_12_27_port, add_in_12_26_port, add_in_12_25_port, 
      add_in_12_24_port, add_in_12_23_port, add_in_12_22_port, 
      add_in_12_21_port, add_in_12_20_port, add_in_12_19_port, 
      add_in_12_18_port, add_in_12_17_port, add_in_12_16_port, 
      add_in_12_15_port, add_in_12_14_port, add_in_12_13_port, 
      add_in_12_12_port, add_in_12_11_port, add_in_12_10_port, add_in_12_9_port
      , add_in_12_8_port, add_in_12_7_port, add_in_12_6_port, add_in_12_5_port,
      add_in_12_4_port, add_in_12_3_port, add_in_12_2_port, add_in_12_1_port, 
      add_in_12_0_port, add_in_11_63_port, add_in_11_62_port, add_in_11_61_port
      , add_in_11_60_port, add_in_11_59_port, add_in_11_58_port, 
      add_in_11_57_port, add_in_11_56_port, add_in_11_55_port, 
      add_in_11_54_port, add_in_11_53_port, add_in_11_52_port, 
      add_in_11_51_port, add_in_11_50_port, add_in_11_49_port, 
      add_in_11_48_port, add_in_11_47_port, add_in_11_46_port, 
      add_in_11_45_port, add_in_11_44_port, add_in_11_43_port, 
      add_in_11_42_port, add_in_11_41_port, add_in_11_40_port, 
      add_in_11_39_port, add_in_11_38_port, add_in_11_37_port, 
      add_in_11_36_port, add_in_11_35_port, add_in_11_34_port, 
      add_in_11_33_port, add_in_11_32_port, add_in_11_31_port, 
      add_in_11_30_port, add_in_11_29_port, add_in_11_28_port, 
      add_in_11_27_port, add_in_11_26_port, add_in_11_25_port, 
      add_in_11_24_port, add_in_11_23_port, add_in_11_22_port, 
      add_in_11_21_port, add_in_11_20_port, add_in_11_19_port, 
      add_in_11_18_port, add_in_11_17_port, add_in_11_16_port, 
      add_in_11_15_port, add_in_11_14_port, add_in_11_13_port, 
      add_in_11_12_port, add_in_11_11_port, add_in_11_10_port, add_in_11_9_port
      , add_in_11_8_port, add_in_11_7_port, add_in_11_6_port, add_in_11_5_port,
      add_in_11_4_port, add_in_11_3_port, add_in_11_2_port, add_in_11_1_port, 
      add_in_11_0_port, add_in_10_63_port, add_in_10_62_port, add_in_10_61_port
      , add_in_10_60_port, add_in_10_59_port, add_in_10_58_port, 
      add_in_10_57_port, add_in_10_56_port, add_in_10_55_port, 
      add_in_10_54_port, add_in_10_53_port, add_in_10_52_port, 
      add_in_10_51_port, add_in_10_50_port, add_in_10_49_port, 
      add_in_10_48_port, add_in_10_47_port, add_in_10_46_port, 
      add_in_10_45_port, add_in_10_44_port, add_in_10_43_port, 
      add_in_10_42_port, add_in_10_41_port, add_in_10_40_port, 
      add_in_10_39_port, add_in_10_38_port, add_in_10_37_port, 
      add_in_10_36_port, add_in_10_35_port, add_in_10_34_port, 
      add_in_10_33_port, add_in_10_32_port, add_in_10_31_port, 
      add_in_10_30_port, add_in_10_29_port, add_in_10_28_port, 
      add_in_10_27_port, add_in_10_26_port, add_in_10_25_port, 
      add_in_10_24_port, add_in_10_23_port, add_in_10_22_port, 
      add_in_10_21_port, add_in_10_20_port, add_in_10_19_port, 
      add_in_10_18_port, add_in_10_17_port, add_in_10_16_port, 
      add_in_10_15_port, add_in_10_14_port, add_in_10_13_port, 
      add_in_10_12_port, add_in_10_11_port, add_in_10_10_port, add_in_10_9_port
      , add_in_10_8_port, add_in_10_7_port, add_in_10_6_port, add_in_10_5_port,
      add_in_10_4_port, add_in_10_3_port, add_in_10_2_port, add_in_10_1_port, 
      add_in_10_0_port, add_in_9_63_port, add_in_9_62_port, add_in_9_61_port, 
      add_in_9_60_port, add_in_9_59_port, add_in_9_58_port, add_in_9_57_port, 
      add_in_9_56_port, add_in_9_55_port, add_in_9_54_port, add_in_9_53_port, 
      add_in_9_52_port, add_in_9_51_port, add_in_9_50_port, add_in_9_49_port, 
      add_in_9_48_port, add_in_9_47_port, add_in_9_46_port, add_in_9_45_port, 
      add_in_9_44_port, add_in_9_43_port, add_in_9_42_port, add_in_9_41_port, 
      add_in_9_40_port, add_in_9_39_port, add_in_9_38_port, add_in_9_37_port, 
      add_in_9_36_port, add_in_9_35_port, add_in_9_34_port, add_in_9_33_port, 
      add_in_9_32_port, add_in_9_31_port, add_in_9_30_port, add_in_9_29_port, 
      add_in_9_28_port, add_in_9_27_port, add_in_9_26_port, add_in_9_25_port, 
      add_in_9_24_port, add_in_9_23_port, add_in_9_22_port, add_in_9_21_port, 
      add_in_9_20_port, add_in_9_19_port, add_in_9_18_port, add_in_9_17_port, 
      add_in_9_16_port, add_in_9_15_port, add_in_9_14_port, add_in_9_13_port, 
      add_in_9_12_port, add_in_9_11_port, add_in_9_10_port, add_in_9_9_port, 
      add_in_9_8_port, add_in_9_7_port, add_in_9_6_port, add_in_9_5_port, 
      add_in_9_4_port, add_in_9_3_port, add_in_9_2_port, add_in_9_1_port, 
      add_in_9_0_port, add_in_8_63_port, add_in_8_62_port, add_in_8_61_port, 
      add_in_8_60_port, add_in_8_59_port, add_in_8_58_port, add_in_8_57_port, 
      add_in_8_56_port, add_in_8_55_port, add_in_8_54_port, add_in_8_53_port, 
      add_in_8_52_port, add_in_8_51_port, add_in_8_50_port, add_in_8_49_port, 
      add_in_8_48_port, add_in_8_47_port, add_in_8_46_port, add_in_8_45_port, 
      add_in_8_44_port, add_in_8_43_port, add_in_8_42_port, add_in_8_41_port, 
      add_in_8_40_port, add_in_8_39_port, add_in_8_38_port, add_in_8_37_port, 
      add_in_8_36_port, add_in_8_35_port, add_in_8_34_port, add_in_8_33_port, 
      add_in_8_32_port, add_in_8_31_port, add_in_8_30_port, add_in_8_29_port, 
      add_in_8_28_port, add_in_8_27_port, add_in_8_26_port, add_in_8_25_port, 
      add_in_8_24_port, add_in_8_23_port, add_in_8_22_port, add_in_8_21_port, 
      add_in_8_20_port, add_in_8_19_port, add_in_8_18_port, add_in_8_17_port, 
      add_in_8_16_port, add_in_8_15_port, add_in_8_14_port, add_in_8_13_port, 
      add_in_8_12_port, add_in_8_11_port, add_in_8_10_port, add_in_8_9_port, 
      add_in_8_8_port, add_in_8_7_port, add_in_8_6_port, add_in_8_5_port, 
      add_in_8_4_port, add_in_8_3_port, add_in_8_2_port, add_in_8_1_port, 
      add_in_8_0_port, net21306, net21307, net21308, net21309, net21310, 
      net21311, net21312, net21313, net21314, net21315, net21316, net21317, 
      net21318, net21319, net21320, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, 
      n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, 
      n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, 
      n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, 
      n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, 
      n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360, 
      n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, 
      n373, n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, 
      n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, 
      n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, 
      n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, 
      n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, 
      n433, n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, 
      n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, 
      n457, n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, 
      n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, 
      n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, 
      n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, 
      n505, n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, 
      n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, 
      n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, 
      n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, 
      n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, 
      n565, n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, 
      n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, 
      n589, n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, 
      n601, n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, 
      n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, 
      n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, 
      n637, n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, 
      n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, 
      n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, 
      n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, 
      n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, 
      net165111 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   enc_i_0 : BOOTH_ENCODER_4 port map( I(2) => B(1), I(1) => B(0), I(0) => 
                           X_Logic0_port, O(2) => encoder_out_2_port, O(1) => 
                           encoder_out_1_port, O(0) => encoder_out_0_port);
   enc_i_1 : BOOTH_ENCODER_19 port map( I(2) => B(3), I(1) => B(2), I(0) => 
                           B(1), O(2) => encoder_out_5_port, O(1) => 
                           encoder_out_4_port, O(0) => encoder_out_3_port);
   enc_i_2 : BOOTH_ENCODER_18 port map( I(2) => B(5), I(1) => B(4), I(0) => 
                           B(3), O(2) => encoder_out_8_port, O(1) => 
                           encoder_out_7_port, O(0) => encoder_out_6_port);
   enc_i_3 : BOOTH_ENCODER_17 port map( I(2) => B(7), I(1) => B(6), I(0) => 
                           B(5), O(2) => encoder_out_11_port, O(1) => 
                           encoder_out_10_port, O(0) => encoder_out_9_port);
   enc_i_4 : BOOTH_ENCODER_16 port map( I(2) => B(9), I(1) => B(8), I(0) => 
                           B(7), O(2) => encoder_out_14_port, O(1) => 
                           encoder_out_13_port, O(0) => encoder_out_12_port);
   enc_i_5 : BOOTH_ENCODER_15 port map( I(2) => B(11), I(1) => B(10), I(0) => 
                           B(9), O(2) => encoder_out_17_port, O(1) => 
                           encoder_out_16_port, O(0) => encoder_out_15_port);
   enc_i_6 : BOOTH_ENCODER_14 port map( I(2) => B(13), I(1) => B(12), I(0) => 
                           B(11), O(2) => encoder_out_20_port, O(1) => 
                           encoder_out_19_port, O(0) => encoder_out_18_port);
   enc_i_7 : BOOTH_ENCODER_13 port map( I(2) => B(15), I(1) => B(14), I(0) => 
                           B(13), O(2) => encoder_out_23_port, O(1) => 
                           encoder_out_22_port, O(0) => encoder_out_21_port);
   enc_i_8 : BOOTH_ENCODER_12 port map( I(2) => B(17), I(1) => B(16), I(0) => 
                           B(15), O(2) => encoder_out_26_port, O(1) => 
                           encoder_out_25_port, O(0) => encoder_out_24_port);
   enc_i_9 : BOOTH_ENCODER_11 port map( I(2) => B(19), I(1) => B(18), I(0) => 
                           B(17), O(2) => encoder_out_29_port, O(1) => 
                           encoder_out_28_port, O(0) => encoder_out_27_port);
   enc_i_10 : BOOTH_ENCODER_10 port map( I(2) => B(21), I(1) => B(20), I(0) => 
                           B(19), O(2) => encoder_out_32_port, O(1) => 
                           encoder_out_31_port, O(0) => encoder_out_30_port);
   enc_i_11 : BOOTH_ENCODER_9 port map( I(2) => B(23), I(1) => B(22), I(0) => 
                           B(21), O(2) => encoder_out_35_port, O(1) => 
                           encoder_out_34_port, O(0) => encoder_out_33_port);
   enc_i_12 : BOOTH_ENCODER_8 port map( I(2) => B(25), I(1) => B(24), I(0) => 
                           B(23), O(2) => encoder_out_38_port, O(1) => 
                           encoder_out_37_port, O(0) => encoder_out_36_port);
   enc_i_13 : BOOTH_ENCODER_7 port map( I(2) => B(27), I(1) => B(26), I(0) => 
                           B(25), O(2) => encoder_out_41_port, O(1) => 
                           encoder_out_40_port, O(0) => encoder_out_39_port);
   enc_i_14 : BOOTH_ENCODER_6 port map( I(2) => B(29), I(1) => B(28), I(0) => 
                           B(27), O(2) => encoder_out_44_port, O(1) => 
                           encoder_out_43_port, O(0) => encoder_out_42_port);
   enc_i_15 : BOOTH_ENCODER_5 port map( I(2) => B(31), I(1) => B(30), I(0) => 
                           B(29), O(2) => encoder_out_47_port, O(1) => 
                           encoder_out_46_port, O(0) => encoder_out_45_port);
   mux_i_0 : MUX51_GENERIC_N64_0 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n587, B(62) => n587, B(61) 
                           => n587, B(60) => n587, B(59) => n587, B(58) => n587
                           , B(57) => n587, B(56) => n586, B(55) => n586, B(54)
                           => n586, B(53) => n586, B(52) => n586, B(51) => n586
                           , B(50) => n586, B(49) => n585, B(48) => n585, B(47)
                           => n585, B(46) => n585, B(45) => n585, B(44) => n585
                           , B(43) => n585, B(42) => n584, B(41) => n584, B(40)
                           => n584, B(39) => n584, B(38) => n584, B(37) => n584
                           , B(36) => n584, B(35) => n583, B(34) => n583, B(33)
                           => n583, B(32) => n583, B(31) => n583, B(30) => n502
                           , B(29) => n492, B(28) => n482, B(27) => n472, B(26)
                           => n462, B(25) => n452, B(24) => n442, B(23) => n432
                           , B(22) => n422, B(21) => n412, B(20) => n402, B(19)
                           => n392, B(18) => n382, B(17) => n372, B(16) => n362
                           , B(15) => n352, B(14) => n342, B(13) => n332, B(12)
                           => n322, B(11) => n312, B(10) => n302, B(9) => n292,
                           B(8) => n282, B(7) => n272, B(6) => n262, B(5) => 
                           n252, B(4) => n242, B(3) => n232, B(2) => n222, B(1)
                           => n212, B(0) => n202, C(63) => n656, C(62) => n659,
                           C(61) => n659, C(60) => n659, C(59) => n659, C(58) 
                           => n659, C(57) => n659, C(56) => n658, C(55) => n658
                           , C(54) => n658, C(53) => n658, C(52) => n658, C(51)
                           => n658, C(50) => n658, C(49) => n658, C(48) => n657
                           , C(47) => n657, C(46) => n657, C(45) => n657, C(44)
                           => n656, C(43) => n656, C(42) => n656, C(41) => n656
                           , C(40) => n656, C(39) => n656, C(38) => n654, C(37)
                           => n654, C(36) => n654, C(35) => n654, C(34) => n654
                           , C(33) => n654, C(32) => n654, C(31) => n654, C(30)
                           => n505, C(29) => n495, C(28) => n485, C(27) => n475
                           , C(26) => n465, C(25) => n455, C(24) => n445, C(23)
                           => n435, C(22) => n425, C(21) => n415, C(20) => n405
                           , C(19) => n395, C(18) => n385, C(17) => n375, C(16)
                           => n365, C(15) => n355, C(14) => n345, C(13) => n335
                           , C(12) => n325, C(11) => n315, C(10) => n305, C(9) 
                           => n295, C(8) => n285, C(7) => n275, C(6) => n265, 
                           C(5) => n255, C(4) => n245, C(3) => n235, C(2) => 
                           n225, C(1) => n215, C(0) => n205, D(63) => n583, 
                           D(62) => n583, D(61) => n582, D(60) => n582, D(59) 
                           => n582, D(58) => n582, D(57) => n582, D(56) => n582
                           , D(55) => n582, D(54) => n581, D(53) => n581, D(52)
                           => n581, D(51) => n581, D(50) => n581, D(49) => n581
                           , D(48) => n581, D(47) => n580, D(46) => n580, D(45)
                           => n580, D(44) => n580, D(43) => n580, D(42) => n580
                           , D(41) => n580, D(40) => n579, D(39) => n579, D(38)
                           => n579, D(37) => n579, D(36) => n579, D(35) => n579
                           , D(34) => n579, D(33) => n578, D(32) => n578, D(31)
                           => n502, D(30) => n492, D(29) => n482, D(28) => n472
                           , D(27) => n462, D(26) => n452, D(25) => n442, D(24)
                           => n432, D(23) => n422, D(22) => n412, D(21) => n402
                           , D(20) => n392, D(19) => n382, D(18) => n372, D(17)
                           => n362, D(16) => n352, D(15) => n342, D(14) => n332
                           , D(13) => n322, D(12) => n312, D(11) => n302, D(10)
                           => n292, D(9) => n282, D(8) => n272, D(7) => n262, 
                           D(6) => n252, D(5) => n242, D(4) => n232, D(3) => 
                           n222, D(2) => n212, D(1) => n202, D(0) => 
                           X_Logic0_port, E(63) => n666, E(62) => n666, E(61) 
                           => n666, E(60) => n665, E(59) => n665, E(58) => n665
                           , E(57) => n665, E(56) => n665, E(55) => n665, E(54)
                           => n665, E(53) => n665, E(52) => n664, E(51) => n664
                           , E(50) => n664, E(49) => n664, E(48) => n664, E(47)
                           => n663, E(46) => n663, E(45) => n663, E(44) => n663
                           , E(43) => n662, E(42) => n662, E(41) => n662, E(40)
                           => n662, E(39) => n662, E(38) => n662, E(37) => n662
                           , E(36) => n662, E(35) => n662, E(34) => n662, E(33)
                           => n662, E(32) => n661, E(31) => n506, E(30) => n496
                           , E(29) => n486, E(28) => n476, E(27) => n466, E(26)
                           => n456, E(25) => n446, E(24) => n436, E(23) => n426
                           , E(22) => n416, E(21) => n406, E(20) => n396, E(19)
                           => n386, E(18) => n376, E(17) => n366, E(16) => n356
                           , E(15) => n346, E(14) => n336, E(13) => n326, E(12)
                           => n316, E(11) => n306, E(10) => n296, E(9) => n286,
                           E(8) => n276, E(7) => n266, E(6) => n256, E(5) => 
                           n246, E(4) => n236, E(3) => n226, E(2) => n216, E(1)
                           => n206, E(0) => X_Logic1_port, SEL(2) => 
                           encoder_out_2_port, SEL(1) => encoder_out_1_port, 
                           SEL(0) => encoder_out_0_port, Y(63) => 
                           add_in_0_63_port, Y(62) => add_in_0_62_port, Y(61) 
                           => add_in_0_61_port, Y(60) => add_in_0_60_port, 
                           Y(59) => add_in_0_59_port, Y(58) => add_in_0_58_port
                           , Y(57) => add_in_0_57_port, Y(56) => 
                           add_in_0_56_port, Y(55) => add_in_0_55_port, Y(54) 
                           => add_in_0_54_port, Y(53) => add_in_0_53_port, 
                           Y(52) => add_in_0_52_port, Y(51) => add_in_0_51_port
                           , Y(50) => add_in_0_50_port, Y(49) => 
                           add_in_0_49_port, Y(48) => add_in_0_48_port, Y(47) 
                           => add_in_0_47_port, Y(46) => add_in_0_46_port, 
                           Y(45) => add_in_0_45_port, Y(44) => add_in_0_44_port
                           , Y(43) => add_in_0_43_port, Y(42) => 
                           add_in_0_42_port, Y(41) => add_in_0_41_port, Y(40) 
                           => add_in_0_40_port, Y(39) => add_in_0_39_port, 
                           Y(38) => add_in_0_38_port, Y(37) => add_in_0_37_port
                           , Y(36) => add_in_0_36_port, Y(35) => 
                           add_in_0_35_port, Y(34) => add_in_0_34_port, Y(33) 
                           => add_in_0_33_port, Y(32) => add_in_0_32_port, 
                           Y(31) => add_in_0_31_port, Y(30) => add_in_0_30_port
                           , Y(29) => add_in_0_29_port, Y(28) => 
                           add_in_0_28_port, Y(27) => add_in_0_27_port, Y(26) 
                           => add_in_0_26_port, Y(25) => add_in_0_25_port, 
                           Y(24) => add_in_0_24_port, Y(23) => add_in_0_23_port
                           , Y(22) => add_in_0_22_port, Y(21) => 
                           add_in_0_21_port, Y(20) => add_in_0_20_port, Y(19) 
                           => add_in_0_19_port, Y(18) => add_in_0_18_port, 
                           Y(17) => add_in_0_17_port, Y(16) => add_in_0_16_port
                           , Y(15) => add_in_0_15_port, Y(14) => 
                           add_in_0_14_port, Y(13) => add_in_0_13_port, Y(12) 
                           => add_in_0_12_port, Y(11) => add_in_0_11_port, 
                           Y(10) => add_in_0_10_port, Y(9) => add_in_0_9_port, 
                           Y(8) => add_in_0_8_port, Y(7) => add_in_0_7_port, 
                           Y(6) => add_in_0_6_port, Y(5) => add_in_0_5_port, 
                           Y(4) => add_in_0_4_port, Y(3) => add_in_0_3_port, 
                           Y(2) => add_in_0_2_port, Y(1) => add_in_0_1_port, 
                           Y(0) => add_in_0_0_port);
   mux_i_1 : MUX51_GENERIC_N64_15 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n516, B(62) => n516, B(61) 
                           => n516, B(60) => n516, B(59) => n516, B(58) => n515
                           , B(57) => n515, B(56) => n515, B(55) => n515, B(54)
                           => n515, B(53) => n515, B(52) => n515, B(51) => n514
                           , B(50) => n514, B(49) => n514, B(48) => n514, B(47)
                           => n514, B(46) => n514, B(45) => n514, B(44) => n513
                           , B(43) => n513, B(42) => n513, B(41) => n513, B(40)
                           => n513, B(39) => n513, B(38) => n513, B(37) => n512
                           , B(36) => n512, B(35) => n512, B(34) => n512, B(33)
                           => n512, B(32) => n498, B(31) => n488, B(30) => n478
                           , B(29) => n468, B(28) => n458, B(27) => n448, B(26)
                           => n438, B(25) => n428, B(24) => n418, B(23) => n408
                           , B(22) => n398, B(21) => n388, B(20) => n378, B(19)
                           => n368, B(18) => n358, B(17) => n348, B(16) => n338
                           , B(15) => n328, B(14) => n318, B(13) => n308, B(12)
                           => n298, B(11) => n288, B(10) => n278, B(9) => n268,
                           B(8) => n258, B(7) => n248, B(6) => n238, B(5) => 
                           n228, B(4) => n218, B(3) => n208, B(2) => n198, B(1)
                           => X_Logic0_port, B(0) => X_Logic0_port, C(63) => 
                           n653, C(62) => n653, C(61) => n653, C(60) => n653, 
                           C(59) => n653, C(58) => n653, C(57) => n653, C(56) 
                           => n653, C(55) => n653, C(54) => n655, C(53) => n655
                           , C(52) => n655, C(51) => n655, C(50) => n655, C(49)
                           => n658, C(48) => n658, C(47) => n658, C(46) => n658
                           , C(45) => n657, C(44) => n657, C(43) => n657, C(42)
                           => n657, C(41) => n657, C(40) => n657, C(39) => n657
                           , C(38) => n657, C(37) => n656, C(36) => n656, C(35)
                           => n656, C(34) => n656, C(33) => n656, C(32) => n505
                           , C(31) => n495, C(30) => n485, C(29) => n475, C(28)
                           => n465, C(27) => n455, C(26) => n445, C(25) => n435
                           , C(24) => n425, C(23) => n415, C(22) => n405, C(21)
                           => n395, C(20) => n385, C(19) => n375, C(18) => n365
                           , C(17) => n355, C(16) => n345, C(15) => n335, C(14)
                           => n325, C(13) => n315, C(12) => n305, C(11) => n295
                           , C(10) => n285, C(9) => n275, C(8) => n265, C(7) =>
                           n255, C(6) => n245, C(5) => n235, C(4) => n225, C(3)
                           => n215, C(2) => n205, C(1) => X_Logic1_port, C(0) 
                           => X_Logic1_port, D(63) => n512, D(62) => n512, 
                           D(61) => n511, D(60) => n511, D(59) => n511, D(58) 
                           => n511, D(57) => n511, D(56) => n511, D(55) => n511
                           , D(54) => n510, D(53) => n510, D(52) => n510, D(51)
                           => n510, D(50) => n510, D(49) => n510, D(48) => n510
                           , D(47) => n509, D(46) => n509, D(45) => n509, D(44)
                           => n509, D(43) => n509, D(42) => n509, D(41) => n509
                           , D(40) => n508, D(39) => n508, D(38) => n508, D(37)
                           => n508, D(36) => n508, D(35) => n508, D(34) => n508
                           , D(33) => n498, D(32) => n488, D(31) => n478, D(30)
                           => n468, D(29) => n458, D(28) => n448, D(27) => n438
                           , D(26) => n428, D(25) => n418, D(24) => n408, D(23)
                           => n398, D(22) => n388, D(21) => n378, D(20) => n368
                           , D(19) => n358, D(18) => n348, D(17) => n338, D(16)
                           => n328, D(15) => n318, D(14) => n308, D(13) => n298
                           , D(12) => n288, D(11) => n278, D(10) => n268, D(9) 
                           => n258, D(8) => n248, D(7) => n238, D(6) => n228, 
                           D(5) => n218, D(4) => n208, D(3) => n198, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(63) => n680, E(62) => n680, E(61) 
                           => n680, E(60) => n680, E(59) => n678, E(58) => n678
                           , E(57) => n678, E(56) => n678, E(55) => n678, E(54)
                           => n678, E(53) => n678, E(52) => n678, E(51) => n678
                           , E(50) => n678, E(49) => n677, E(48) => n677, E(47)
                           => n677, E(46) => n677, E(45) => n677, E(44) => n677
                           , E(43) => n677, E(42) => n677, E(41) => n677, E(40)
                           => n677, E(39) => n677, E(38) => n675, E(37) => n675
                           , E(36) => n674, E(35) => n674, E(34) => n674, E(33)
                           => n507, E(32) => n497, E(31) => n487, E(30) => n477
                           , E(29) => n467, E(28) => n457, E(27) => n447, E(26)
                           => n437, E(25) => n427, E(24) => n417, E(23) => n407
                           , E(22) => n397, E(21) => n387, E(20) => n377, E(19)
                           => n367, E(18) => n357, E(17) => n347, E(16) => n337
                           , E(15) => n327, E(14) => n317, E(13) => n307, E(12)
                           => n297, E(11) => n287, E(10) => n277, E(9) => n267,
                           E(8) => n257, E(7) => n247, E(6) => n237, E(5) => 
                           n227, E(4) => n217, E(3) => n207, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_5_port, SEL(1) 
                           => encoder_out_4_port, SEL(0) => encoder_out_3_port,
                           Y(63) => mux_out_1_63_port, Y(62) => 
                           mux_out_1_62_port, Y(61) => mux_out_1_61_port, Y(60)
                           => mux_out_1_60_port, Y(59) => mux_out_1_59_port, 
                           Y(58) => mux_out_1_58_port, Y(57) => 
                           mux_out_1_57_port, Y(56) => mux_out_1_56_port, Y(55)
                           => mux_out_1_55_port, Y(54) => mux_out_1_54_port, 
                           Y(53) => mux_out_1_53_port, Y(52) => 
                           mux_out_1_52_port, Y(51) => mux_out_1_51_port, Y(50)
                           => mux_out_1_50_port, Y(49) => mux_out_1_49_port, 
                           Y(48) => mux_out_1_48_port, Y(47) => 
                           mux_out_1_47_port, Y(46) => mux_out_1_46_port, Y(45)
                           => mux_out_1_45_port, Y(44) => mux_out_1_44_port, 
                           Y(43) => mux_out_1_43_port, Y(42) => 
                           mux_out_1_42_port, Y(41) => mux_out_1_41_port, Y(40)
                           => mux_out_1_40_port, Y(39) => mux_out_1_39_port, 
                           Y(38) => mux_out_1_38_port, Y(37) => 
                           mux_out_1_37_port, Y(36) => mux_out_1_36_port, Y(35)
                           => mux_out_1_35_port, Y(34) => mux_out_1_34_port, 
                           Y(33) => mux_out_1_33_port, Y(32) => 
                           mux_out_1_32_port, Y(31) => mux_out_1_31_port, Y(30)
                           => mux_out_1_30_port, Y(29) => mux_out_1_29_port, 
                           Y(28) => mux_out_1_28_port, Y(27) => 
                           mux_out_1_27_port, Y(26) => mux_out_1_26_port, Y(25)
                           => mux_out_1_25_port, Y(24) => mux_out_1_24_port, 
                           Y(23) => mux_out_1_23_port, Y(22) => 
                           mux_out_1_22_port, Y(21) => mux_out_1_21_port, Y(20)
                           => mux_out_1_20_port, Y(19) => mux_out_1_19_port, 
                           Y(18) => mux_out_1_18_port, Y(17) => 
                           mux_out_1_17_port, Y(16) => mux_out_1_16_port, Y(15)
                           => mux_out_1_15_port, Y(14) => mux_out_1_14_port, 
                           Y(13) => mux_out_1_13_port, Y(12) => 
                           mux_out_1_12_port, Y(11) => mux_out_1_11_port, Y(10)
                           => mux_out_1_10_port, Y(9) => mux_out_1_9_port, Y(8)
                           => mux_out_1_8_port, Y(7) => mux_out_1_7_port, Y(6) 
                           => mux_out_1_6_port, Y(5) => mux_out_1_5_port, Y(4) 
                           => mux_out_1_4_port, Y(3) => mux_out_1_3_port, Y(2) 
                           => mux_out_1_2_port, Y(1) => mux_out_1_1_port, Y(0) 
                           => mux_out_1_0_port);
   mux_i_2 : MUX51_GENERIC_N64_14 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n524, B(62) => n524, B(61) 
                           => n524, B(60) => n524, B(59) => n524, B(58) => n524
                           , B(57) => n523, B(56) => n523, B(55) => n523, B(54)
                           => n523, B(53) => n523, B(52) => n523, B(51) => n523
                           , B(50) => n522, B(49) => n522, B(48) => n522, B(47)
                           => n522, B(46) => n522, B(45) => n522, B(44) => n522
                           , B(43) => n521, B(42) => n521, B(41) => n521, B(40)
                           => n521, B(39) => n521, B(38) => n521, B(37) => n521
                           , B(36) => n520, B(35) => n520, B(34) => n498, B(33)
                           => n488, B(32) => n478, B(31) => n468, B(30) => n458
                           , B(29) => n448, B(28) => n438, B(27) => n428, B(26)
                           => n418, B(25) => n408, B(24) => n398, B(23) => n388
                           , B(22) => n378, B(21) => n368, B(20) => n358, B(19)
                           => n348, B(18) => n338, B(17) => n328, B(16) => n318
                           , B(15) => n308, B(14) => n298, B(13) => n288, B(12)
                           => n278, B(11) => n268, B(10) => n258, B(9) => n248,
                           B(8) => n238, B(7) => n228, B(6) => n218, B(5) => 
                           n208, B(4) => n198, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, C(63) => n651, C(62) => n651, C(61) 
                           => n651, C(60) => n652, C(59) => n652, C(58) => n652
                           , C(57) => n652, C(56) => n652, C(55) => n652, C(54)
                           => n652, C(53) => n652, C(52) => n652, C(51) => n652
                           , C(50) => n652, C(49) => n652, C(48) => n653, C(47)
                           => n653, C(46) => n653, C(45) => n654, C(44) => n654
                           , C(43) => n654, C(42) => n654, C(41) => n655, C(40)
                           => n655, C(39) => n655, C(38) => n655, C(37) => n655
                           , C(36) => n655, C(35) => n655, C(34) => n505, C(33)
                           => n495, C(32) => n485, C(31) => n475, C(30) => n465
                           , C(29) => n455, C(28) => n445, C(27) => n435, C(26)
                           => n425, C(25) => n415, C(24) => n405, C(23) => n395
                           , C(22) => n385, C(21) => n375, C(20) => n365, C(19)
                           => n355, C(18) => n345, C(17) => n335, C(16) => n325
                           , C(15) => n315, C(14) => n305, C(13) => n295, C(12)
                           => n285, C(11) => n275, C(10) => n265, C(9) => n255,
                           C(8) => n245, C(7) => n235, C(6) => n225, C(5) => 
                           n215, C(4) => n205, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n520, D(62) => n520, D(61) 
                           => n520, D(60) => n520, D(59) => n520, D(58) => n519
                           , D(57) => n519, D(56) => n519, D(55) => n519, D(54)
                           => n519, D(53) => n519, D(52) => n519, D(51) => n518
                           , D(50) => n518, D(49) => n518, D(48) => n518, D(47)
                           => n518, D(46) => n518, D(45) => n518, D(44) => n517
                           , D(43) => n517, D(42) => n517, D(41) => n517, D(40)
                           => n517, D(39) => n517, D(38) => n517, D(37) => n516
                           , D(36) => n516, D(35) => n498, D(34) => n488, D(33)
                           => n478, D(32) => n468, D(31) => n458, D(30) => n448
                           , D(29) => n438, D(28) => n428, D(27) => n418, D(26)
                           => n408, D(25) => n398, D(24) => n388, D(23) => n378
                           , D(22) => n368, D(21) => n358, D(20) => n348, D(19)
                           => n338, D(18) => n328, D(17) => n318, D(16) => n308
                           , D(15) => n298, D(14) => n288, D(13) => n278, D(12)
                           => n268, D(11) => n258, D(10) => n248, D(9) => n238,
                           D(8) => n228, D(7) => n218, D(6) => n208, D(5) => 
                           n198, D(4) => X_Logic0_port, D(3) => X_Logic0_port, 
                           D(2) => X_Logic0_port, D(1) => X_Logic0_port, D(0) 
                           => X_Logic0_port, E(63) => n668, E(62) => n668, 
                           E(61) => n647, E(60) => n667, E(59) => n666, E(58) 
                           => n650, E(57) => n649, E(56) => n648, E(55) => n651
                           , E(54) => n672, E(53) => n672, E(52) => n672, E(51)
                           => n672, E(50) => n672, E(49) => n670, E(48) => n670
                           , E(47) => n670, E(46) => n670, E(45) => n670, E(44)
                           => n669, E(43) => n669, E(42) => n669, E(41) => n669
                           , E(40) => n669, E(39) => n669, E(38) => n669, E(37)
                           => n675, E(36) => n660, E(35) => n507, E(34) => n497
                           , E(33) => n487, E(32) => n477, E(31) => n467, E(30)
                           => n457, E(29) => n447, E(28) => n437, E(27) => n427
                           , E(26) => n417, E(25) => n407, E(24) => n397, E(23)
                           => n387, E(22) => n377, E(21) => n367, E(20) => n357
                           , E(19) => n347, E(18) => n337, E(17) => n327, E(16)
                           => n317, E(15) => n307, E(14) => n297, E(13) => n287
                           , E(12) => n277, E(11) => n267, E(10) => n257, E(9) 
                           => n247, E(8) => n237, E(7) => n227, E(6) => n217, 
                           E(5) => n207, E(4) => X_Logic1_port, E(3) => 
                           X_Logic1_port, E(2) => X_Logic1_port, E(1) => 
                           X_Logic1_port, E(0) => X_Logic1_port, SEL(2) => 
                           encoder_out_8_port, SEL(1) => encoder_out_7_port, 
                           SEL(0) => encoder_out_6_port, Y(63) => 
                           mux_out_2_63_port, Y(62) => mux_out_2_62_port, Y(61)
                           => mux_out_2_61_port, Y(60) => mux_out_2_60_port, 
                           Y(59) => mux_out_2_59_port, Y(58) => 
                           mux_out_2_58_port, Y(57) => mux_out_2_57_port, Y(56)
                           => mux_out_2_56_port, Y(55) => mux_out_2_55_port, 
                           Y(54) => mux_out_2_54_port, Y(53) => 
                           mux_out_2_53_port, Y(52) => mux_out_2_52_port, Y(51)
                           => mux_out_2_51_port, Y(50) => mux_out_2_50_port, 
                           Y(49) => mux_out_2_49_port, Y(48) => 
                           mux_out_2_48_port, Y(47) => mux_out_2_47_port, Y(46)
                           => mux_out_2_46_port, Y(45) => mux_out_2_45_port, 
                           Y(44) => mux_out_2_44_port, Y(43) => 
                           mux_out_2_43_port, Y(42) => mux_out_2_42_port, Y(41)
                           => mux_out_2_41_port, Y(40) => mux_out_2_40_port, 
                           Y(39) => mux_out_2_39_port, Y(38) => 
                           mux_out_2_38_port, Y(37) => mux_out_2_37_port, Y(36)
                           => mux_out_2_36_port, Y(35) => mux_out_2_35_port, 
                           Y(34) => mux_out_2_34_port, Y(33) => 
                           mux_out_2_33_port, Y(32) => mux_out_2_32_port, Y(31)
                           => mux_out_2_31_port, Y(30) => mux_out_2_30_port, 
                           Y(29) => mux_out_2_29_port, Y(28) => 
                           mux_out_2_28_port, Y(27) => mux_out_2_27_port, Y(26)
                           => mux_out_2_26_port, Y(25) => mux_out_2_25_port, 
                           Y(24) => mux_out_2_24_port, Y(23) => 
                           mux_out_2_23_port, Y(22) => mux_out_2_22_port, Y(21)
                           => mux_out_2_21_port, Y(20) => mux_out_2_20_port, 
                           Y(19) => mux_out_2_19_port, Y(18) => 
                           mux_out_2_18_port, Y(17) => mux_out_2_17_port, Y(16)
                           => mux_out_2_16_port, Y(15) => mux_out_2_15_port, 
                           Y(14) => mux_out_2_14_port, Y(13) => 
                           mux_out_2_13_port, Y(12) => mux_out_2_12_port, Y(11)
                           => mux_out_2_11_port, Y(10) => mux_out_2_10_port, 
                           Y(9) => mux_out_2_9_port, Y(8) => mux_out_2_8_port, 
                           Y(7) => mux_out_2_7_port, Y(6) => mux_out_2_6_port, 
                           Y(5) => mux_out_2_5_port, Y(4) => mux_out_2_4_port, 
                           Y(3) => mux_out_2_3_port, Y(2) => mux_out_2_2_port, 
                           Y(1) => mux_out_2_1_port, Y(0) => mux_out_2_0_port);
   mux_i_3 : MUX51_GENERIC_N64_13 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n532, B(62) => n532, B(61) 
                           => n532, B(60) => n531, B(59) => n531, B(58) => n531
                           , B(57) => n531, B(56) => n531, B(55) => n531, B(54)
                           => n531, B(53) => n530, B(52) => n530, B(51) => n530
                           , B(50) => n530, B(49) => n530, B(48) => n530, B(47)
                           => n530, B(46) => n529, B(45) => n529, B(44) => n529
                           , B(43) => n529, B(42) => n529, B(41) => n529, B(40)
                           => n529, B(39) => n528, B(38) => n528, B(37) => n528
                           , B(36) => n498, B(35) => n488, B(34) => n478, B(33)
                           => n468, B(32) => n458, B(31) => n448, B(30) => n438
                           , B(29) => n428, B(28) => n418, B(27) => n408, B(26)
                           => n398, B(25) => n388, B(24) => n378, B(23) => n368
                           , B(22) => n358, B(21) => n348, B(20) => n338, B(19)
                           => n328, B(18) => n318, B(17) => n308, B(16) => n298
                           , B(15) => n288, B(14) => n278, B(13) => n268, B(12)
                           => n258, B(11) => n248, B(10) => n238, B(9) => n228,
                           B(8) => n218, B(7) => n208, B(6) => n198, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(63) => n659,
                           C(62) => n659, C(61) => n659, C(60) => n659, C(59) 
                           => n659, C(58) => n659, C(57) => n643, C(56) => n636
                           , C(55) => n636, C(54) => n636, C(53) => n636, C(52)
                           => n636, C(51) => n636, C(50) => n636, C(49) => n636
                           , C(48) => n636, C(47) => n636, C(46) => n636, C(45)
                           => n637, C(44) => n637, C(43) => n637, C(42) => n637
                           , C(41) => n637, C(40) => n637, C(39) => n637, C(38)
                           => n637, C(37) => n637, C(36) => n505, C(35) => n495
                           , C(34) => n485, C(33) => n475, C(32) => n465, C(31)
                           => n455, C(30) => n445, C(29) => n435, C(28) => n425
                           , C(27) => n415, C(26) => n405, C(25) => n395, C(24)
                           => n385, C(23) => n375, C(22) => n365, C(21) => n355
                           , C(20) => n345, C(19) => n335, C(18) => n325, C(17)
                           => n315, C(16) => n305, C(15) => n295, C(14) => n285
                           , C(13) => n275, C(12) => n265, C(11) => n255, C(10)
                           => n245, C(9) => n235, C(8) => n225, C(7) => n215, 
                           C(6) => n205, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n528, D(62) => n528, D(61) 
                           => n528, D(60) => n528, D(59) => n527, D(58) => n527
                           , D(57) => n527, D(56) => n527, D(55) => n527, D(54)
                           => n527, D(53) => n527, D(52) => n526, D(51) => n526
                           , D(50) => n526, D(49) => n526, D(48) => n526, D(47)
                           => n526, D(46) => n526, D(45) => n525, D(44) => n525
                           , D(43) => n525, D(42) => n525, D(41) => n525, D(40)
                           => n525, D(39) => n525, D(38) => n524, D(37) => n498
                           , D(36) => n488, D(35) => n478, D(34) => n468, D(33)
                           => n458, D(32) => n448, D(31) => n438, D(30) => n428
                           , D(29) => n418, D(28) => n408, D(27) => n398, D(26)
                           => n388, D(25) => n378, D(24) => n368, D(23) => n358
                           , D(22) => n348, D(21) => n338, D(20) => n328, D(19)
                           => n318, D(18) => n308, D(17) => n298, D(16) => n288
                           , D(15) => n278, D(14) => n268, D(13) => n258, D(12)
                           => n248, D(11) => n238, D(10) => n228, D(9) => n218,
                           D(8) => n208, D(7) => n198, D(6) => X_Logic0_port, 
                           D(5) => X_Logic0_port, D(4) => X_Logic0_port, D(3) 
                           => X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, E(63) => n670,
                           E(62) => n670, E(61) => n670, E(60) => n670, E(59) 
                           => n670, E(58) => n670, E(57) => n670, E(56) => n671
                           , E(55) => n671, E(54) => n671, E(53) => n671, E(52)
                           => n671, E(51) => n671, E(50) => n671, E(49) => n671
                           , E(48) => n671, E(47) => n671, E(46) => n671, E(45)
                           => n671, E(44) => n672, E(43) => n672, E(42) => n672
                           , E(41) => n672, E(40) => n672, E(39) => n672, E(38)
                           => n672, E(37) => n507, E(36) => n497, E(35) => n487
                           , E(34) => n477, E(33) => n467, E(32) => n457, E(31)
                           => n447, E(30) => n437, E(29) => n427, E(28) => n417
                           , E(27) => n407, E(26) => n397, E(25) => n387, E(24)
                           => n377, E(23) => n367, E(22) => n357, E(21) => n347
                           , E(20) => n337, E(19) => n327, E(18) => n317, E(17)
                           => n307, E(16) => n297, E(15) => n287, E(14) => n277
                           , E(13) => n267, E(12) => n257, E(11) => n247, E(10)
                           => n237, E(9) => n227, E(8) => n217, E(7) => n207, 
                           E(6) => X_Logic1_port, E(5) => X_Logic1_port, E(4) 
                           => X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_11_port, SEL(1)
                           => encoder_out_10_port, SEL(0) => encoder_out_9_port
                           , Y(63) => mux_out_3_63_port, Y(62) => 
                           mux_out_3_62_port, Y(61) => mux_out_3_61_port, Y(60)
                           => mux_out_3_60_port, Y(59) => mux_out_3_59_port, 
                           Y(58) => mux_out_3_58_port, Y(57) => 
                           mux_out_3_57_port, Y(56) => mux_out_3_56_port, Y(55)
                           => mux_out_3_55_port, Y(54) => mux_out_3_54_port, 
                           Y(53) => mux_out_3_53_port, Y(52) => 
                           mux_out_3_52_port, Y(51) => mux_out_3_51_port, Y(50)
                           => mux_out_3_50_port, Y(49) => mux_out_3_49_port, 
                           Y(48) => mux_out_3_48_port, Y(47) => 
                           mux_out_3_47_port, Y(46) => mux_out_3_46_port, Y(45)
                           => mux_out_3_45_port, Y(44) => mux_out_3_44_port, 
                           Y(43) => mux_out_3_43_port, Y(42) => 
                           mux_out_3_42_port, Y(41) => mux_out_3_41_port, Y(40)
                           => mux_out_3_40_port, Y(39) => mux_out_3_39_port, 
                           Y(38) => mux_out_3_38_port, Y(37) => 
                           mux_out_3_37_port, Y(36) => mux_out_3_36_port, Y(35)
                           => mux_out_3_35_port, Y(34) => mux_out_3_34_port, 
                           Y(33) => mux_out_3_33_port, Y(32) => 
                           mux_out_3_32_port, Y(31) => mux_out_3_31_port, Y(30)
                           => mux_out_3_30_port, Y(29) => mux_out_3_29_port, 
                           Y(28) => mux_out_3_28_port, Y(27) => 
                           mux_out_3_27_port, Y(26) => mux_out_3_26_port, Y(25)
                           => mux_out_3_25_port, Y(24) => mux_out_3_24_port, 
                           Y(23) => mux_out_3_23_port, Y(22) => 
                           mux_out_3_22_port, Y(21) => mux_out_3_21_port, Y(20)
                           => mux_out_3_20_port, Y(19) => mux_out_3_19_port, 
                           Y(18) => mux_out_3_18_port, Y(17) => 
                           mux_out_3_17_port, Y(16) => mux_out_3_16_port, Y(15)
                           => mux_out_3_15_port, Y(14) => mux_out_3_14_port, 
                           Y(13) => mux_out_3_13_port, Y(12) => 
                           mux_out_3_12_port, Y(11) => mux_out_3_11_port, Y(10)
                           => mux_out_3_10_port, Y(9) => mux_out_3_9_port, Y(8)
                           => mux_out_3_8_port, Y(7) => mux_out_3_7_port, Y(6) 
                           => mux_out_3_6_port, Y(5) => mux_out_3_5_port, Y(4) 
                           => mux_out_3_4_port, Y(3) => mux_out_3_3_port, Y(2) 
                           => mux_out_3_2_port, Y(1) => mux_out_3_1_port, Y(0) 
                           => mux_out_3_0_port);
   mux_i_4 : MUX51_GENERIC_N64_12 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n539, B(62) => n539, B(61) 
                           => n539, B(60) => n538, B(59) => n538, B(58) => n538
                           , B(57) => n538, B(56) => n538, B(55) => n538, B(54)
                           => n538, B(53) => n537, B(52) => n537, B(51) => n537
                           , B(50) => n537, B(49) => n537, B(48) => n537, B(47)
                           => n537, B(46) => n536, B(45) => n536, B(44) => n536
                           , B(43) => n536, B(42) => n536, B(41) => n536, B(40)
                           => n536, B(39) => n535, B(38) => n499, B(37) => n489
                           , B(36) => n479, B(35) => n469, B(34) => n459, B(33)
                           => n449, B(32) => n439, B(31) => n429, B(30) => n419
                           , B(29) => n409, B(28) => n399, B(27) => n389, B(26)
                           => n379, B(25) => n369, B(24) => n359, B(23) => n349
                           , B(22) => n339, B(21) => n329, B(20) => n319, B(19)
                           => n309, B(18) => n299, B(17) => n289, B(16) => n279
                           , B(15) => n269, B(14) => n259, B(13) => n249, B(12)
                           => n239, B(11) => n229, B(10) => n219, B(9) => n209,
                           B(8) => n199, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, C(63) => n637, C(62) => n637, C(61) 
                           => n637, C(60) => n638, C(59) => n638, C(58) => n638
                           , C(57) => n638, C(56) => n638, C(55) => n638, C(54)
                           => n638, C(53) => n638, C(52) => n638, C(51) => n638
                           , C(50) => n638, C(49) => n638, C(48) => n639, C(47)
                           => n639, C(46) => n639, C(45) => n639, C(44) => n639
                           , C(43) => n639, C(42) => n639, C(41) => n639, C(40)
                           => n639, C(39) => n639, C(38) => n505, C(37) => n495
                           , C(36) => n485, C(35) => n475, C(34) => n465, C(33)
                           => n455, C(32) => n445, C(31) => n435, C(30) => n425
                           , C(29) => n415, C(28) => n405, C(27) => n395, C(26)
                           => n385, C(25) => n375, C(24) => n365, C(23) => n355
                           , C(22) => n345, C(21) => n335, C(20) => n325, C(19)
                           => n315, C(18) => n305, C(17) => n295, C(16) => n285
                           , C(15) => n275, C(14) => n265, C(13) => n255, C(12)
                           => n245, C(11) => n235, C(10) => n225, C(9) => n215,
                           C(8) => n205, C(7) => X_Logic1_port, C(6) => 
                           X_Logic1_port, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n535, D(62) => n535, D(61) 
                           => n535, D(60) => n535, D(59) => n535, D(58) => n535
                           , D(57) => n534, D(56) => n534, D(55) => n534, D(54)
                           => n534, D(53) => n534, D(52) => n534, D(51) => n534
                           , D(50) => n533, D(49) => n533, D(48) => n533, D(47)
                           => n533, D(46) => n533, D(45) => n533, D(44) => n533
                           , D(43) => n532, D(42) => n532, D(41) => n532, D(40)
                           => n532, D(39) => n498, D(38) => n488, D(37) => n478
                           , D(36) => n468, D(35) => n458, D(34) => n448, D(33)
                           => n438, D(32) => n428, D(31) => n418, D(30) => n408
                           , D(29) => n398, D(28) => n388, D(27) => n378, D(26)
                           => n368, D(25) => n358, D(24) => n348, D(23) => n338
                           , D(22) => n328, D(21) => n318, D(20) => n308, D(19)
                           => n298, D(18) => n288, D(17) => n278, D(16) => n268
                           , D(15) => n258, D(14) => n248, D(13) => n238, D(12)
                           => n228, D(11) => n218, D(10) => n208, D(9) => n198,
                           D(8) => X_Logic0_port, D(7) => X_Logic0_port, D(6) 
                           => X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(63) => n668, E(62) => n668, E(61) 
                           => n668, E(60) => n673, E(59) => n673, E(58) => n673
                           , E(57) => n673, E(56) => n673, E(55) => n673, E(54)
                           => n673, E(53) => n673, E(52) => n673, E(51) => n673
                           , E(50) => n673, E(49) => n673, E(48) => n674, E(47)
                           => n674, E(46) => n674, E(45) => n674, E(44) => n674
                           , E(43) => n674, E(42) => n674, E(41) => n674, E(40)
                           => n674, E(39) => n507, E(38) => n497, E(37) => n487
                           , E(36) => n477, E(35) => n467, E(34) => n457, E(33)
                           => n447, E(32) => n437, E(31) => n427, E(30) => n417
                           , E(29) => n407, E(28) => n397, E(27) => n387, E(26)
                           => n377, E(25) => n367, E(24) => n357, E(23) => n347
                           , E(22) => n337, E(21) => n327, E(20) => n317, E(19)
                           => n307, E(18) => n297, E(17) => n287, E(16) => n277
                           , E(15) => n267, E(14) => n257, E(13) => n247, E(12)
                           => n237, E(11) => n227, E(10) => n217, E(9) => n207,
                           E(8) => X_Logic1_port, E(7) => X_Logic1_port, E(6) 
                           => X_Logic1_port, E(5) => X_Logic1_port, E(4) => 
                           X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_14_port, SEL(1)
                           => encoder_out_13_port, SEL(0) => 
                           encoder_out_12_port, Y(63) => mux_out_4_63_port, 
                           Y(62) => mux_out_4_62_port, Y(61) => 
                           mux_out_4_61_port, Y(60) => mux_out_4_60_port, Y(59)
                           => mux_out_4_59_port, Y(58) => mux_out_4_58_port, 
                           Y(57) => mux_out_4_57_port, Y(56) => 
                           mux_out_4_56_port, Y(55) => mux_out_4_55_port, Y(54)
                           => mux_out_4_54_port, Y(53) => mux_out_4_53_port, 
                           Y(52) => mux_out_4_52_port, Y(51) => 
                           mux_out_4_51_port, Y(50) => mux_out_4_50_port, Y(49)
                           => mux_out_4_49_port, Y(48) => mux_out_4_48_port, 
                           Y(47) => mux_out_4_47_port, Y(46) => 
                           mux_out_4_46_port, Y(45) => mux_out_4_45_port, Y(44)
                           => mux_out_4_44_port, Y(43) => mux_out_4_43_port, 
                           Y(42) => mux_out_4_42_port, Y(41) => 
                           mux_out_4_41_port, Y(40) => mux_out_4_40_port, Y(39)
                           => mux_out_4_39_port, Y(38) => mux_out_4_38_port, 
                           Y(37) => mux_out_4_37_port, Y(36) => 
                           mux_out_4_36_port, Y(35) => mux_out_4_35_port, Y(34)
                           => mux_out_4_34_port, Y(33) => mux_out_4_33_port, 
                           Y(32) => mux_out_4_32_port, Y(31) => 
                           mux_out_4_31_port, Y(30) => mux_out_4_30_port, Y(29)
                           => mux_out_4_29_port, Y(28) => mux_out_4_28_port, 
                           Y(27) => mux_out_4_27_port, Y(26) => 
                           mux_out_4_26_port, Y(25) => mux_out_4_25_port, Y(24)
                           => mux_out_4_24_port, Y(23) => mux_out_4_23_port, 
                           Y(22) => mux_out_4_22_port, Y(21) => 
                           mux_out_4_21_port, Y(20) => mux_out_4_20_port, Y(19)
                           => mux_out_4_19_port, Y(18) => mux_out_4_18_port, 
                           Y(17) => mux_out_4_17_port, Y(16) => 
                           mux_out_4_16_port, Y(15) => mux_out_4_15_port, Y(14)
                           => mux_out_4_14_port, Y(13) => mux_out_4_13_port, 
                           Y(12) => mux_out_4_12_port, Y(11) => 
                           mux_out_4_11_port, Y(10) => mux_out_4_10_port, Y(9) 
                           => mux_out_4_9_port, Y(8) => mux_out_4_8_port, Y(7) 
                           => mux_out_4_7_port, Y(6) => mux_out_4_6_port, Y(5) 
                           => mux_out_4_5_port, Y(4) => mux_out_4_4_port, Y(3) 
                           => mux_out_4_3_port, Y(2) => mux_out_4_2_port, Y(1) 
                           => mux_out_4_1_port, Y(0) => mux_out_4_0_port);
   mux_i_5 : MUX51_GENERIC_N64_11 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n545, B(62) => n545, B(61) 
                           => n545, B(60) => n545, B(59) => n545, B(58) => n545
                           , B(57) => n544, B(56) => n544, B(55) => n544, B(54)
                           => n544, B(53) => n544, B(52) => n544, B(51) => n544
                           , B(50) => n543, B(49) => n543, B(48) => n543, B(47)
                           => n543, B(46) => n543, B(45) => n543, B(44) => n543
                           , B(43) => n542, B(42) => n542, B(41) => n542, B(40)
                           => n499, B(39) => n489, B(38) => n479, B(37) => n469
                           , B(36) => n459, B(35) => n449, B(34) => n439, B(33)
                           => n429, B(32) => n419, B(31) => n409, B(30) => n399
                           , B(29) => n389, B(28) => n379, B(27) => n369, B(26)
                           => n359, B(25) => n349, B(24) => n339, B(23) => n329
                           , B(22) => n319, B(21) => n309, B(20) => n299, B(19)
                           => n289, B(18) => n279, B(17) => n269, B(16) => n259
                           , B(15) => n249, B(14) => n239, B(13) => n229, B(12)
                           => n219, B(11) => n209, B(10) => n199, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(63) => n639,
                           C(62) => n639, C(61) => n640, C(60) => n640, C(59) 
                           => n640, C(58) => n640, C(57) => n640, C(56) => n640
                           , C(55) => n640, C(54) => n640, C(53) => n640, C(52)
                           => n640, C(51) => n640, C(50) => n640, C(49) => n641
                           , C(48) => n641, C(47) => n641, C(46) => n641, C(45)
                           => n641, C(44) => n641, C(43) => n641, C(42) => n641
                           , C(41) => n641, C(40) => n505, C(39) => n495, C(38)
                           => n485, C(37) => n475, C(36) => n465, C(35) => n455
                           , C(34) => n445, C(33) => n435, C(32) => n425, C(31)
                           => n415, C(30) => n405, C(29) => n395, C(28) => n385
                           , C(27) => n375, C(26) => n365, C(25) => n355, C(24)
                           => n345, C(23) => n335, C(22) => n325, C(21) => n315
                           , C(20) => n305, C(19) => n295, C(18) => n285, C(17)
                           => n275, C(16) => n265, C(15) => n255, C(14) => n245
                           , C(13) => n235, C(12) => n225, C(11) => n215, C(10)
                           => n205, C(9) => X_Logic1_port, C(8) => 
                           X_Logic1_port, C(7) => X_Logic1_port, C(6) => 
                           X_Logic1_port, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n542, D(62) => n542, D(61) 
                           => n542, D(60) => n542, D(59) => n541, D(58) => n541
                           , D(57) => n541, D(56) => n541, D(55) => n541, D(54)
                           => n541, D(53) => n541, D(52) => n540, D(51) => n540
                           , D(50) => n540, D(49) => n540, D(48) => n540, D(47)
                           => n540, D(46) => n540, D(45) => n539, D(44) => n539
                           , D(43) => n539, D(42) => n539, D(41) => n499, D(40)
                           => n489, D(39) => n479, D(38) => n469, D(37) => n459
                           , D(36) => n449, D(35) => n439, D(34) => n429, D(33)
                           => n419, D(32) => n409, D(31) => n399, D(30) => n389
                           , D(29) => n379, D(28) => n369, D(27) => n359, D(26)
                           => n349, D(25) => n339, D(24) => n329, D(23) => n319
                           , D(22) => n309, D(21) => n299, D(20) => n289, D(19)
                           => n279, D(18) => n269, D(17) => n259, D(16) => n249
                           , D(15) => n239, D(14) => n229, D(13) => n219, D(12)
                           => n209, D(11) => n199, D(10) => X_Logic0_port, D(9)
                           => X_Logic0_port, D(8) => X_Logic0_port, D(7) => 
                           X_Logic0_port, D(6) => X_Logic0_port, D(5) => 
                           X_Logic0_port, D(4) => X_Logic0_port, D(3) => 
                           X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, E(63) => n675,
                           E(62) => n675, E(61) => n675, E(60) => n675, E(59) 
                           => n675, E(58) => n675, E(57) => n675, E(56) => n675
                           , E(55) => n675, E(54) => n676, E(53) => n676, E(52)
                           => n676, E(51) => n676, E(50) => n676, E(49) => n676
                           , E(48) => n676, E(47) => n676, E(46) => n676, E(45)
                           => n676, E(44) => n676, E(43) => n676, E(42) => n677
                           , E(41) => n507, E(40) => n497, E(39) => n487, E(38)
                           => n477, E(37) => n467, E(36) => n457, E(35) => n447
                           , E(34) => n437, E(33) => n427, E(32) => n417, E(31)
                           => n407, E(30) => n397, E(29) => n387, E(28) => n377
                           , E(27) => n367, E(26) => n357, E(25) => n347, E(24)
                           => n337, E(23) => n327, E(22) => n317, E(21) => n307
                           , E(20) => n297, E(19) => n287, E(18) => n277, E(17)
                           => n267, E(16) => n257, E(15) => n247, E(14) => n237
                           , E(13) => n227, E(12) => n217, E(11) => n207, E(10)
                           => X_Logic1_port, E(9) => X_Logic1_port, E(8) => 
                           X_Logic1_port, E(7) => X_Logic1_port, E(6) => 
                           X_Logic1_port, E(5) => X_Logic1_port, E(4) => 
                           X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_17_port, SEL(1)
                           => encoder_out_16_port, SEL(0) => 
                           encoder_out_15_port, Y(63) => mux_out_5_63_port, 
                           Y(62) => mux_out_5_62_port, Y(61) => 
                           mux_out_5_61_port, Y(60) => mux_out_5_60_port, Y(59)
                           => mux_out_5_59_port, Y(58) => mux_out_5_58_port, 
                           Y(57) => mux_out_5_57_port, Y(56) => 
                           mux_out_5_56_port, Y(55) => mux_out_5_55_port, Y(54)
                           => mux_out_5_54_port, Y(53) => mux_out_5_53_port, 
                           Y(52) => mux_out_5_52_port, Y(51) => 
                           mux_out_5_51_port, Y(50) => mux_out_5_50_port, Y(49)
                           => mux_out_5_49_port, Y(48) => mux_out_5_48_port, 
                           Y(47) => mux_out_5_47_port, Y(46) => 
                           mux_out_5_46_port, Y(45) => mux_out_5_45_port, Y(44)
                           => mux_out_5_44_port, Y(43) => mux_out_5_43_port, 
                           Y(42) => mux_out_5_42_port, Y(41) => 
                           mux_out_5_41_port, Y(40) => mux_out_5_40_port, Y(39)
                           => mux_out_5_39_port, Y(38) => mux_out_5_38_port, 
                           Y(37) => mux_out_5_37_port, Y(36) => 
                           mux_out_5_36_port, Y(35) => mux_out_5_35_port, Y(34)
                           => mux_out_5_34_port, Y(33) => mux_out_5_33_port, 
                           Y(32) => mux_out_5_32_port, Y(31) => 
                           mux_out_5_31_port, Y(30) => mux_out_5_30_port, Y(29)
                           => mux_out_5_29_port, Y(28) => mux_out_5_28_port, 
                           Y(27) => mux_out_5_27_port, Y(26) => 
                           mux_out_5_26_port, Y(25) => mux_out_5_25_port, Y(24)
                           => mux_out_5_24_port, Y(23) => mux_out_5_23_port, 
                           Y(22) => mux_out_5_22_port, Y(21) => 
                           mux_out_5_21_port, Y(20) => mux_out_5_20_port, Y(19)
                           => mux_out_5_19_port, Y(18) => mux_out_5_18_port, 
                           Y(17) => mux_out_5_17_port, Y(16) => 
                           mux_out_5_16_port, Y(15) => mux_out_5_15_port, Y(14)
                           => mux_out_5_14_port, Y(13) => mux_out_5_13_port, 
                           Y(12) => mux_out_5_12_port, Y(11) => 
                           mux_out_5_11_port, Y(10) => mux_out_5_10_port, Y(9) 
                           => mux_out_5_9_port, Y(8) => mux_out_5_8_port, Y(7) 
                           => mux_out_5_7_port, Y(6) => mux_out_5_6_port, Y(5) 
                           => mux_out_5_5_port, Y(4) => mux_out_5_4_port, Y(3) 
                           => mux_out_5_3_port, Y(2) => mux_out_5_2_port, Y(1) 
                           => mux_out_5_1_port, Y(0) => mux_out_5_0_port);
   mux_i_6 : MUX51_GENERIC_N64_10 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n551, B(62) => n551, B(61) 
                           => n551, B(60) => n551, B(59) => n551, B(58) => n550
                           , B(57) => n550, B(56) => n550, B(55) => n550, B(54)
                           => n550, B(53) => n550, B(52) => n550, B(51) => n549
                           , B(50) => n549, B(49) => n549, B(48) => n549, B(47)
                           => n549, B(46) => n549, B(45) => n549, B(44) => n548
                           , B(43) => n548, B(42) => n499, B(41) => n489, B(40)
                           => n479, B(39) => n469, B(38) => n459, B(37) => n449
                           , B(36) => n439, B(35) => n429, B(34) => n419, B(33)
                           => n409, B(32) => n399, B(31) => n389, B(30) => n379
                           , B(29) => n369, B(28) => n359, B(27) => n349, B(26)
                           => n339, B(25) => n329, B(24) => n319, B(23) => n309
                           , B(22) => n299, B(21) => n289, B(20) => n279, B(19)
                           => n269, B(18) => n259, B(17) => n249, B(16) => n239
                           , B(15) => n229, B(14) => n219, B(13) => n209, B(12)
                           => n199, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, C(63) => n641, C(62) => n641, C(61) 
                           => n641, C(60) => n642, C(59) => n642, C(58) => n642
                           , C(57) => n642, C(56) => n642, C(55) => n642, C(54)
                           => n642, C(53) => n642, C(52) => n642, C(51) => n642
                           , C(50) => n642, C(49) => n642, C(48) => n643, C(47)
                           => n643, C(46) => n643, C(45) => n643, C(44) => n643
                           , C(43) => n643, C(42) => n505, C(41) => n495, C(40)
                           => n485, C(39) => n475, C(38) => n465, C(37) => n455
                           , C(36) => n445, C(35) => n435, C(34) => n425, C(33)
                           => n415, C(32) => n405, C(31) => n395, C(30) => n385
                           , C(29) => n375, C(28) => n365, C(27) => n355, C(26)
                           => n345, C(25) => n335, C(24) => n325, C(23) => n315
                           , C(22) => n305, C(21) => n295, C(20) => n285, C(19)
                           => n275, C(18) => n265, C(17) => n255, C(16) => n245
                           , C(15) => n235, C(14) => n225, C(13) => n215, C(12)
                           => n205, C(11) => X_Logic1_port, C(10) => 
                           X_Logic1_port, C(9) => X_Logic1_port, C(8) => 
                           X_Logic1_port, C(7) => X_Logic1_port, C(6) => 
                           X_Logic1_port, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n548, D(62) => n548, D(61) 
                           => n548, D(60) => n548, D(59) => n548, D(58) => n547
                           , D(57) => n547, D(56) => n547, D(55) => n547, D(54)
                           => n547, D(53) => n547, D(52) => n547, D(51) => n546
                           , D(50) => n546, D(49) => n546, D(48) => n546, D(47)
                           => n546, D(46) => n546, D(45) => n546, D(44) => n545
                           , D(43) => n499, D(42) => n489, D(41) => n479, D(40)
                           => n469, D(39) => n459, D(38) => n449, D(37) => n439
                           , D(36) => n429, D(35) => n419, D(34) => n409, D(33)
                           => n399, D(32) => n389, D(31) => n379, D(30) => n369
                           , D(29) => n359, D(28) => n349, D(27) => n339, D(26)
                           => n329, D(25) => n319, D(24) => n309, D(23) => n299
                           , D(22) => n289, D(21) => n279, D(20) => n269, D(19)
                           => n259, D(18) => n249, D(17) => n239, D(16) => n229
                           , D(15) => n219, D(14) => n209, D(13) => n199, D(12)
                           => X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(63) => n678, E(62) => n678, E(61) 
                           => n679, E(60) => n679, E(59) => n679, E(58) => n679
                           , E(57) => n679, E(56) => n679, E(55) => n679, E(54)
                           => n679, E(53) => n679, E(52) => n679, E(51) => n679
                           , E(50) => n679, E(49) => n680, E(48) => n680, E(47)
                           => n680, E(46) => n680, E(45) => n680, E(44) => n680
                           , E(43) => n507, E(42) => n497, E(41) => n487, E(40)
                           => n477, E(39) => n467, E(38) => n457, E(37) => n447
                           , E(36) => n437, E(35) => n427, E(34) => n417, E(33)
                           => n407, E(32) => n397, E(31) => n387, E(30) => n377
                           , E(29) => n367, E(28) => n357, E(27) => n347, E(26)
                           => n337, E(25) => n327, E(24) => n317, E(23) => n307
                           , E(22) => n297, E(21) => n287, E(20) => n277, E(19)
                           => n267, E(18) => n257, E(17) => n247, E(16) => n237
                           , E(15) => n227, E(14) => n217, E(13) => n207, E(12)
                           => X_Logic1_port, E(11) => X_Logic1_port, E(10) => 
                           X_Logic1_port, E(9) => X_Logic1_port, E(8) => 
                           X_Logic1_port, E(7) => X_Logic1_port, E(6) => 
                           X_Logic1_port, E(5) => X_Logic1_port, E(4) => 
                           X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_20_port, SEL(1)
                           => encoder_out_19_port, SEL(0) => 
                           encoder_out_18_port, Y(63) => mux_out_6_63_port, 
                           Y(62) => mux_out_6_62_port, Y(61) => 
                           mux_out_6_61_port, Y(60) => mux_out_6_60_port, Y(59)
                           => mux_out_6_59_port, Y(58) => mux_out_6_58_port, 
                           Y(57) => mux_out_6_57_port, Y(56) => 
                           mux_out_6_56_port, Y(55) => mux_out_6_55_port, Y(54)
                           => mux_out_6_54_port, Y(53) => mux_out_6_53_port, 
                           Y(52) => mux_out_6_52_port, Y(51) => 
                           mux_out_6_51_port, Y(50) => mux_out_6_50_port, Y(49)
                           => mux_out_6_49_port, Y(48) => mux_out_6_48_port, 
                           Y(47) => mux_out_6_47_port, Y(46) => 
                           mux_out_6_46_port, Y(45) => mux_out_6_45_port, Y(44)
                           => mux_out_6_44_port, Y(43) => mux_out_6_43_port, 
                           Y(42) => mux_out_6_42_port, Y(41) => 
                           mux_out_6_41_port, Y(40) => mux_out_6_40_port, Y(39)
                           => mux_out_6_39_port, Y(38) => mux_out_6_38_port, 
                           Y(37) => mux_out_6_37_port, Y(36) => 
                           mux_out_6_36_port, Y(35) => mux_out_6_35_port, Y(34)
                           => mux_out_6_34_port, Y(33) => mux_out_6_33_port, 
                           Y(32) => mux_out_6_32_port, Y(31) => 
                           mux_out_6_31_port, Y(30) => mux_out_6_30_port, Y(29)
                           => mux_out_6_29_port, Y(28) => mux_out_6_28_port, 
                           Y(27) => mux_out_6_27_port, Y(26) => 
                           mux_out_6_26_port, Y(25) => mux_out_6_25_port, Y(24)
                           => mux_out_6_24_port, Y(23) => mux_out_6_23_port, 
                           Y(22) => mux_out_6_22_port, Y(21) => 
                           mux_out_6_21_port, Y(20) => mux_out_6_20_port, Y(19)
                           => mux_out_6_19_port, Y(18) => mux_out_6_18_port, 
                           Y(17) => mux_out_6_17_port, Y(16) => 
                           mux_out_6_16_port, Y(15) => mux_out_6_15_port, Y(14)
                           => mux_out_6_14_port, Y(13) => mux_out_6_13_port, 
                           Y(12) => mux_out_6_12_port, Y(11) => 
                           mux_out_6_11_port, Y(10) => mux_out_6_10_port, Y(9) 
                           => mux_out_6_9_port, Y(8) => mux_out_6_8_port, Y(7) 
                           => mux_out_6_7_port, Y(6) => mux_out_6_6_port, Y(5) 
                           => mux_out_6_5_port, Y(4) => mux_out_6_4_port, Y(3) 
                           => mux_out_6_3_port, Y(2) => mux_out_6_2_port, Y(1) 
                           => mux_out_6_1_port, Y(0) => mux_out_6_0_port);
   mux_i_7 : MUX51_GENERIC_N64_9 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n556, B(62) => n556, B(61) 
                           => n556, B(60) => n556, B(59) => n556, B(58) => n556
                           , B(57) => n556, B(56) => n555, B(55) => n555, B(54)
                           => n555, B(53) => n555, B(52) => n555, B(51) => n555
                           , B(50) => n555, B(49) => n554, B(48) => n554, B(47)
                           => n554, B(46) => n554, B(45) => n554, B(44) => n499
                           , B(43) => n489, B(42) => n479, B(41) => n469, B(40)
                           => n459, B(39) => n449, B(38) => n439, B(37) => n429
                           , B(36) => n419, B(35) => n409, B(34) => n399, B(33)
                           => n389, B(32) => n379, B(31) => n369, B(30) => n359
                           , B(29) => n349, B(28) => n339, B(27) => n329, B(26)
                           => n319, B(25) => n309, B(24) => n299, B(23) => n289
                           , B(22) => n279, B(21) => n269, B(20) => n259, B(19)
                           => n249, B(18) => n239, B(17) => n229, B(16) => n219
                           , B(15) => n209, B(14) => n199, B(13) => 
                           X_Logic0_port, B(12) => X_Logic0_port, B(11) => 
                           X_Logic0_port, B(10) => X_Logic0_port, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(63) => n643,
                           C(62) => n643, C(61) => n643, C(60) => n643, C(59) 
                           => n643, C(58) => n644, C(57) => n644, C(56) => n644
                           , C(55) => n644, C(54) => n644, C(53) => n644, C(52)
                           => n644, C(51) => n644, C(50) => n644, C(49) => n644
                           , C(48) => n644, C(47) => n644, C(46) => n645, C(45)
                           => n645, C(44) => n505, C(43) => n495, C(42) => n485
                           , C(41) => n475, C(40) => n465, C(39) => n455, C(38)
                           => n445, C(37) => n435, C(36) => n425, C(35) => n415
                           , C(34) => n405, C(33) => n395, C(32) => n385, C(31)
                           => n375, C(30) => n365, C(29) => n355, C(28) => n345
                           , C(27) => n335, C(26) => n325, C(25) => n315, C(24)
                           => n305, C(23) => n295, C(22) => n285, C(21) => n275
                           , C(20) => n265, C(19) => n255, C(18) => n245, C(17)
                           => n235, C(16) => n225, C(15) => n215, C(14) => n205
                           , C(13) => X_Logic1_port, C(12) => X_Logic1_port, 
                           C(11) => X_Logic1_port, C(10) => X_Logic1_port, C(9)
                           => X_Logic1_port, C(8) => X_Logic1_port, C(7) => 
                           X_Logic1_port, C(6) => X_Logic1_port, C(5) => 
                           X_Logic1_port, C(4) => X_Logic1_port, C(3) => 
                           X_Logic1_port, C(2) => X_Logic1_port, C(1) => 
                           X_Logic1_port, C(0) => X_Logic1_port, D(63) => n554,
                           D(62) => n554, D(61) => n553, D(60) => n553, D(59) 
                           => n553, D(58) => n553, D(57) => n553, D(56) => n553
                           , D(55) => n553, D(54) => n552, D(53) => n552, D(52)
                           => n552, D(51) => n552, D(50) => n552, D(49) => n552
                           , D(48) => n552, D(47) => n551, D(46) => n551, D(45)
                           => n499, D(44) => n489, D(43) => n479, D(42) => n469
                           , D(41) => n459, D(40) => n449, D(39) => n439, D(38)
                           => n429, D(37) => n419, D(36) => n409, D(35) => n399
                           , D(34) => n389, D(33) => n379, D(32) => n369, D(31)
                           => n359, D(30) => n349, D(29) => n339, D(28) => n329
                           , D(27) => n319, D(26) => n309, D(25) => n299, D(24)
                           => n289, D(23) => n279, D(22) => n269, D(21) => n259
                           , D(20) => n249, D(19) => n239, D(18) => n229, D(17)
                           => n219, D(16) => n209, D(15) => n199, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(63) => n680, E(62) => n680, E(61) 
                           => n668, E(60) => n668, E(59) => n668, E(58) => n668
                           , E(57) => n668, E(56) => n668, E(55) => n668, E(54)
                           => n650, E(53) => n663, E(52) => n660, E(51) => n661
                           , E(50) => n660, E(49) => n660, E(48) => n661, E(47)
                           => n660, E(46) => n660, E(45) => n507, E(44) => n497
                           , E(43) => n487, E(42) => n477, E(41) => n467, E(40)
                           => n457, E(39) => n447, E(38) => n437, E(37) => n427
                           , E(36) => n417, E(35) => n407, E(34) => n397, E(33)
                           => n387, E(32) => n377, E(31) => n367, E(30) => n357
                           , E(29) => n347, E(28) => n337, E(27) => n327, E(26)
                           => n317, E(25) => n307, E(24) => n297, E(23) => n287
                           , E(22) => n277, E(21) => n267, E(20) => n257, E(19)
                           => n247, E(18) => n237, E(17) => n227, E(16) => n217
                           , E(15) => n207, E(14) => X_Logic1_port, E(13) => 
                           X_Logic1_port, E(12) => X_Logic1_port, E(11) => 
                           X_Logic1_port, E(10) => X_Logic1_port, E(9) => 
                           X_Logic1_port, E(8) => X_Logic1_port, E(7) => 
                           X_Logic1_port, E(6) => X_Logic1_port, E(5) => 
                           X_Logic1_port, E(4) => X_Logic1_port, E(3) => 
                           X_Logic1_port, E(2) => X_Logic1_port, E(1) => 
                           X_Logic1_port, E(0) => X_Logic1_port, SEL(2) => 
                           encoder_out_23_port, SEL(1) => encoder_out_22_port, 
                           SEL(0) => encoder_out_21_port, Y(63) => 
                           mux_out_7_63_port, Y(62) => mux_out_7_62_port, Y(61)
                           => mux_out_7_61_port, Y(60) => mux_out_7_60_port, 
                           Y(59) => mux_out_7_59_port, Y(58) => 
                           mux_out_7_58_port, Y(57) => mux_out_7_57_port, Y(56)
                           => mux_out_7_56_port, Y(55) => mux_out_7_55_port, 
                           Y(54) => mux_out_7_54_port, Y(53) => 
                           mux_out_7_53_port, Y(52) => mux_out_7_52_port, Y(51)
                           => mux_out_7_51_port, Y(50) => mux_out_7_50_port, 
                           Y(49) => mux_out_7_49_port, Y(48) => 
                           mux_out_7_48_port, Y(47) => mux_out_7_47_port, Y(46)
                           => mux_out_7_46_port, Y(45) => mux_out_7_45_port, 
                           Y(44) => mux_out_7_44_port, Y(43) => 
                           mux_out_7_43_port, Y(42) => mux_out_7_42_port, Y(41)
                           => mux_out_7_41_port, Y(40) => mux_out_7_40_port, 
                           Y(39) => mux_out_7_39_port, Y(38) => 
                           mux_out_7_38_port, Y(37) => mux_out_7_37_port, Y(36)
                           => mux_out_7_36_port, Y(35) => mux_out_7_35_port, 
                           Y(34) => mux_out_7_34_port, Y(33) => 
                           mux_out_7_33_port, Y(32) => mux_out_7_32_port, Y(31)
                           => mux_out_7_31_port, Y(30) => mux_out_7_30_port, 
                           Y(29) => mux_out_7_29_port, Y(28) => 
                           mux_out_7_28_port, Y(27) => mux_out_7_27_port, Y(26)
                           => mux_out_7_26_port, Y(25) => mux_out_7_25_port, 
                           Y(24) => mux_out_7_24_port, Y(23) => 
                           mux_out_7_23_port, Y(22) => mux_out_7_22_port, Y(21)
                           => mux_out_7_21_port, Y(20) => mux_out_7_20_port, 
                           Y(19) => mux_out_7_19_port, Y(18) => 
                           mux_out_7_18_port, Y(17) => mux_out_7_17_port, Y(16)
                           => mux_out_7_16_port, Y(15) => mux_out_7_15_port, 
                           Y(14) => mux_out_7_14_port, Y(13) => 
                           mux_out_7_13_port, Y(12) => mux_out_7_12_port, Y(11)
                           => mux_out_7_11_port, Y(10) => mux_out_7_10_port, 
                           Y(9) => mux_out_7_9_port, Y(8) => mux_out_7_8_port, 
                           Y(7) => mux_out_7_7_port, Y(6) => mux_out_7_6_port, 
                           Y(5) => mux_out_7_5_port, Y(4) => mux_out_7_4_port, 
                           Y(3) => mux_out_7_3_port, Y(2) => mux_out_7_2_port, 
                           Y(1) => mux_out_7_1_port, Y(0) => mux_out_7_0_port);
   mux_i_8 : MUX51_GENERIC_N64_8 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n561, B(62) => n561, B(61) 
                           => n561, B(60) => n561, B(59) => n561, B(58) => n560
                           , B(57) => n560, B(56) => n560, B(55) => n560, B(54)
                           => n560, B(53) => n560, B(52) => n560, B(51) => n559
                           , B(50) => n559, B(49) => n559, B(48) => n559, B(47)
                           => n559, B(46) => n500, B(45) => n490, B(44) => n480
                           , B(43) => n470, B(42) => n460, B(41) => n450, B(40)
                           => n440, B(39) => n430, B(38) => n420, B(37) => n410
                           , B(36) => n400, B(35) => n390, B(34) => n380, B(33)
                           => n370, B(32) => n360, B(31) => n350, B(30) => n340
                           , B(29) => n330, B(28) => n320, B(27) => n310, B(26)
                           => n300, B(25) => n290, B(24) => n280, B(23) => n270
                           , B(22) => n260, B(21) => n250, B(20) => n240, B(19)
                           => n230, B(18) => n220, B(17) => n210, B(16) => n200
                           , B(15) => X_Logic0_port, B(14) => X_Logic0_port, 
                           B(13) => X_Logic0_port, B(12) => X_Logic0_port, 
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(63) => n645,
                           C(62) => n645, C(61) => n645, C(60) => n645, C(59) 
                           => n645, C(58) => n645, C(57) => n645, C(56) => n645
                           , C(55) => n645, C(54) => n645, C(53) => n646, C(52)
                           => n646, C(51) => n646, C(50) => n646, C(49) => n646
                           , C(48) => n646, C(47) => n646, C(46) => n506, C(45)
                           => n496, C(44) => n486, C(43) => n476, C(42) => n466
                           , C(41) => n456, C(40) => n446, C(39) => n436, C(38)
                           => n426, C(37) => n416, C(36) => n406, C(35) => n396
                           , C(34) => n386, C(33) => n376, C(32) => n366, C(31)
                           => n356, C(30) => n346, C(29) => n336, C(28) => n326
                           , C(27) => n316, C(26) => n306, C(25) => n296, C(24)
                           => n286, C(23) => n276, C(22) => n266, C(21) => n256
                           , C(20) => n246, C(19) => n236, C(18) => n226, C(17)
                           => n216, C(16) => n206, C(15) => X_Logic1_port, 
                           C(14) => X_Logic1_port, C(13) => X_Logic1_port, 
                           C(12) => X_Logic1_port, C(11) => X_Logic1_port, 
                           C(10) => X_Logic1_port, C(9) => X_Logic1_port, C(8) 
                           => X_Logic1_port, C(7) => X_Logic1_port, C(6) => 
                           X_Logic1_port, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n559, D(62) => n559, D(61) 
                           => n558, D(60) => n558, D(59) => n558, D(58) => n558
                           , D(57) => n558, D(56) => n558, D(55) => n558, D(54)
                           => n557, D(53) => n557, D(52) => n557, D(51) => n557
                           , D(50) => n557, D(49) => n557, D(48) => n557, D(47)
                           => n500, D(46) => n490, D(45) => n480, D(44) => n470
                           , D(43) => n460, D(42) => n450, D(41) => n440, D(40)
                           => n430, D(39) => n420, D(38) => n410, D(37) => n400
                           , D(36) => n390, D(35) => n380, D(34) => n370, D(33)
                           => n360, D(32) => n350, D(31) => n340, D(30) => n330
                           , D(29) => n320, D(28) => n310, D(27) => n300, D(26)
                           => n290, D(25) => n280, D(24) => n270, D(23) => n260
                           , D(22) => n250, D(21) => n240, D(20) => n230, D(19)
                           => n220, D(18) => n210, D(17) => n200, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(63) => n660, E(62) => n660, E(61) 
                           => n660, E(60) => n660, E(59) => n660, E(58) => n660
                           , E(57) => n661, E(56) => n661, E(55) => n661, E(54)
                           => n661, E(53) => n661, E(52) => n661, E(51) => n661
                           , E(50) => n661, E(49) => n661, E(48) => n662, E(47)
                           => n507, E(46) => n497, E(45) => n487, E(44) => n477
                           , E(43) => n467, E(42) => n457, E(41) => n447, E(40)
                           => n437, E(39) => n427, E(38) => n417, E(37) => n407
                           , E(36) => n397, E(35) => n387, E(34) => n377, E(33)
                           => n367, E(32) => n357, E(31) => n347, E(30) => n337
                           , E(29) => n327, E(28) => n317, E(27) => n307, E(26)
                           => n297, E(25) => n287, E(24) => n277, E(23) => n267
                           , E(22) => n257, E(21) => n247, E(20) => n237, E(19)
                           => n227, E(18) => n217, E(17) => n207, E(16) => 
                           X_Logic1_port, E(15) => X_Logic1_port, E(14) => 
                           X_Logic1_port, E(13) => X_Logic1_port, E(12) => 
                           X_Logic1_port, E(11) => X_Logic1_port, E(10) => 
                           X_Logic1_port, E(9) => X_Logic1_port, E(8) => 
                           X_Logic1_port, E(7) => X_Logic1_port, E(6) => 
                           X_Logic1_port, E(5) => X_Logic1_port, E(4) => 
                           X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_26_port, SEL(1)
                           => encoder_out_25_port, SEL(0) => 
                           encoder_out_24_port, Y(63) => mux_out_8_63_port, 
                           Y(62) => mux_out_8_62_port, Y(61) => 
                           mux_out_8_61_port, Y(60) => mux_out_8_60_port, Y(59)
                           => mux_out_8_59_port, Y(58) => mux_out_8_58_port, 
                           Y(57) => mux_out_8_57_port, Y(56) => 
                           mux_out_8_56_port, Y(55) => mux_out_8_55_port, Y(54)
                           => mux_out_8_54_port, Y(53) => mux_out_8_53_port, 
                           Y(52) => mux_out_8_52_port, Y(51) => 
                           mux_out_8_51_port, Y(50) => mux_out_8_50_port, Y(49)
                           => mux_out_8_49_port, Y(48) => mux_out_8_48_port, 
                           Y(47) => mux_out_8_47_port, Y(46) => 
                           mux_out_8_46_port, Y(45) => mux_out_8_45_port, Y(44)
                           => mux_out_8_44_port, Y(43) => mux_out_8_43_port, 
                           Y(42) => mux_out_8_42_port, Y(41) => 
                           mux_out_8_41_port, Y(40) => mux_out_8_40_port, Y(39)
                           => mux_out_8_39_port, Y(38) => mux_out_8_38_port, 
                           Y(37) => mux_out_8_37_port, Y(36) => 
                           mux_out_8_36_port, Y(35) => mux_out_8_35_port, Y(34)
                           => mux_out_8_34_port, Y(33) => mux_out_8_33_port, 
                           Y(32) => mux_out_8_32_port, Y(31) => 
                           mux_out_8_31_port, Y(30) => mux_out_8_30_port, Y(29)
                           => mux_out_8_29_port, Y(28) => mux_out_8_28_port, 
                           Y(27) => mux_out_8_27_port, Y(26) => 
                           mux_out_8_26_port, Y(25) => mux_out_8_25_port, Y(24)
                           => mux_out_8_24_port, Y(23) => mux_out_8_23_port, 
                           Y(22) => mux_out_8_22_port, Y(21) => 
                           mux_out_8_21_port, Y(20) => mux_out_8_20_port, Y(19)
                           => mux_out_8_19_port, Y(18) => mux_out_8_18_port, 
                           Y(17) => mux_out_8_17_port, Y(16) => 
                           mux_out_8_16_port, Y(15) => mux_out_8_15_port, Y(14)
                           => mux_out_8_14_port, Y(13) => mux_out_8_13_port, 
                           Y(12) => mux_out_8_12_port, Y(11) => 
                           mux_out_8_11_port, Y(10) => mux_out_8_10_port, Y(9) 
                           => mux_out_8_9_port, Y(8) => mux_out_8_8_port, Y(7) 
                           => mux_out_8_7_port, Y(6) => mux_out_8_6_port, Y(5) 
                           => mux_out_8_5_port, Y(4) => mux_out_8_4_port, Y(3) 
                           => mux_out_8_3_port, Y(2) => mux_out_8_2_port, Y(1) 
                           => mux_out_8_1_port, Y(0) => mux_out_8_0_port);
   mux_i_9 : MUX51_GENERIC_N64_7 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n565, B(62) => n565, B(61) 
                           => n565, B(60) => n565, B(59) => n565, B(58) => n565
                           , B(57) => n564, B(56) => n564, B(55) => n564, B(54)
                           => n564, B(53) => n564, B(52) => n564, B(51) => n564
                           , B(50) => n563, B(49) => n563, B(48) => n500, B(47)
                           => n490, B(46) => n480, B(45) => n470, B(44) => n460
                           , B(43) => n450, B(42) => n440, B(41) => n430, B(40)
                           => n420, B(39) => n410, B(38) => n400, B(37) => n390
                           , B(36) => n380, B(35) => n370, B(34) => n360, B(33)
                           => n350, B(32) => n340, B(31) => n330, B(30) => n320
                           , B(29) => n310, B(28) => n300, B(27) => n290, B(26)
                           => n280, B(25) => n270, B(24) => n260, B(23) => n250
                           , B(22) => n240, B(21) => n230, B(20) => n220, B(19)
                           => n210, B(18) => n200, B(17) => X_Logic0_port, 
                           B(16) => X_Logic0_port, B(15) => X_Logic0_port, 
                           B(14) => X_Logic0_port, B(13) => X_Logic0_port, 
                           B(12) => X_Logic0_port, B(11) => X_Logic0_port, 
                           B(10) => X_Logic0_port, B(9) => X_Logic0_port, B(8) 
                           => X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, C(63) => n646, C(62) => n646, C(61) 
                           => n646, C(60) => n646, C(59) => n646, C(58) => n647
                           , C(57) => n647, C(56) => n647, C(55) => n647, C(54)
                           => n647, C(53) => n647, C(52) => n647, C(51) => n647
                           , C(50) => n647, C(49) => n647, C(48) => n506, C(47)
                           => n496, C(46) => n486, C(45) => n476, C(44) => n466
                           , C(43) => n456, C(42) => n446, C(41) => n436, C(40)
                           => n426, C(39) => n416, C(38) => n406, C(37) => n396
                           , C(36) => n386, C(35) => n376, C(34) => n366, C(33)
                           => n356, C(32) => n346, C(31) => n336, C(30) => n326
                           , C(29) => n316, C(28) => n306, C(27) => n296, C(26)
                           => n286, C(25) => n276, C(24) => n266, C(23) => n256
                           , C(22) => n246, C(21) => n236, C(20) => n226, C(19)
                           => n216, C(18) => n206, C(17) => X_Logic1_port, 
                           C(16) => X_Logic1_port, C(15) => X_Logic1_port, 
                           C(14) => X_Logic1_port, C(13) => X_Logic1_port, 
                           C(12) => X_Logic1_port, C(11) => X_Logic1_port, 
                           C(10) => X_Logic1_port, C(9) => X_Logic1_port, C(8) 
                           => X_Logic1_port, C(7) => X_Logic1_port, C(6) => 
                           X_Logic1_port, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n563, D(62) => n563, D(61) 
                           => n563, D(60) => n563, D(59) => n563, D(58) => n562
                           , D(57) => n562, D(56) => n562, D(55) => n562, D(54)
                           => n562, D(53) => n562, D(52) => n562, D(51) => n561
                           , D(50) => n561, D(49) => n500, D(48) => n490, D(47)
                           => n480, D(46) => n470, D(45) => n460, D(44) => n450
                           , D(43) => n440, D(42) => n430, D(41) => n420, D(40)
                           => n410, D(39) => n400, D(38) => n390, D(37) => n380
                           , D(36) => n370, D(35) => n360, D(34) => n350, D(33)
                           => n340, D(32) => n330, D(31) => n320, D(30) => n310
                           , D(29) => n300, D(28) => n290, D(27) => n280, D(26)
                           => n270, D(25) => n260, D(24) => n250, D(23) => n240
                           , D(22) => n230, D(21) => n220, D(20) => n210, D(19)
                           => n200, D(18) => X_Logic0_port, D(17) => 
                           X_Logic0_port, D(16) => X_Logic0_port, D(15) => 
                           X_Logic0_port, D(14) => X_Logic0_port, D(13) => 
                           X_Logic0_port, D(12) => X_Logic0_port, D(11) => 
                           X_Logic0_port, D(10) => X_Logic0_port, D(9) => 
                           X_Logic0_port, D(8) => X_Logic0_port, D(7) => 
                           X_Logic0_port, D(6) => X_Logic0_port, D(5) => 
                           X_Logic0_port, D(4) => X_Logic0_port, D(3) => 
                           X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, E(63) => n663,
                           E(62) => n663, E(61) => n663, E(60) => n663, E(59) 
                           => n663, E(58) => n663, E(57) => n663, E(56) => n664
                           , E(55) => n664, E(54) => n664, E(53) => n664, E(52)
                           => n664, E(51) => n664, E(50) => n664, E(49) => n506
                           , E(48) => n496, E(47) => n486, E(46) => n476, E(45)
                           => n466, E(44) => n456, E(43) => n446, E(42) => n436
                           , E(41) => n426, E(40) => n416, E(39) => n406, E(38)
                           => n396, E(37) => n386, E(36) => n376, E(35) => n366
                           , E(34) => n356, E(33) => n346, E(32) => n336, E(31)
                           => n326, E(30) => n316, E(29) => n306, E(28) => n296
                           , E(27) => n286, E(26) => n276, E(25) => n266, E(24)
                           => n256, E(23) => n246, E(22) => n236, E(21) => n226
                           , E(20) => n216, E(19) => n206, E(18) => 
                           X_Logic1_port, E(17) => X_Logic1_port, E(16) => 
                           X_Logic1_port, E(15) => X_Logic1_port, E(14) => 
                           X_Logic1_port, E(13) => X_Logic1_port, E(12) => 
                           X_Logic1_port, E(11) => X_Logic1_port, E(10) => 
                           X_Logic1_port, E(9) => X_Logic1_port, E(8) => 
                           X_Logic1_port, E(7) => X_Logic1_port, E(6) => 
                           X_Logic1_port, E(5) => X_Logic1_port, E(4) => 
                           X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_29_port, SEL(1)
                           => encoder_out_28_port, SEL(0) => 
                           encoder_out_27_port, Y(63) => mux_out_9_63_port, 
                           Y(62) => mux_out_9_62_port, Y(61) => 
                           mux_out_9_61_port, Y(60) => mux_out_9_60_port, Y(59)
                           => mux_out_9_59_port, Y(58) => mux_out_9_58_port, 
                           Y(57) => mux_out_9_57_port, Y(56) => 
                           mux_out_9_56_port, Y(55) => mux_out_9_55_port, Y(54)
                           => mux_out_9_54_port, Y(53) => mux_out_9_53_port, 
                           Y(52) => mux_out_9_52_port, Y(51) => 
                           mux_out_9_51_port, Y(50) => mux_out_9_50_port, Y(49)
                           => mux_out_9_49_port, Y(48) => mux_out_9_48_port, 
                           Y(47) => mux_out_9_47_port, Y(46) => 
                           mux_out_9_46_port, Y(45) => mux_out_9_45_port, Y(44)
                           => mux_out_9_44_port, Y(43) => mux_out_9_43_port, 
                           Y(42) => mux_out_9_42_port, Y(41) => 
                           mux_out_9_41_port, Y(40) => mux_out_9_40_port, Y(39)
                           => mux_out_9_39_port, Y(38) => mux_out_9_38_port, 
                           Y(37) => mux_out_9_37_port, Y(36) => 
                           mux_out_9_36_port, Y(35) => mux_out_9_35_port, Y(34)
                           => mux_out_9_34_port, Y(33) => mux_out_9_33_port, 
                           Y(32) => mux_out_9_32_port, Y(31) => 
                           mux_out_9_31_port, Y(30) => mux_out_9_30_port, Y(29)
                           => mux_out_9_29_port, Y(28) => mux_out_9_28_port, 
                           Y(27) => mux_out_9_27_port, Y(26) => 
                           mux_out_9_26_port, Y(25) => mux_out_9_25_port, Y(24)
                           => mux_out_9_24_port, Y(23) => mux_out_9_23_port, 
                           Y(22) => mux_out_9_22_port, Y(21) => 
                           mux_out_9_21_port, Y(20) => mux_out_9_20_port, Y(19)
                           => mux_out_9_19_port, Y(18) => mux_out_9_18_port, 
                           Y(17) => mux_out_9_17_port, Y(16) => 
                           mux_out_9_16_port, Y(15) => mux_out_9_15_port, Y(14)
                           => mux_out_9_14_port, Y(13) => mux_out_9_13_port, 
                           Y(12) => mux_out_9_12_port, Y(11) => 
                           mux_out_9_11_port, Y(10) => mux_out_9_10_port, Y(9) 
                           => mux_out_9_9_port, Y(8) => mux_out_9_8_port, Y(7) 
                           => mux_out_9_7_port, Y(6) => mux_out_9_6_port, Y(5) 
                           => mux_out_9_5_port, Y(4) => mux_out_9_4_port, Y(3) 
                           => mux_out_9_3_port, Y(2) => mux_out_9_2_port, Y(1) 
                           => mux_out_9_1_port, Y(0) => mux_out_9_0_port);
   mux_i_10 : MUX51_GENERIC_N64_6 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n569, B(62) => n569, B(61) 
                           => n569, B(60) => n568, B(59) => n568, B(58) => n568
                           , B(57) => n568, B(56) => n568, B(55) => n568, B(54)
                           => n568, B(53) => n567, B(52) => n567, B(51) => n567
                           , B(50) => n500, B(49) => n490, B(48) => n480, B(47)
                           => n470, B(46) => n460, B(45) => n450, B(44) => n440
                           , B(43) => n430, B(42) => n420, B(41) => n410, B(40)
                           => n400, B(39) => n390, B(38) => n380, B(37) => n370
                           , B(36) => n360, B(35) => n350, B(34) => n340, B(33)
                           => n330, B(32) => n320, B(31) => n310, B(30) => n300
                           , B(29) => n290, B(28) => n280, B(27) => n270, B(26)
                           => n260, B(25) => n250, B(24) => n240, B(23) => n230
                           , B(22) => n220, B(21) => n210, B(20) => n200, B(19)
                           => X_Logic0_port, B(18) => X_Logic0_port, B(17) => 
                           X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
                           X_Logic0_port, B(14) => X_Logic0_port, B(13) => 
                           X_Logic0_port, B(12) => X_Logic0_port, B(11) => 
                           X_Logic0_port, B(10) => X_Logic0_port, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(63) => n647,
                           C(62) => n647, C(61) => n648, C(60) => n648, C(59) 
                           => n648, C(58) => n648, C(57) => n648, C(56) => n648
                           , C(55) => n648, C(54) => n648, C(53) => n648, C(52)
                           => n648, C(51) => n648, C(50) => n506, C(49) => n496
                           , C(48) => n486, C(47) => n476, C(46) => n466, C(45)
                           => n456, C(44) => n446, C(43) => n436, C(42) => n426
                           , C(41) => n416, C(40) => n406, C(39) => n396, C(38)
                           => n386, C(37) => n376, C(36) => n366, C(35) => n356
                           , C(34) => n346, C(33) => n336, C(32) => n326, C(31)
                           => n316, C(30) => n306, C(29) => n296, C(28) => n286
                           , C(27) => n276, C(26) => n266, C(25) => n256, C(24)
                           => n246, C(23) => n236, C(22) => n226, C(21) => n216
                           , C(20) => n206, C(19) => X_Logic1_port, C(18) => 
                           X_Logic1_port, C(17) => X_Logic1_port, C(16) => 
                           X_Logic1_port, C(15) => X_Logic1_port, C(14) => 
                           X_Logic1_port, C(13) => X_Logic1_port, C(12) => 
                           X_Logic1_port, C(11) => X_Logic1_port, C(10) => 
                           X_Logic1_port, C(9) => X_Logic1_port, C(8) => 
                           X_Logic1_port, C(7) => X_Logic1_port, C(6) => 
                           X_Logic1_port, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n567, D(62) => n567, D(61) 
                           => n567, D(60) => n567, D(59) => n566, D(58) => n566
                           , D(57) => n566, D(56) => n566, D(55) => n566, D(54)
                           => n566, D(53) => n566, D(52) => n565, D(51) => n500
                           , D(50) => n490, D(49) => n480, D(48) => n470, D(47)
                           => n460, D(46) => n450, D(45) => n440, D(44) => n430
                           , D(43) => n420, D(42) => n410, D(41) => n400, D(40)
                           => n390, D(39) => n380, D(38) => n370, D(37) => n360
                           , D(36) => n350, D(35) => n340, D(34) => n330, D(33)
                           => n320, D(32) => n310, D(31) => n300, D(30) => n290
                           , D(29) => n280, D(28) => n270, D(27) => n260, D(26)
                           => n250, D(25) => n240, D(24) => n230, D(23) => n220
                           , D(22) => n210, D(21) => n200, D(20) => 
                           X_Logic0_port, D(19) => X_Logic0_port, D(18) => 
                           X_Logic0_port, D(17) => X_Logic0_port, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(63) => n665, E(62) => n665, E(61) 
                           => n665, E(60) => n665, E(59) => n666, E(58) => n666
                           , E(57) => n666, E(56) => n666, E(55) => n666, E(54)
                           => n666, E(53) => n666, E(52) => n666, E(51) => n506
                           , E(50) => n496, E(49) => n486, E(48) => n476, E(47)
                           => n466, E(46) => n456, E(45) => n446, E(44) => n436
                           , E(43) => n426, E(42) => n416, E(41) => n406, E(40)
                           => n396, E(39) => n386, E(38) => n376, E(37) => n366
                           , E(36) => n356, E(35) => n346, E(34) => n336, E(33)
                           => n326, E(32) => n316, E(31) => n306, E(30) => n296
                           , E(29) => n286, E(28) => n276, E(27) => n266, E(26)
                           => n256, E(25) => n246, E(24) => n236, E(23) => n226
                           , E(22) => n216, E(21) => n206, E(20) => 
                           X_Logic1_port, E(19) => X_Logic1_port, E(18) => 
                           X_Logic1_port, E(17) => X_Logic1_port, E(16) => 
                           X_Logic1_port, E(15) => X_Logic1_port, E(14) => 
                           X_Logic1_port, E(13) => X_Logic1_port, E(12) => 
                           X_Logic1_port, E(11) => X_Logic1_port, E(10) => 
                           X_Logic1_port, E(9) => X_Logic1_port, E(8) => 
                           X_Logic1_port, E(7) => X_Logic1_port, E(6) => 
                           X_Logic1_port, E(5) => X_Logic1_port, E(4) => 
                           X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_32_port, SEL(1)
                           => encoder_out_31_port, SEL(0) => 
                           encoder_out_30_port, Y(63) => mux_out_10_63_port, 
                           Y(62) => mux_out_10_62_port, Y(61) => 
                           mux_out_10_61_port, Y(60) => mux_out_10_60_port, 
                           Y(59) => mux_out_10_59_port, Y(58) => 
                           mux_out_10_58_port, Y(57) => mux_out_10_57_port, 
                           Y(56) => mux_out_10_56_port, Y(55) => 
                           mux_out_10_55_port, Y(54) => mux_out_10_54_port, 
                           Y(53) => mux_out_10_53_port, Y(52) => 
                           mux_out_10_52_port, Y(51) => mux_out_10_51_port, 
                           Y(50) => mux_out_10_50_port, Y(49) => 
                           mux_out_10_49_port, Y(48) => mux_out_10_48_port, 
                           Y(47) => mux_out_10_47_port, Y(46) => 
                           mux_out_10_46_port, Y(45) => mux_out_10_45_port, 
                           Y(44) => mux_out_10_44_port, Y(43) => 
                           mux_out_10_43_port, Y(42) => mux_out_10_42_port, 
                           Y(41) => mux_out_10_41_port, Y(40) => 
                           mux_out_10_40_port, Y(39) => mux_out_10_39_port, 
                           Y(38) => mux_out_10_38_port, Y(37) => 
                           mux_out_10_37_port, Y(36) => mux_out_10_36_port, 
                           Y(35) => mux_out_10_35_port, Y(34) => 
                           mux_out_10_34_port, Y(33) => mux_out_10_33_port, 
                           Y(32) => mux_out_10_32_port, Y(31) => 
                           mux_out_10_31_port, Y(30) => mux_out_10_30_port, 
                           Y(29) => mux_out_10_29_port, Y(28) => 
                           mux_out_10_28_port, Y(27) => mux_out_10_27_port, 
                           Y(26) => mux_out_10_26_port, Y(25) => 
                           mux_out_10_25_port, Y(24) => mux_out_10_24_port, 
                           Y(23) => mux_out_10_23_port, Y(22) => 
                           mux_out_10_22_port, Y(21) => mux_out_10_21_port, 
                           Y(20) => mux_out_10_20_port, Y(19) => 
                           mux_out_10_19_port, Y(18) => mux_out_10_18_port, 
                           Y(17) => mux_out_10_17_port, Y(16) => 
                           mux_out_10_16_port, Y(15) => mux_out_10_15_port, 
                           Y(14) => mux_out_10_14_port, Y(13) => 
                           mux_out_10_13_port, Y(12) => mux_out_10_12_port, 
                           Y(11) => mux_out_10_11_port, Y(10) => 
                           mux_out_10_10_port, Y(9) => mux_out_10_9_port, Y(8) 
                           => mux_out_10_8_port, Y(7) => mux_out_10_7_port, 
                           Y(6) => mux_out_10_6_port, Y(5) => mux_out_10_5_port
                           , Y(4) => mux_out_10_4_port, Y(3) => 
                           mux_out_10_3_port, Y(2) => mux_out_10_2_port, Y(1) 
                           => mux_out_10_1_port, Y(0) => mux_out_10_0_port);
   mux_i_11 : MUX51_GENERIC_N64_5 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n572, B(62) => n572, B(61) 
                           => n572, B(60) => n571, B(59) => n571, B(58) => n571
                           , B(57) => n571, B(56) => n571, B(55) => n571, B(54)
                           => n571, B(53) => n570, B(52) => n501, B(51) => n491
                           , B(50) => n481, B(49) => n471, B(48) => n461, B(47)
                           => n451, B(46) => n441, B(45) => n431, B(44) => n421
                           , B(43) => n411, B(42) => n401, B(41) => n391, B(40)
                           => n381, B(39) => n371, B(38) => n361, B(37) => n351
                           , B(36) => n341, B(35) => n331, B(34) => n321, B(33)
                           => n311, B(32) => n301, B(31) => n291, B(30) => n281
                           , B(29) => n271, B(28) => n261, B(27) => n251, B(26)
                           => n241, B(25) => n231, B(24) => n221, B(23) => n211
                           , B(22) => n201, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, C(63) => n648, C(62) => n649, C(61) 
                           => n649, C(60) => n649, C(59) => n649, C(58) => n649
                           , C(57) => n649, C(56) => n649, C(55) => n649, C(54)
                           => n649, C(53) => n649, C(52) => n506, C(51) => n496
                           , C(50) => n486, C(49) => n476, C(48) => n466, C(47)
                           => n456, C(46) => n446, C(45) => n436, C(44) => n426
                           , C(43) => n416, C(42) => n406, C(41) => n396, C(40)
                           => n386, C(39) => n376, C(38) => n366, C(37) => n356
                           , C(36) => n346, C(35) => n336, C(34) => n326, C(33)
                           => n316, C(32) => n306, C(31) => n296, C(30) => n286
                           , C(29) => n276, C(28) => n266, C(27) => n256, C(26)
                           => n246, C(25) => n236, C(24) => n226, C(23) => n216
                           , C(22) => n206, C(21) => X_Logic1_port, C(20) => 
                           X_Logic1_port, C(19) => X_Logic1_port, C(18) => 
                           X_Logic1_port, C(17) => X_Logic1_port, C(16) => 
                           X_Logic1_port, C(15) => X_Logic1_port, C(14) => 
                           X_Logic1_port, C(13) => X_Logic1_port, C(12) => 
                           X_Logic1_port, C(11) => X_Logic1_port, C(10) => 
                           X_Logic1_port, C(9) => X_Logic1_port, C(8) => 
                           X_Logic1_port, C(7) => X_Logic1_port, C(6) => 
                           X_Logic1_port, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n570, D(62) => n570, D(61) 
                           => n570, D(60) => n570, D(59) => n570, D(58) => n570
                           , D(57) => n569, D(56) => n569, D(55) => n569, D(54)
                           => n569, D(53) => n500, D(52) => n490, D(51) => n480
                           , D(50) => n470, D(49) => n460, D(48) => n450, D(47)
                           => n440, D(46) => n430, D(45) => n420, D(44) => n410
                           , D(43) => n400, D(42) => n390, D(41) => n380, D(40)
                           => n370, D(39) => n360, D(38) => n350, D(37) => n340
                           , D(36) => n330, D(35) => n320, D(34) => n310, D(33)
                           => n300, D(32) => n290, D(31) => n280, D(30) => n270
                           , D(29) => n260, D(28) => n250, D(27) => n240, D(26)
                           => n230, D(25) => n220, D(24) => n210, D(23) => n200
                           , D(22) => X_Logic0_port, D(21) => X_Logic0_port, 
                           D(20) => X_Logic0_port, D(19) => X_Logic0_port, 
                           D(18) => X_Logic0_port, D(17) => X_Logic0_port, 
                           D(16) => X_Logic0_port, D(15) => X_Logic0_port, 
                           D(14) => X_Logic0_port, D(13) => X_Logic0_port, 
                           D(12) => X_Logic0_port, D(11) => X_Logic0_port, 
                           D(10) => X_Logic0_port, D(9) => X_Logic0_port, D(8) 
                           => X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(63) => n666, E(62) => n667, E(61) 
                           => n667, E(60) => n667, E(59) => n667, E(58) => n667
                           , E(57) => n667, E(56) => n667, E(55) => n667, E(54)
                           => n667, E(53) => n506, E(52) => n496, E(51) => n486
                           , E(50) => n476, E(49) => n466, E(48) => n456, E(47)
                           => n446, E(46) => n436, E(45) => n426, E(44) => n416
                           , E(43) => n406, E(42) => n396, E(41) => n386, E(40)
                           => n376, E(39) => n366, E(38) => n356, E(37) => n346
                           , E(36) => n336, E(35) => n326, E(34) => n316, E(33)
                           => n306, E(32) => n296, E(31) => n286, E(30) => n276
                           , E(29) => n266, E(28) => n256, E(27) => n246, E(26)
                           => n236, E(25) => n226, E(24) => n216, E(23) => n206
                           , E(22) => X_Logic1_port, E(21) => X_Logic1_port, 
                           E(20) => X_Logic1_port, E(19) => X_Logic1_port, 
                           E(18) => X_Logic1_port, E(17) => X_Logic1_port, 
                           E(16) => X_Logic1_port, E(15) => X_Logic1_port, 
                           E(14) => X_Logic1_port, E(13) => X_Logic1_port, 
                           E(12) => X_Logic1_port, E(11) => X_Logic1_port, 
                           E(10) => X_Logic1_port, E(9) => X_Logic1_port, E(8) 
                           => X_Logic1_port, E(7) => X_Logic1_port, E(6) => 
                           X_Logic1_port, E(5) => X_Logic1_port, E(4) => 
                           X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_35_port, SEL(1)
                           => encoder_out_34_port, SEL(0) => 
                           encoder_out_33_port, Y(63) => mux_out_11_63_port, 
                           Y(62) => mux_out_11_62_port, Y(61) => 
                           mux_out_11_61_port, Y(60) => mux_out_11_60_port, 
                           Y(59) => mux_out_11_59_port, Y(58) => 
                           mux_out_11_58_port, Y(57) => mux_out_11_57_port, 
                           Y(56) => mux_out_11_56_port, Y(55) => 
                           mux_out_11_55_port, Y(54) => mux_out_11_54_port, 
                           Y(53) => mux_out_11_53_port, Y(52) => 
                           mux_out_11_52_port, Y(51) => mux_out_11_51_port, 
                           Y(50) => mux_out_11_50_port, Y(49) => 
                           mux_out_11_49_port, Y(48) => mux_out_11_48_port, 
                           Y(47) => mux_out_11_47_port, Y(46) => 
                           mux_out_11_46_port, Y(45) => mux_out_11_45_port, 
                           Y(44) => mux_out_11_44_port, Y(43) => 
                           mux_out_11_43_port, Y(42) => mux_out_11_42_port, 
                           Y(41) => mux_out_11_41_port, Y(40) => 
                           mux_out_11_40_port, Y(39) => mux_out_11_39_port, 
                           Y(38) => mux_out_11_38_port, Y(37) => 
                           mux_out_11_37_port, Y(36) => mux_out_11_36_port, 
                           Y(35) => mux_out_11_35_port, Y(34) => 
                           mux_out_11_34_port, Y(33) => mux_out_11_33_port, 
                           Y(32) => mux_out_11_32_port, Y(31) => 
                           mux_out_11_31_port, Y(30) => mux_out_11_30_port, 
                           Y(29) => mux_out_11_29_port, Y(28) => 
                           mux_out_11_28_port, Y(27) => mux_out_11_27_port, 
                           Y(26) => mux_out_11_26_port, Y(25) => 
                           mux_out_11_25_port, Y(24) => mux_out_11_24_port, 
                           Y(23) => mux_out_11_23_port, Y(22) => 
                           mux_out_11_22_port, Y(21) => mux_out_11_21_port, 
                           Y(20) => mux_out_11_20_port, Y(19) => 
                           mux_out_11_19_port, Y(18) => mux_out_11_18_port, 
                           Y(17) => mux_out_11_17_port, Y(16) => 
                           mux_out_11_16_port, Y(15) => mux_out_11_15_port, 
                           Y(14) => mux_out_11_14_port, Y(13) => 
                           mux_out_11_13_port, Y(12) => mux_out_11_12_port, 
                           Y(11) => mux_out_11_11_port, Y(10) => 
                           mux_out_11_10_port, Y(9) => mux_out_11_9_port, Y(8) 
                           => mux_out_11_8_port, Y(7) => mux_out_11_7_port, 
                           Y(6) => mux_out_11_6_port, Y(5) => mux_out_11_5_port
                           , Y(4) => mux_out_11_4_port, Y(3) => 
                           mux_out_11_3_port, Y(2) => mux_out_11_2_port, Y(1) 
                           => mux_out_11_1_port, Y(0) => mux_out_11_0_port);
   mux_i_12 : MUX51_GENERIC_N64_4 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n574, B(62) => n574, B(61) 
                           => n574, B(60) => n574, B(59) => n574, B(58) => n574
                           , B(57) => n573, B(56) => n573, B(55) => n573, B(54)
                           => n501, B(53) => n491, B(52) => n481, B(51) => n471
                           , B(50) => n461, B(49) => n451, B(48) => n441, B(47)
                           => n431, B(46) => n421, B(45) => n411, B(44) => n401
                           , B(43) => n391, B(42) => n381, B(41) => n371, B(40)
                           => n361, B(39) => n351, B(38) => n341, B(37) => n331
                           , B(36) => n321, B(35) => n311, B(34) => n301, B(33)
                           => n291, B(32) => n281, B(31) => n271, B(30) => n261
                           , B(29) => n251, B(28) => n241, B(27) => n231, B(26)
                           => n221, B(25) => n211, B(24) => n201, B(23) => 
                           X_Logic0_port, B(22) => X_Logic0_port, B(21) => 
                           X_Logic0_port, B(20) => X_Logic0_port, B(19) => 
                           X_Logic0_port, B(18) => X_Logic0_port, B(17) => 
                           X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
                           X_Logic0_port, B(14) => X_Logic0_port, B(13) => 
                           X_Logic0_port, B(12) => X_Logic0_port, B(11) => 
                           X_Logic0_port, B(10) => X_Logic0_port, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(63) => n649,
                           C(62) => n649, C(61) => n650, C(60) => n650, C(59) 
                           => n650, C(58) => n650, C(57) => n650, C(56) => n650
                           , C(55) => n650, C(54) => n505, C(53) => n495, C(52)
                           => n485, C(51) => n475, C(50) => n465, C(49) => n455
                           , C(48) => n445, C(47) => n435, C(46) => n425, C(45)
                           => n415, C(44) => n405, C(43) => n395, C(42) => n385
                           , C(41) => n375, C(40) => n365, C(39) => n355, C(38)
                           => n345, C(37) => n335, C(36) => n325, C(35) => n315
                           , C(34) => n305, C(33) => n295, C(32) => n285, C(31)
                           => n275, C(30) => n265, C(29) => n255, C(28) => n245
                           , C(27) => n235, C(26) => n225, C(25) => n215, C(24)
                           => n205, C(23) => X_Logic1_port, C(22) => 
                           X_Logic1_port, C(21) => X_Logic1_port, C(20) => 
                           X_Logic1_port, C(19) => X_Logic1_port, C(18) => 
                           X_Logic1_port, C(17) => X_Logic1_port, C(16) => 
                           X_Logic1_port, C(15) => X_Logic1_port, C(14) => 
                           X_Logic1_port, C(13) => X_Logic1_port, C(12) => 
                           X_Logic1_port, C(11) => X_Logic1_port, C(10) => 
                           X_Logic1_port, C(9) => X_Logic1_port, C(8) => 
                           X_Logic1_port, C(7) => X_Logic1_port, C(6) => 
                           X_Logic1_port, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n573, D(62) => n573, D(61) 
                           => n573, D(60) => n573, D(59) => n572, D(58) => n572
                           , D(57) => n572, D(56) => n572, D(55) => n501, D(54)
                           => n491, D(53) => n481, D(52) => n471, D(51) => n461
                           , D(50) => n451, D(49) => n441, D(48) => n431, D(47)
                           => n421, D(46) => n411, D(45) => n401, D(44) => n391
                           , D(43) => n381, D(42) => n371, D(41) => n361, D(40)
                           => n351, D(39) => n341, D(38) => n331, D(37) => n321
                           , D(36) => n311, D(35) => n301, D(34) => n291, D(33)
                           => n281, D(32) => n271, D(31) => n261, D(30) => n251
                           , D(29) => n241, D(28) => n231, D(27) => n221, D(26)
                           => n211, D(25) => n201, D(24) => X_Logic0_port, 
                           D(23) => X_Logic0_port, D(22) => X_Logic0_port, 
                           D(21) => X_Logic0_port, D(20) => X_Logic0_port, 
                           D(19) => X_Logic0_port, D(18) => X_Logic0_port, 
                           D(17) => X_Logic0_port, D(16) => X_Logic0_port, 
                           D(15) => X_Logic0_port, D(14) => X_Logic0_port, 
                           D(13) => X_Logic0_port, D(12) => X_Logic0_port, 
                           D(11) => X_Logic0_port, D(10) => X_Logic0_port, D(9)
                           => X_Logic0_port, D(8) => X_Logic0_port, D(7) => 
                           X_Logic0_port, D(6) => X_Logic0_port, D(5) => 
                           X_Logic0_port, D(4) => X_Logic0_port, D(3) => 
                           X_Logic0_port, D(2) => X_Logic0_port, D(1) => 
                           X_Logic0_port, D(0) => X_Logic0_port, E(63) => n667,
                           E(62) => n667, E(61) => n667, E(60) => n668, E(59) 
                           => n668, E(58) => n668, E(57) => n668, E(56) => n668
                           , E(55) => n506, E(54) => n496, E(53) => n486, E(52)
                           => n476, E(51) => n466, E(50) => n456, E(49) => n446
                           , E(48) => n436, E(47) => n426, E(46) => n416, E(45)
                           => n406, E(44) => n396, E(43) => n386, E(42) => n376
                           , E(41) => n366, E(40) => n356, E(39) => n346, E(38)
                           => n336, E(37) => n326, E(36) => n316, E(35) => n306
                           , E(34) => n296, E(33) => n286, E(32) => n276, E(31)
                           => n266, E(30) => n256, E(29) => n246, E(28) => n236
                           , E(27) => n226, E(26) => n216, E(25) => n206, E(24)
                           => X_Logic1_port, E(23) => X_Logic1_port, E(22) => 
                           X_Logic1_port, E(21) => X_Logic1_port, E(20) => 
                           X_Logic1_port, E(19) => X_Logic1_port, E(18) => 
                           X_Logic1_port, E(17) => X_Logic1_port, E(16) => 
                           X_Logic1_port, E(15) => X_Logic1_port, E(14) => 
                           X_Logic1_port, E(13) => X_Logic1_port, E(12) => 
                           X_Logic1_port, E(11) => X_Logic1_port, E(10) => 
                           X_Logic1_port, E(9) => X_Logic1_port, E(8) => 
                           X_Logic1_port, E(7) => X_Logic1_port, E(6) => 
                           X_Logic1_port, E(5) => X_Logic1_port, E(4) => 
                           X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_38_port, SEL(1)
                           => encoder_out_37_port, SEL(0) => 
                           encoder_out_36_port, Y(63) => mux_out_12_63_port, 
                           Y(62) => mux_out_12_62_port, Y(61) => 
                           mux_out_12_61_port, Y(60) => mux_out_12_60_port, 
                           Y(59) => mux_out_12_59_port, Y(58) => 
                           mux_out_12_58_port, Y(57) => mux_out_12_57_port, 
                           Y(56) => mux_out_12_56_port, Y(55) => 
                           mux_out_12_55_port, Y(54) => mux_out_12_54_port, 
                           Y(53) => mux_out_12_53_port, Y(52) => 
                           mux_out_12_52_port, Y(51) => mux_out_12_51_port, 
                           Y(50) => mux_out_12_50_port, Y(49) => 
                           mux_out_12_49_port, Y(48) => mux_out_12_48_port, 
                           Y(47) => mux_out_12_47_port, Y(46) => 
                           mux_out_12_46_port, Y(45) => mux_out_12_45_port, 
                           Y(44) => mux_out_12_44_port, Y(43) => 
                           mux_out_12_43_port, Y(42) => mux_out_12_42_port, 
                           Y(41) => mux_out_12_41_port, Y(40) => 
                           mux_out_12_40_port, Y(39) => mux_out_12_39_port, 
                           Y(38) => mux_out_12_38_port, Y(37) => 
                           mux_out_12_37_port, Y(36) => mux_out_12_36_port, 
                           Y(35) => mux_out_12_35_port, Y(34) => 
                           mux_out_12_34_port, Y(33) => mux_out_12_33_port, 
                           Y(32) => mux_out_12_32_port, Y(31) => 
                           mux_out_12_31_port, Y(30) => mux_out_12_30_port, 
                           Y(29) => mux_out_12_29_port, Y(28) => 
                           mux_out_12_28_port, Y(27) => mux_out_12_27_port, 
                           Y(26) => mux_out_12_26_port, Y(25) => 
                           mux_out_12_25_port, Y(24) => mux_out_12_24_port, 
                           Y(23) => mux_out_12_23_port, Y(22) => 
                           mux_out_12_22_port, Y(21) => mux_out_12_21_port, 
                           Y(20) => mux_out_12_20_port, Y(19) => 
                           mux_out_12_19_port, Y(18) => mux_out_12_18_port, 
                           Y(17) => mux_out_12_17_port, Y(16) => 
                           mux_out_12_16_port, Y(15) => mux_out_12_15_port, 
                           Y(14) => mux_out_12_14_port, Y(13) => 
                           mux_out_12_13_port, Y(12) => mux_out_12_12_port, 
                           Y(11) => mux_out_12_11_port, Y(10) => 
                           mux_out_12_10_port, Y(9) => mux_out_12_9_port, Y(8) 
                           => mux_out_12_8_port, Y(7) => mux_out_12_7_port, 
                           Y(6) => mux_out_12_6_port, Y(5) => mux_out_12_5_port
                           , Y(4) => mux_out_12_4_port, Y(3) => 
                           mux_out_12_3_port, Y(2) => mux_out_12_2_port, Y(1) 
                           => mux_out_12_1_port, Y(0) => mux_out_12_0_port);
   mux_i_13 : MUX51_GENERIC_N64_3 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n576, B(62) => n576, B(61) 
                           => n576, B(60) => n576, B(59) => n576, B(58) => n575
                           , B(57) => n575, B(56) => n501, B(55) => n491, B(54)
                           => n481, B(53) => n471, B(52) => n461, B(51) => n451
                           , B(50) => n441, B(49) => n431, B(48) => n421, B(47)
                           => n411, B(46) => n401, B(45) => n391, B(44) => n381
                           , B(43) => n371, B(42) => n361, B(41) => n351, B(40)
                           => n341, B(39) => n331, B(38) => n321, B(37) => n311
                           , B(36) => n301, B(35) => n291, B(34) => n281, B(33)
                           => n271, B(32) => n261, B(31) => n251, B(30) => n241
                           , B(29) => n231, B(28) => n221, B(27) => n211, B(26)
                           => n201, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic0_port, C(63) => n650, C(62) => n650, C(61) 
                           => n650, C(60) => n650, C(59) => n650, C(58) => n651
                           , C(57) => n651, C(56) => n505, C(55) => n495, C(54)
                           => n485, C(53) => n475, C(52) => n465, C(51) => n455
                           , C(50) => n445, C(49) => n435, C(48) => n425, C(47)
                           => n415, C(46) => n405, C(45) => n395, C(44) => n385
                           , C(43) => n375, C(42) => n365, C(41) => n355, C(40)
                           => n345, C(39) => n335, C(38) => n325, C(37) => n315
                           , C(36) => n305, C(35) => n295, C(34) => n285, C(33)
                           => n275, C(32) => n265, C(31) => n255, C(30) => n245
                           , C(29) => n235, C(28) => n225, C(27) => n215, C(26)
                           => n205, C(25) => X_Logic1_port, C(24) => 
                           X_Logic1_port, C(23) => X_Logic1_port, C(22) => 
                           X_Logic1_port, C(21) => X_Logic1_port, C(20) => 
                           X_Logic1_port, C(19) => X_Logic1_port, C(18) => 
                           X_Logic1_port, C(17) => X_Logic1_port, C(16) => 
                           X_Logic1_port, C(15) => X_Logic1_port, C(14) => 
                           X_Logic1_port, C(13) => X_Logic1_port, C(12) => 
                           X_Logic1_port, C(11) => X_Logic1_port, C(10) => 
                           X_Logic1_port, C(9) => X_Logic1_port, C(8) => 
                           X_Logic1_port, C(7) => X_Logic1_port, C(6) => 
                           X_Logic1_port, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n575, D(62) => n575, D(61) 
                           => n575, D(60) => n575, D(59) => n575, D(58) => n574
                           , D(57) => n501, D(56) => n491, D(55) => n481, D(54)
                           => n471, D(53) => n461, D(52) => n451, D(51) => n441
                           , D(50) => n431, D(49) => n421, D(48) => n411, D(47)
                           => n401, D(46) => n391, D(45) => n381, D(44) => n371
                           , D(43) => n361, D(42) => n351, D(41) => n341, D(40)
                           => n331, D(39) => n321, D(38) => n311, D(37) => n301
                           , D(36) => n291, D(35) => n281, D(34) => n271, D(33)
                           => n261, D(32) => n251, D(31) => n241, D(30) => n231
                           , D(29) => n221, D(28) => n211, D(27) => n201, D(26)
                           => X_Logic0_port, D(25) => X_Logic0_port, D(24) => 
                           X_Logic0_port, D(23) => X_Logic0_port, D(22) => 
                           X_Logic0_port, D(21) => X_Logic0_port, D(20) => 
                           X_Logic0_port, D(19) => X_Logic0_port, D(18) => 
                           X_Logic0_port, D(17) => X_Logic0_port, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(63) => n668, E(62) => n668, E(61) 
                           => n668, E(60) => n668, E(59) => n668, E(58) => n668
                           , E(57) => n506, E(56) => n496, E(55) => n486, E(54)
                           => n476, E(53) => n466, E(52) => n456, E(51) => n446
                           , E(50) => n436, E(49) => n426, E(48) => n416, E(47)
                           => n406, E(46) => n396, E(45) => n386, E(44) => n376
                           , E(43) => n366, E(42) => n356, E(41) => n346, E(40)
                           => n336, E(39) => n326, E(38) => n316, E(37) => n306
                           , E(36) => n296, E(35) => n286, E(34) => n276, E(33)
                           => n266, E(32) => n256, E(31) => n246, E(30) => n236
                           , E(29) => n226, E(28) => n216, E(27) => n206, E(26)
                           => X_Logic1_port, E(25) => X_Logic1_port, E(24) => 
                           X_Logic1_port, E(23) => X_Logic1_port, E(22) => 
                           X_Logic1_port, E(21) => X_Logic1_port, E(20) => 
                           X_Logic1_port, E(19) => X_Logic1_port, E(18) => 
                           X_Logic1_port, E(17) => X_Logic1_port, E(16) => 
                           X_Logic1_port, E(15) => X_Logic1_port, E(14) => 
                           X_Logic1_port, E(13) => X_Logic1_port, E(12) => 
                           X_Logic1_port, E(11) => X_Logic1_port, E(10) => 
                           X_Logic1_port, E(9) => X_Logic1_port, E(8) => 
                           X_Logic1_port, E(7) => X_Logic1_port, E(6) => 
                           X_Logic1_port, E(5) => X_Logic1_port, E(4) => 
                           X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_41_port, SEL(1)
                           => encoder_out_40_port, SEL(0) => 
                           encoder_out_39_port, Y(63) => mux_out_13_63_port, 
                           Y(62) => mux_out_13_62_port, Y(61) => 
                           mux_out_13_61_port, Y(60) => mux_out_13_60_port, 
                           Y(59) => mux_out_13_59_port, Y(58) => 
                           mux_out_13_58_port, Y(57) => mux_out_13_57_port, 
                           Y(56) => mux_out_13_56_port, Y(55) => 
                           mux_out_13_55_port, Y(54) => mux_out_13_54_port, 
                           Y(53) => mux_out_13_53_port, Y(52) => 
                           mux_out_13_52_port, Y(51) => mux_out_13_51_port, 
                           Y(50) => mux_out_13_50_port, Y(49) => 
                           mux_out_13_49_port, Y(48) => mux_out_13_48_port, 
                           Y(47) => mux_out_13_47_port, Y(46) => 
                           mux_out_13_46_port, Y(45) => mux_out_13_45_port, 
                           Y(44) => mux_out_13_44_port, Y(43) => 
                           mux_out_13_43_port, Y(42) => mux_out_13_42_port, 
                           Y(41) => mux_out_13_41_port, Y(40) => 
                           mux_out_13_40_port, Y(39) => mux_out_13_39_port, 
                           Y(38) => mux_out_13_38_port, Y(37) => 
                           mux_out_13_37_port, Y(36) => mux_out_13_36_port, 
                           Y(35) => mux_out_13_35_port, Y(34) => 
                           mux_out_13_34_port, Y(33) => mux_out_13_33_port, 
                           Y(32) => mux_out_13_32_port, Y(31) => 
                           mux_out_13_31_port, Y(30) => mux_out_13_30_port, 
                           Y(29) => mux_out_13_29_port, Y(28) => 
                           mux_out_13_28_port, Y(27) => mux_out_13_27_port, 
                           Y(26) => mux_out_13_26_port, Y(25) => 
                           mux_out_13_25_port, Y(24) => mux_out_13_24_port, 
                           Y(23) => mux_out_13_23_port, Y(22) => 
                           mux_out_13_22_port, Y(21) => mux_out_13_21_port, 
                           Y(20) => mux_out_13_20_port, Y(19) => 
                           mux_out_13_19_port, Y(18) => mux_out_13_18_port, 
                           Y(17) => mux_out_13_17_port, Y(16) => 
                           mux_out_13_16_port, Y(15) => mux_out_13_15_port, 
                           Y(14) => mux_out_13_14_port, Y(13) => 
                           mux_out_13_13_port, Y(12) => mux_out_13_12_port, 
                           Y(11) => mux_out_13_11_port, Y(10) => 
                           mux_out_13_10_port, Y(9) => mux_out_13_9_port, Y(8) 
                           => mux_out_13_8_port, Y(7) => mux_out_13_7_port, 
                           Y(6) => mux_out_13_6_port, Y(5) => mux_out_13_5_port
                           , Y(4) => mux_out_13_4_port, Y(3) => 
                           mux_out_13_3_port, Y(2) => mux_out_13_2_port, Y(1) 
                           => mux_out_13_1_port, Y(0) => mux_out_13_0_port);
   mux_i_14 : MUX51_GENERIC_N64_2 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n577, B(62) => n577, B(61) 
                           => n577, B(60) => n577, B(59) => n577, B(58) => n501
                           , B(57) => n491, B(56) => n481, B(55) => n471, B(54)
                           => n461, B(53) => n451, B(52) => n441, B(51) => n431
                           , B(50) => n421, B(49) => n411, B(48) => n401, B(47)
                           => n391, B(46) => n381, B(45) => n371, B(44) => n361
                           , B(43) => n351, B(42) => n341, B(41) => n331, B(40)
                           => n321, B(39) => n311, B(38) => n301, B(37) => n291
                           , B(36) => n281, B(35) => n271, B(34) => n261, B(33)
                           => n251, B(32) => n241, B(31) => n231, B(30) => n221
                           , B(29) => n211, B(28) => n201, B(27) => 
                           X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
                           X_Logic0_port, B(24) => X_Logic0_port, B(23) => 
                           X_Logic0_port, B(22) => X_Logic0_port, B(21) => 
                           X_Logic0_port, B(20) => X_Logic0_port, B(19) => 
                           X_Logic0_port, B(18) => X_Logic0_port, B(17) => 
                           X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
                           X_Logic0_port, B(14) => X_Logic0_port, B(13) => 
                           X_Logic0_port, B(12) => X_Logic0_port, B(11) => 
                           X_Logic0_port, B(10) => X_Logic0_port, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(63) => n651,
                           C(62) => n651, C(61) => n651, C(60) => n651, C(59) 
                           => n651, C(58) => n505, C(57) => n495, C(56) => n485
                           , C(55) => n475, C(54) => n465, C(53) => n455, C(52)
                           => n445, C(51) => n435, C(50) => n425, C(49) => n415
                           , C(48) => n405, C(47) => n395, C(46) => n385, C(45)
                           => n375, C(44) => n365, C(43) => n355, C(42) => n345
                           , C(41) => n335, C(40) => n325, C(39) => n315, C(38)
                           => n305, C(37) => n295, C(36) => n285, C(35) => n275
                           , C(34) => n265, C(33) => n255, C(32) => n245, C(31)
                           => n235, C(30) => n225, C(29) => n215, C(28) => n205
                           , C(27) => X_Logic1_port, C(26) => X_Logic1_port, 
                           C(25) => X_Logic1_port, C(24) => X_Logic1_port, 
                           C(23) => X_Logic1_port, C(22) => X_Logic1_port, 
                           C(21) => X_Logic1_port, C(20) => X_Logic1_port, 
                           C(19) => X_Logic1_port, C(18) => X_Logic1_port, 
                           C(17) => X_Logic1_port, C(16) => X_Logic1_port, 
                           C(15) => X_Logic1_port, C(14) => X_Logic1_port, 
                           C(13) => X_Logic1_port, C(12) => X_Logic1_port, 
                           C(11) => X_Logic1_port, C(10) => X_Logic1_port, C(9)
                           => X_Logic1_port, C(8) => X_Logic1_port, C(7) => 
                           X_Logic1_port, C(6) => X_Logic1_port, C(5) => 
                           X_Logic1_port, C(4) => X_Logic1_port, C(3) => 
                           X_Logic1_port, C(2) => X_Logic1_port, C(1) => 
                           X_Logic1_port, C(0) => X_Logic1_port, D(63) => n577,
                           D(62) => n577, D(61) => n576, D(60) => n576, D(59) 
                           => n501, D(58) => n491, D(57) => n481, D(56) => n471
                           , D(55) => n461, D(54) => n451, D(53) => n441, D(52)
                           => n431, D(51) => n421, D(50) => n411, D(49) => n401
                           , D(48) => n391, D(47) => n381, D(46) => n371, D(45)
                           => n361, D(44) => n351, D(43) => n341, D(42) => n331
                           , D(41) => n321, D(40) => n311, D(39) => n301, D(38)
                           => n291, D(37) => n281, D(36) => n271, D(35) => n261
                           , D(34) => n251, D(33) => n241, D(32) => n231, D(31)
                           => n221, D(30) => n211, D(29) => n201, D(28) => 
                           X_Logic0_port, D(27) => X_Logic0_port, D(26) => 
                           X_Logic0_port, D(25) => X_Logic0_port, D(24) => 
                           X_Logic0_port, D(23) => X_Logic0_port, D(22) => 
                           X_Logic0_port, D(21) => X_Logic0_port, D(20) => 
                           X_Logic0_port, D(19) => X_Logic0_port, D(18) => 
                           X_Logic0_port, D(17) => X_Logic0_port, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(63) => n668, E(62) => n669, E(61) 
                           => n669, E(60) => n669, E(59) => n506, E(58) => n496
                           , E(57) => n486, E(56) => n476, E(55) => n466, E(54)
                           => n456, E(53) => n446, E(52) => n436, E(51) => n426
                           , E(50) => n416, E(49) => n406, E(48) => n396, E(47)
                           => n386, E(46) => n376, E(45) => n366, E(44) => n356
                           , E(43) => n346, E(42) => n336, E(41) => n326, E(40)
                           => n316, E(39) => n306, E(38) => n296, E(37) => n286
                           , E(36) => n276, E(35) => n266, E(34) => n256, E(33)
                           => n246, E(32) => n236, E(31) => n226, E(30) => n216
                           , E(29) => n206, E(28) => X_Logic1_port, E(27) => 
                           X_Logic1_port, E(26) => X_Logic1_port, E(25) => 
                           X_Logic1_port, E(24) => X_Logic1_port, E(23) => 
                           X_Logic1_port, E(22) => X_Logic1_port, E(21) => 
                           X_Logic1_port, E(20) => X_Logic1_port, E(19) => 
                           X_Logic1_port, E(18) => X_Logic1_port, E(17) => 
                           X_Logic1_port, E(16) => X_Logic1_port, E(15) => 
                           X_Logic1_port, E(14) => X_Logic1_port, E(13) => 
                           X_Logic1_port, E(12) => X_Logic1_port, E(11) => 
                           X_Logic1_port, E(10) => X_Logic1_port, E(9) => 
                           X_Logic1_port, E(8) => X_Logic1_port, E(7) => 
                           X_Logic1_port, E(6) => X_Logic1_port, E(5) => 
                           X_Logic1_port, E(4) => X_Logic1_port, E(3) => 
                           X_Logic1_port, E(2) => X_Logic1_port, E(1) => 
                           X_Logic1_port, E(0) => X_Logic1_port, SEL(2) => 
                           encoder_out_44_port, SEL(1) => encoder_out_43_port, 
                           SEL(0) => encoder_out_42_port, Y(63) => 
                           mux_out_14_63_port, Y(62) => mux_out_14_62_port, 
                           Y(61) => mux_out_14_61_port, Y(60) => 
                           mux_out_14_60_port, Y(59) => mux_out_14_59_port, 
                           Y(58) => mux_out_14_58_port, Y(57) => 
                           mux_out_14_57_port, Y(56) => mux_out_14_56_port, 
                           Y(55) => mux_out_14_55_port, Y(54) => 
                           mux_out_14_54_port, Y(53) => mux_out_14_53_port, 
                           Y(52) => mux_out_14_52_port, Y(51) => 
                           mux_out_14_51_port, Y(50) => mux_out_14_50_port, 
                           Y(49) => mux_out_14_49_port, Y(48) => 
                           mux_out_14_48_port, Y(47) => mux_out_14_47_port, 
                           Y(46) => mux_out_14_46_port, Y(45) => 
                           mux_out_14_45_port, Y(44) => mux_out_14_44_port, 
                           Y(43) => mux_out_14_43_port, Y(42) => 
                           mux_out_14_42_port, Y(41) => mux_out_14_41_port, 
                           Y(40) => mux_out_14_40_port, Y(39) => 
                           mux_out_14_39_port, Y(38) => mux_out_14_38_port, 
                           Y(37) => mux_out_14_37_port, Y(36) => 
                           mux_out_14_36_port, Y(35) => mux_out_14_35_port, 
                           Y(34) => mux_out_14_34_port, Y(33) => 
                           mux_out_14_33_port, Y(32) => mux_out_14_32_port, 
                           Y(31) => mux_out_14_31_port, Y(30) => 
                           mux_out_14_30_port, Y(29) => mux_out_14_29_port, 
                           Y(28) => mux_out_14_28_port, Y(27) => 
                           mux_out_14_27_port, Y(26) => mux_out_14_26_port, 
                           Y(25) => mux_out_14_25_port, Y(24) => 
                           mux_out_14_24_port, Y(23) => mux_out_14_23_port, 
                           Y(22) => mux_out_14_22_port, Y(21) => 
                           mux_out_14_21_port, Y(20) => mux_out_14_20_port, 
                           Y(19) => mux_out_14_19_port, Y(18) => 
                           mux_out_14_18_port, Y(17) => mux_out_14_17_port, 
                           Y(16) => mux_out_14_16_port, Y(15) => 
                           mux_out_14_15_port, Y(14) => mux_out_14_14_port, 
                           Y(13) => mux_out_14_13_port, Y(12) => 
                           mux_out_14_12_port, Y(11) => mux_out_14_11_port, 
                           Y(10) => mux_out_14_10_port, Y(9) => 
                           mux_out_14_9_port, Y(8) => mux_out_14_8_port, Y(7) 
                           => mux_out_14_7_port, Y(6) => mux_out_14_6_port, 
                           Y(5) => mux_out_14_5_port, Y(4) => mux_out_14_4_port
                           , Y(3) => mux_out_14_3_port, Y(2) => 
                           mux_out_14_2_port, Y(1) => mux_out_14_1_port, Y(0) 
                           => mux_out_14_0_port);
   mux_i_15 : MUX51_GENERIC_N64_1 port map( A(63) => X_Logic0_port, A(62) => 
                           X_Logic0_port, A(61) => X_Logic0_port, A(60) => 
                           X_Logic0_port, A(59) => X_Logic0_port, A(58) => 
                           X_Logic0_port, A(57) => X_Logic0_port, A(56) => 
                           X_Logic0_port, A(55) => X_Logic0_port, A(54) => 
                           X_Logic0_port, A(53) => X_Logic0_port, A(52) => 
                           X_Logic0_port, A(51) => X_Logic0_port, A(50) => 
                           X_Logic0_port, A(49) => X_Logic0_port, A(48) => 
                           X_Logic0_port, A(47) => X_Logic0_port, A(46) => 
                           X_Logic0_port, A(45) => X_Logic0_port, A(44) => 
                           X_Logic0_port, A(43) => X_Logic0_port, A(42) => 
                           X_Logic0_port, A(41) => X_Logic0_port, A(40) => 
                           X_Logic0_port, A(39) => X_Logic0_port, A(38) => 
                           X_Logic0_port, A(37) => X_Logic0_port, A(36) => 
                           X_Logic0_port, A(35) => X_Logic0_port, A(34) => 
                           X_Logic0_port, A(33) => X_Logic0_port, A(32) => 
                           X_Logic0_port, A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(63) => n578, B(62) => n578, B(61) 
                           => n578, B(60) => n502, B(59) => n492, B(58) => n482
                           , B(57) => n472, B(56) => n462, B(55) => n452, B(54)
                           => n442, B(53) => n432, B(52) => n422, B(51) => n412
                           , B(50) => n402, B(49) => n392, B(48) => n382, B(47)
                           => n372, B(46) => n362, B(45) => n352, B(44) => n342
                           , B(43) => n332, B(42) => n322, B(41) => n312, B(40)
                           => n302, B(39) => n292, B(38) => n282, B(37) => n272
                           , B(36) => n262, B(35) => n252, B(34) => n242, B(33)
                           => n232, B(32) => n222, B(31) => n212, B(30) => n202
                           , B(29) => X_Logic0_port, B(28) => X_Logic0_port, 
                           B(27) => X_Logic0_port, B(26) => X_Logic0_port, 
                           B(25) => X_Logic0_port, B(24) => X_Logic0_port, 
                           B(23) => X_Logic0_port, B(22) => X_Logic0_port, 
                           B(21) => X_Logic0_port, B(20) => X_Logic0_port, 
                           B(19) => X_Logic0_port, B(18) => X_Logic0_port, 
                           B(17) => X_Logic0_port, B(16) => X_Logic0_port, 
                           B(15) => X_Logic0_port, B(14) => X_Logic0_port, 
                           B(13) => X_Logic0_port, B(12) => X_Logic0_port, 
                           B(11) => X_Logic0_port, B(10) => X_Logic0_port, B(9)
                           => X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic0_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, C(63) => n651,
                           C(62) => n651, C(61) => n636, C(60) => n505, C(59) 
                           => n495, C(58) => n485, C(57) => n475, C(56) => n465
                           , C(55) => n455, C(54) => n445, C(53) => n435, C(52)
                           => n425, C(51) => n415, C(50) => n405, C(49) => n395
                           , C(48) => n385, C(47) => n375, C(46) => n365, C(45)
                           => n355, C(44) => n345, C(43) => n335, C(42) => n325
                           , C(41) => n315, C(40) => n305, C(39) => n295, C(38)
                           => n285, C(37) => n275, C(36) => n265, C(35) => n255
                           , C(34) => n245, C(33) => n235, C(32) => n225, C(31)
                           => n215, C(30) => n205, C(29) => X_Logic1_port, 
                           C(28) => X_Logic1_port, C(27) => X_Logic1_port, 
                           C(26) => X_Logic1_port, C(25) => X_Logic1_port, 
                           C(24) => X_Logic1_port, C(23) => X_Logic1_port, 
                           C(22) => X_Logic1_port, C(21) => X_Logic1_port, 
                           C(20) => X_Logic1_port, C(19) => X_Logic1_port, 
                           C(18) => X_Logic1_port, C(17) => X_Logic1_port, 
                           C(16) => X_Logic1_port, C(15) => X_Logic1_port, 
                           C(14) => X_Logic1_port, C(13) => X_Logic1_port, 
                           C(12) => X_Logic1_port, C(11) => X_Logic1_port, 
                           C(10) => X_Logic1_port, C(9) => X_Logic1_port, C(8) 
                           => X_Logic1_port, C(7) => X_Logic1_port, C(6) => 
                           X_Logic1_port, C(5) => X_Logic1_port, C(4) => 
                           X_Logic1_port, C(3) => X_Logic1_port, C(2) => 
                           X_Logic1_port, C(1) => X_Logic1_port, C(0) => 
                           X_Logic1_port, D(63) => n578, D(62) => n578, D(61) 
                           => n502, D(60) => n492, D(59) => n482, D(58) => n472
                           , D(57) => n462, D(56) => n452, D(55) => n442, D(54)
                           => n432, D(53) => n422, D(52) => n412, D(51) => n402
                           , D(50) => n392, D(49) => n382, D(48) => n372, D(47)
                           => n362, D(46) => n352, D(45) => n342, D(44) => n332
                           , D(43) => n322, D(42) => n312, D(41) => n302, D(40)
                           => n292, D(39) => n282, D(38) => n272, D(37) => n262
                           , D(36) => n252, D(35) => n242, D(34) => n232, D(33)
                           => n222, D(32) => n212, D(31) => n202, D(30) => 
                           X_Logic0_port, D(29) => X_Logic0_port, D(28) => 
                           X_Logic0_port, D(27) => X_Logic0_port, D(26) => 
                           X_Logic0_port, D(25) => X_Logic0_port, D(24) => 
                           X_Logic0_port, D(23) => X_Logic0_port, D(22) => 
                           X_Logic0_port, D(21) => X_Logic0_port, D(20) => 
                           X_Logic0_port, D(19) => X_Logic0_port, D(18) => 
                           X_Logic0_port, D(17) => X_Logic0_port, D(16) => 
                           X_Logic0_port, D(15) => X_Logic0_port, D(14) => 
                           X_Logic0_port, D(13) => X_Logic0_port, D(12) => 
                           X_Logic0_port, D(11) => X_Logic0_port, D(10) => 
                           X_Logic0_port, D(9) => X_Logic0_port, D(8) => 
                           X_Logic0_port, D(7) => X_Logic0_port, D(6) => 
                           X_Logic0_port, D(5) => X_Logic0_port, D(4) => 
                           X_Logic0_port, D(3) => X_Logic0_port, D(2) => 
                           X_Logic0_port, D(1) => X_Logic0_port, D(0) => 
                           X_Logic0_port, E(63) => n669, E(62) => n669, E(61) 
                           => n506, E(60) => n496, E(59) => n486, E(58) => n476
                           , E(57) => n466, E(56) => n456, E(55) => n446, E(54)
                           => n436, E(53) => n426, E(52) => n416, E(51) => n406
                           , E(50) => n396, E(49) => n386, E(48) => n376, E(47)
                           => n366, E(46) => n356, E(45) => n346, E(44) => n336
                           , E(43) => n326, E(42) => n316, E(41) => n306, E(40)
                           => n296, E(39) => n286, E(38) => n276, E(37) => n266
                           , E(36) => n256, E(35) => n246, E(34) => n236, E(33)
                           => n226, E(32) => n216, E(31) => n206, E(30) => 
                           X_Logic1_port, E(29) => X_Logic1_port, E(28) => 
                           X_Logic1_port, E(27) => X_Logic1_port, E(26) => 
                           X_Logic1_port, E(25) => X_Logic1_port, E(24) => 
                           X_Logic1_port, E(23) => X_Logic1_port, E(22) => 
                           X_Logic1_port, E(21) => X_Logic1_port, E(20) => 
                           X_Logic1_port, E(19) => X_Logic1_port, E(18) => 
                           X_Logic1_port, E(17) => X_Logic1_port, E(16) => 
                           X_Logic1_port, E(15) => X_Logic1_port, E(14) => 
                           X_Logic1_port, E(13) => X_Logic1_port, E(12) => 
                           X_Logic1_port, E(11) => X_Logic1_port, E(10) => 
                           X_Logic1_port, E(9) => X_Logic1_port, E(8) => 
                           X_Logic1_port, E(7) => X_Logic1_port, E(6) => 
                           X_Logic1_port, E(5) => X_Logic1_port, E(4) => 
                           X_Logic1_port, E(3) => X_Logic1_port, E(2) => 
                           X_Logic1_port, E(1) => X_Logic1_port, E(0) => 
                           X_Logic1_port, SEL(2) => encoder_out_47_port, SEL(1)
                           => encoder_out_46_port, SEL(0) => 
                           encoder_out_45_port, Y(63) => mux_out_15_63_port, 
                           Y(62) => mux_out_15_62_port, Y(61) => 
                           mux_out_15_61_port, Y(60) => mux_out_15_60_port, 
                           Y(59) => mux_out_15_59_port, Y(58) => 
                           mux_out_15_58_port, Y(57) => mux_out_15_57_port, 
                           Y(56) => mux_out_15_56_port, Y(55) => 
                           mux_out_15_55_port, Y(54) => mux_out_15_54_port, 
                           Y(53) => mux_out_15_53_port, Y(52) => 
                           mux_out_15_52_port, Y(51) => mux_out_15_51_port, 
                           Y(50) => mux_out_15_50_port, Y(49) => 
                           mux_out_15_49_port, Y(48) => mux_out_15_48_port, 
                           Y(47) => mux_out_15_47_port, Y(46) => 
                           mux_out_15_46_port, Y(45) => mux_out_15_45_port, 
                           Y(44) => mux_out_15_44_port, Y(43) => 
                           mux_out_15_43_port, Y(42) => mux_out_15_42_port, 
                           Y(41) => mux_out_15_41_port, Y(40) => 
                           mux_out_15_40_port, Y(39) => mux_out_15_39_port, 
                           Y(38) => mux_out_15_38_port, Y(37) => 
                           mux_out_15_37_port, Y(36) => mux_out_15_36_port, 
                           Y(35) => mux_out_15_35_port, Y(34) => 
                           mux_out_15_34_port, Y(33) => mux_out_15_33_port, 
                           Y(32) => mux_out_15_32_port, Y(31) => 
                           mux_out_15_31_port, Y(30) => mux_out_15_30_port, 
                           Y(29) => mux_out_15_29_port, Y(28) => 
                           mux_out_15_28_port, Y(27) => mux_out_15_27_port, 
                           Y(26) => mux_out_15_26_port, Y(25) => 
                           mux_out_15_25_port, Y(24) => mux_out_15_24_port, 
                           Y(23) => mux_out_15_23_port, Y(22) => 
                           mux_out_15_22_port, Y(21) => mux_out_15_21_port, 
                           Y(20) => mux_out_15_20_port, Y(19) => 
                           mux_out_15_19_port, Y(18) => mux_out_15_18_port, 
                           Y(17) => mux_out_15_17_port, Y(16) => 
                           mux_out_15_16_port, Y(15) => mux_out_15_15_port, 
                           Y(14) => mux_out_15_14_port, Y(13) => 
                           mux_out_15_13_port, Y(12) => mux_out_15_12_port, 
                           Y(11) => mux_out_15_11_port, Y(10) => 
                           mux_out_15_10_port, Y(9) => mux_out_15_9_port, Y(8) 
                           => mux_out_15_8_port, Y(7) => mux_out_15_7_port, 
                           Y(6) => mux_out_15_6_port, Y(5) => mux_out_15_5_port
                           , Y(4) => mux_out_15_4_port, Y(3) => 
                           mux_out_15_3_port, Y(2) => mux_out_15_2_port, Y(1) 
                           => mux_out_15_1_port, Y(0) => mux_out_15_0_port);
   add_i_0 : RCA_generic_N64_0 port map( A(63) => mux_out_1_63_port, A(62) => 
                           mux_out_1_62_port, A(61) => mux_out_1_61_port, A(60)
                           => mux_out_1_60_port, A(59) => mux_out_1_59_port, 
                           A(58) => mux_out_1_58_port, A(57) => 
                           mux_out_1_57_port, A(56) => mux_out_1_56_port, A(55)
                           => mux_out_1_55_port, A(54) => mux_out_1_54_port, 
                           A(53) => mux_out_1_53_port, A(52) => 
                           mux_out_1_52_port, A(51) => mux_out_1_51_port, A(50)
                           => mux_out_1_50_port, A(49) => mux_out_1_49_port, 
                           A(48) => mux_out_1_48_port, A(47) => 
                           mux_out_1_47_port, A(46) => mux_out_1_46_port, A(45)
                           => mux_out_1_45_port, A(44) => mux_out_1_44_port, 
                           A(43) => mux_out_1_43_port, A(42) => 
                           mux_out_1_42_port, A(41) => mux_out_1_41_port, A(40)
                           => mux_out_1_40_port, A(39) => mux_out_1_39_port, 
                           A(38) => mux_out_1_38_port, A(37) => 
                           mux_out_1_37_port, A(36) => mux_out_1_36_port, A(35)
                           => mux_out_1_35_port, A(34) => mux_out_1_34_port, 
                           A(33) => mux_out_1_33_port, A(32) => 
                           mux_out_1_32_port, A(31) => mux_out_1_31_port, A(30)
                           => mux_out_1_30_port, A(29) => mux_out_1_29_port, 
                           A(28) => mux_out_1_28_port, A(27) => 
                           mux_out_1_27_port, A(26) => mux_out_1_26_port, A(25)
                           => mux_out_1_25_port, A(24) => mux_out_1_24_port, 
                           A(23) => mux_out_1_23_port, A(22) => 
                           mux_out_1_22_port, A(21) => mux_out_1_21_port, A(20)
                           => mux_out_1_20_port, A(19) => mux_out_1_19_port, 
                           A(18) => mux_out_1_18_port, A(17) => 
                           mux_out_1_17_port, A(16) => mux_out_1_16_port, A(15)
                           => mux_out_1_15_port, A(14) => mux_out_1_14_port, 
                           A(13) => mux_out_1_13_port, A(12) => 
                           mux_out_1_12_port, A(11) => mux_out_1_11_port, A(10)
                           => mux_out_1_10_port, A(9) => mux_out_1_9_port, A(8)
                           => mux_out_1_8_port, A(7) => mux_out_1_7_port, A(6) 
                           => mux_out_1_6_port, A(5) => mux_out_1_5_port, A(4) 
                           => mux_out_1_4_port, A(3) => mux_out_1_3_port, A(2) 
                           => mux_out_1_2_port, A(1) => mux_out_1_1_port, A(0) 
                           => mux_out_1_0_port, B(63) => add_in_0_63_port, 
                           B(62) => add_in_0_62_port, B(61) => add_in_0_61_port
                           , B(60) => add_in_0_60_port, B(59) => 
                           add_in_0_59_port, B(58) => add_in_0_58_port, B(57) 
                           => add_in_0_57_port, B(56) => add_in_0_56_port, 
                           B(55) => add_in_0_55_port, B(54) => add_in_0_54_port
                           , B(53) => add_in_0_53_port, B(52) => 
                           add_in_0_52_port, B(51) => add_in_0_51_port, B(50) 
                           => add_in_0_50_port, B(49) => add_in_0_49_port, 
                           B(48) => add_in_0_48_port, B(47) => add_in_0_47_port
                           , B(46) => add_in_0_46_port, B(45) => 
                           add_in_0_45_port, B(44) => add_in_0_44_port, B(43) 
                           => add_in_0_43_port, B(42) => add_in_0_42_port, 
                           B(41) => add_in_0_41_port, B(40) => add_in_0_40_port
                           , B(39) => add_in_0_39_port, B(38) => 
                           add_in_0_38_port, B(37) => add_in_0_37_port, B(36) 
                           => add_in_0_36_port, B(35) => add_in_0_35_port, 
                           B(34) => add_in_0_34_port, B(33) => add_in_0_33_port
                           , B(32) => add_in_0_32_port, B(31) => 
                           add_in_0_31_port, B(30) => add_in_0_30_port, B(29) 
                           => add_in_0_29_port, B(28) => add_in_0_28_port, 
                           B(27) => add_in_0_27_port, B(26) => add_in_0_26_port
                           , B(25) => add_in_0_25_port, B(24) => 
                           add_in_0_24_port, B(23) => add_in_0_23_port, B(22) 
                           => add_in_0_22_port, B(21) => add_in_0_21_port, 
                           B(20) => add_in_0_20_port, B(19) => add_in_0_19_port
                           , B(18) => add_in_0_18_port, B(17) => 
                           add_in_0_17_port, B(16) => add_in_0_16_port, B(15) 
                           => add_in_0_15_port, B(14) => add_in_0_14_port, 
                           B(13) => add_in_0_13_port, B(12) => add_in_0_12_port
                           , B(11) => add_in_0_11_port, B(10) => 
                           add_in_0_10_port, B(9) => add_in_0_9_port, B(8) => 
                           add_in_0_8_port, B(7) => add_in_0_7_port, B(6) => 
                           add_in_0_6_port, B(5) => add_in_0_5_port, B(4) => 
                           add_in_0_4_port, B(3) => add_in_0_3_port, B(2) => 
                           add_in_0_2_port, B(1) => add_in_0_1_port, B(0) => 
                           add_in_0_0_port, Ci => B(1), S(63) => 
                           add_in_1_63_port, S(62) => add_in_1_62_port, S(61) 
                           => add_in_1_61_port, S(60) => add_in_1_60_port, 
                           S(59) => add_in_1_59_port, S(58) => add_in_1_58_port
                           , S(57) => add_in_1_57_port, S(56) => 
                           add_in_1_56_port, S(55) => add_in_1_55_port, S(54) 
                           => add_in_1_54_port, S(53) => add_in_1_53_port, 
                           S(52) => add_in_1_52_port, S(51) => add_in_1_51_port
                           , S(50) => add_in_1_50_port, S(49) => 
                           add_in_1_49_port, S(48) => add_in_1_48_port, S(47) 
                           => add_in_1_47_port, S(46) => add_in_1_46_port, 
                           S(45) => add_in_1_45_port, S(44) => add_in_1_44_port
                           , S(43) => add_in_1_43_port, S(42) => 
                           add_in_1_42_port, S(41) => add_in_1_41_port, S(40) 
                           => add_in_1_40_port, S(39) => add_in_1_39_port, 
                           S(38) => add_in_1_38_port, S(37) => add_in_1_37_port
                           , S(36) => add_in_1_36_port, S(35) => 
                           add_in_1_35_port, S(34) => add_in_1_34_port, S(33) 
                           => add_in_1_33_port, S(32) => add_in_1_32_port, 
                           S(31) => add_in_1_31_port, S(30) => add_in_1_30_port
                           , S(29) => add_in_1_29_port, S(28) => 
                           add_in_1_28_port, S(27) => add_in_1_27_port, S(26) 
                           => add_in_1_26_port, S(25) => add_in_1_25_port, 
                           S(24) => add_in_1_24_port, S(23) => add_in_1_23_port
                           , S(22) => add_in_1_22_port, S(21) => 
                           add_in_1_21_port, S(20) => add_in_1_20_port, S(19) 
                           => add_in_1_19_port, S(18) => add_in_1_18_port, 
                           S(17) => add_in_1_17_port, S(16) => add_in_1_16_port
                           , S(15) => add_in_1_15_port, S(14) => 
                           add_in_1_14_port, S(13) => add_in_1_13_port, S(12) 
                           => add_in_1_12_port, S(11) => add_in_1_11_port, 
                           S(10) => add_in_1_10_port, S(9) => add_in_1_9_port, 
                           S(8) => add_in_1_8_port, S(7) => add_in_1_7_port, 
                           S(6) => add_in_1_6_port, S(5) => add_in_1_5_port, 
                           S(4) => add_in_1_4_port, S(3) => add_in_1_3_port, 
                           S(2) => add_in_1_2_port, S(1) => add_in_1_1_port, 
                           S(0) => add_in_1_0_port, Co => net21320);
   add_i_1 : RCA_generic_N64_14 port map( A(63) => mux_out_2_63_port, A(62) => 
                           mux_out_2_62_port, A(61) => mux_out_2_61_port, A(60)
                           => mux_out_2_60_port, A(59) => mux_out_2_59_port, 
                           A(58) => mux_out_2_58_port, A(57) => 
                           mux_out_2_57_port, A(56) => mux_out_2_56_port, A(55)
                           => mux_out_2_55_port, A(54) => mux_out_2_54_port, 
                           A(53) => mux_out_2_53_port, A(52) => 
                           mux_out_2_52_port, A(51) => mux_out_2_51_port, A(50)
                           => mux_out_2_50_port, A(49) => mux_out_2_49_port, 
                           A(48) => mux_out_2_48_port, A(47) => 
                           mux_out_2_47_port, A(46) => mux_out_2_46_port, A(45)
                           => mux_out_2_45_port, A(44) => mux_out_2_44_port, 
                           A(43) => mux_out_2_43_port, A(42) => 
                           mux_out_2_42_port, A(41) => mux_out_2_41_port, A(40)
                           => mux_out_2_40_port, A(39) => mux_out_2_39_port, 
                           A(38) => mux_out_2_38_port, A(37) => 
                           mux_out_2_37_port, A(36) => mux_out_2_36_port, A(35)
                           => mux_out_2_35_port, A(34) => mux_out_2_34_port, 
                           A(33) => mux_out_2_33_port, A(32) => 
                           mux_out_2_32_port, A(31) => mux_out_2_31_port, A(30)
                           => mux_out_2_30_port, A(29) => mux_out_2_29_port, 
                           A(28) => mux_out_2_28_port, A(27) => 
                           mux_out_2_27_port, A(26) => mux_out_2_26_port, A(25)
                           => mux_out_2_25_port, A(24) => mux_out_2_24_port, 
                           A(23) => mux_out_2_23_port, A(22) => 
                           mux_out_2_22_port, A(21) => mux_out_2_21_port, A(20)
                           => mux_out_2_20_port, A(19) => mux_out_2_19_port, 
                           A(18) => mux_out_2_18_port, A(17) => 
                           mux_out_2_17_port, A(16) => mux_out_2_16_port, A(15)
                           => mux_out_2_15_port, A(14) => mux_out_2_14_port, 
                           A(13) => mux_out_2_13_port, A(12) => 
                           mux_out_2_12_port, A(11) => mux_out_2_11_port, A(10)
                           => mux_out_2_10_port, A(9) => mux_out_2_9_port, A(8)
                           => mux_out_2_8_port, A(7) => mux_out_2_7_port, A(6) 
                           => mux_out_2_6_port, A(5) => mux_out_2_5_port, A(4) 
                           => mux_out_2_4_port, A(3) => mux_out_2_3_port, A(2) 
                           => mux_out_2_2_port, A(1) => mux_out_2_1_port, A(0) 
                           => mux_out_2_0_port, B(63) => add_in_1_63_port, 
                           B(62) => add_in_1_62_port, B(61) => add_in_1_61_port
                           , B(60) => add_in_1_60_port, B(59) => 
                           add_in_1_59_port, B(58) => add_in_1_58_port, B(57) 
                           => add_in_1_57_port, B(56) => add_in_1_56_port, 
                           B(55) => add_in_1_55_port, B(54) => add_in_1_54_port
                           , B(53) => add_in_1_53_port, B(52) => 
                           add_in_1_52_port, B(51) => add_in_1_51_port, B(50) 
                           => add_in_1_50_port, B(49) => add_in_1_49_port, 
                           B(48) => add_in_1_48_port, B(47) => add_in_1_47_port
                           , B(46) => add_in_1_46_port, B(45) => 
                           add_in_1_45_port, B(44) => add_in_1_44_port, B(43) 
                           => add_in_1_43_port, B(42) => add_in_1_42_port, 
                           B(41) => add_in_1_41_port, B(40) => add_in_1_40_port
                           , B(39) => add_in_1_39_port, B(38) => 
                           add_in_1_38_port, B(37) => add_in_1_37_port, B(36) 
                           => add_in_1_36_port, B(35) => add_in_1_35_port, 
                           B(34) => add_in_1_34_port, B(33) => add_in_1_33_port
                           , B(32) => add_in_1_32_port, B(31) => 
                           add_in_1_31_port, B(30) => add_in_1_30_port, B(29) 
                           => add_in_1_29_port, B(28) => add_in_1_28_port, 
                           B(27) => add_in_1_27_port, B(26) => add_in_1_26_port
                           , B(25) => add_in_1_25_port, B(24) => 
                           add_in_1_24_port, B(23) => add_in_1_23_port, B(22) 
                           => add_in_1_22_port, B(21) => add_in_1_21_port, 
                           B(20) => add_in_1_20_port, B(19) => add_in_1_19_port
                           , B(18) => add_in_1_18_port, B(17) => 
                           add_in_1_17_port, B(16) => add_in_1_16_port, B(15) 
                           => add_in_1_15_port, B(14) => add_in_1_14_port, 
                           B(13) => add_in_1_13_port, B(12) => add_in_1_12_port
                           , B(11) => add_in_1_11_port, B(10) => 
                           add_in_1_10_port, B(9) => add_in_1_9_port, B(8) => 
                           add_in_1_8_port, B(7) => add_in_1_7_port, B(6) => 
                           add_in_1_6_port, B(5) => add_in_1_5_port, B(4) => 
                           add_in_1_4_port, B(3) => add_in_1_3_port, B(2) => 
                           add_in_1_2_port, B(1) => add_in_1_1_port, B(0) => 
                           add_in_1_0_port, Ci => mode_1_port, S(63) => 
                           add_in_2_63_port, S(62) => add_in_2_62_port, S(61) 
                           => add_in_2_61_port, S(60) => add_in_2_60_port, 
                           S(59) => add_in_2_59_port, S(58) => add_in_2_58_port
                           , S(57) => add_in_2_57_port, S(56) => 
                           add_in_2_56_port, S(55) => add_in_2_55_port, S(54) 
                           => add_in_2_54_port, S(53) => add_in_2_53_port, 
                           S(52) => add_in_2_52_port, S(51) => add_in_2_51_port
                           , S(50) => add_in_2_50_port, S(49) => 
                           add_in_2_49_port, S(48) => add_in_2_48_port, S(47) 
                           => add_in_2_47_port, S(46) => add_in_2_46_port, 
                           S(45) => add_in_2_45_port, S(44) => add_in_2_44_port
                           , S(43) => add_in_2_43_port, S(42) => 
                           add_in_2_42_port, S(41) => add_in_2_41_port, S(40) 
                           => add_in_2_40_port, S(39) => add_in_2_39_port, 
                           S(38) => add_in_2_38_port, S(37) => add_in_2_37_port
                           , S(36) => add_in_2_36_port, S(35) => 
                           add_in_2_35_port, S(34) => add_in_2_34_port, S(33) 
                           => add_in_2_33_port, S(32) => add_in_2_32_port, 
                           S(31) => add_in_2_31_port, S(30) => add_in_2_30_port
                           , S(29) => add_in_2_29_port, S(28) => 
                           add_in_2_28_port, S(27) => add_in_2_27_port, S(26) 
                           => add_in_2_26_port, S(25) => add_in_2_25_port, 
                           S(24) => add_in_2_24_port, S(23) => add_in_2_23_port
                           , S(22) => add_in_2_22_port, S(21) => 
                           add_in_2_21_port, S(20) => add_in_2_20_port, S(19) 
                           => add_in_2_19_port, S(18) => add_in_2_18_port, 
                           S(17) => add_in_2_17_port, S(16) => add_in_2_16_port
                           , S(15) => add_in_2_15_port, S(14) => 
                           add_in_2_14_port, S(13) => add_in_2_13_port, S(12) 
                           => add_in_2_12_port, S(11) => add_in_2_11_port, 
                           S(10) => add_in_2_10_port, S(9) => add_in_2_9_port, 
                           S(8) => add_in_2_8_port, S(7) => add_in_2_7_port, 
                           S(6) => add_in_2_6_port, S(5) => add_in_2_5_port, 
                           S(4) => add_in_2_4_port, S(3) => add_in_2_3_port, 
                           S(2) => add_in_2_2_port, S(1) => add_in_2_1_port, 
                           S(0) => add_in_2_0_port, Co => net21319);
   add_i_2 : RCA_generic_N64_13 port map( A(63) => mux_out_3_63_port, A(62) => 
                           mux_out_3_62_port, A(61) => mux_out_3_61_port, A(60)
                           => mux_out_3_60_port, A(59) => mux_out_3_59_port, 
                           A(58) => mux_out_3_58_port, A(57) => 
                           mux_out_3_57_port, A(56) => mux_out_3_56_port, A(55)
                           => mux_out_3_55_port, A(54) => mux_out_3_54_port, 
                           A(53) => mux_out_3_53_port, A(52) => 
                           mux_out_3_52_port, A(51) => mux_out_3_51_port, A(50)
                           => mux_out_3_50_port, A(49) => mux_out_3_49_port, 
                           A(48) => mux_out_3_48_port, A(47) => 
                           mux_out_3_47_port, A(46) => mux_out_3_46_port, A(45)
                           => mux_out_3_45_port, A(44) => mux_out_3_44_port, 
                           A(43) => mux_out_3_43_port, A(42) => 
                           mux_out_3_42_port, A(41) => mux_out_3_41_port, A(40)
                           => mux_out_3_40_port, A(39) => mux_out_3_39_port, 
                           A(38) => mux_out_3_38_port, A(37) => 
                           mux_out_3_37_port, A(36) => mux_out_3_36_port, A(35)
                           => mux_out_3_35_port, A(34) => mux_out_3_34_port, 
                           A(33) => mux_out_3_33_port, A(32) => 
                           mux_out_3_32_port, A(31) => mux_out_3_31_port, A(30)
                           => mux_out_3_30_port, A(29) => mux_out_3_29_port, 
                           A(28) => mux_out_3_28_port, A(27) => 
                           mux_out_3_27_port, A(26) => mux_out_3_26_port, A(25)
                           => mux_out_3_25_port, A(24) => mux_out_3_24_port, 
                           A(23) => mux_out_3_23_port, A(22) => 
                           mux_out_3_22_port, A(21) => mux_out_3_21_port, A(20)
                           => mux_out_3_20_port, A(19) => mux_out_3_19_port, 
                           A(18) => mux_out_3_18_port, A(17) => 
                           mux_out_3_17_port, A(16) => mux_out_3_16_port, A(15)
                           => mux_out_3_15_port, A(14) => mux_out_3_14_port, 
                           A(13) => mux_out_3_13_port, A(12) => 
                           mux_out_3_12_port, A(11) => mux_out_3_11_port, A(10)
                           => mux_out_3_10_port, A(9) => mux_out_3_9_port, A(8)
                           => mux_out_3_8_port, A(7) => mux_out_3_7_port, A(6) 
                           => mux_out_3_6_port, A(5) => mux_out_3_5_port, A(4) 
                           => mux_out_3_4_port, A(3) => mux_out_3_3_port, A(2) 
                           => mux_out_3_2_port, A(1) => mux_out_3_1_port, A(0) 
                           => mux_out_3_0_port, B(63) => add_in_2_63_port, 
                           B(62) => add_in_2_62_port, B(61) => add_in_2_61_port
                           , B(60) => add_in_2_60_port, B(59) => 
                           add_in_2_59_port, B(58) => add_in_2_58_port, B(57) 
                           => add_in_2_57_port, B(56) => add_in_2_56_port, 
                           B(55) => add_in_2_55_port, B(54) => add_in_2_54_port
                           , B(53) => add_in_2_53_port, B(52) => 
                           add_in_2_52_port, B(51) => add_in_2_51_port, B(50) 
                           => add_in_2_50_port, B(49) => add_in_2_49_port, 
                           B(48) => add_in_2_48_port, B(47) => add_in_2_47_port
                           , B(46) => add_in_2_46_port, B(45) => 
                           add_in_2_45_port, B(44) => add_in_2_44_port, B(43) 
                           => add_in_2_43_port, B(42) => add_in_2_42_port, 
                           B(41) => add_in_2_41_port, B(40) => add_in_2_40_port
                           , B(39) => add_in_2_39_port, B(38) => 
                           add_in_2_38_port, B(37) => add_in_2_37_port, B(36) 
                           => add_in_2_36_port, B(35) => add_in_2_35_port, 
                           B(34) => add_in_2_34_port, B(33) => add_in_2_33_port
                           , B(32) => add_in_2_32_port, B(31) => 
                           add_in_2_31_port, B(30) => add_in_2_30_port, B(29) 
                           => add_in_2_29_port, B(28) => add_in_2_28_port, 
                           B(27) => add_in_2_27_port, B(26) => add_in_2_26_port
                           , B(25) => add_in_2_25_port, B(24) => 
                           add_in_2_24_port, B(23) => add_in_2_23_port, B(22) 
                           => add_in_2_22_port, B(21) => add_in_2_21_port, 
                           B(20) => add_in_2_20_port, B(19) => add_in_2_19_port
                           , B(18) => add_in_2_18_port, B(17) => 
                           add_in_2_17_port, B(16) => add_in_2_16_port, B(15) 
                           => add_in_2_15_port, B(14) => add_in_2_14_port, 
                           B(13) => add_in_2_13_port, B(12) => add_in_2_12_port
                           , B(11) => add_in_2_11_port, B(10) => 
                           add_in_2_10_port, B(9) => add_in_2_9_port, B(8) => 
                           add_in_2_8_port, B(7) => add_in_2_7_port, B(6) => 
                           add_in_2_6_port, B(5) => add_in_2_5_port, B(4) => 
                           add_in_2_4_port, B(3) => add_in_2_3_port, B(2) => 
                           add_in_2_2_port, B(1) => add_in_2_1_port, B(0) => 
                           add_in_2_0_port, Ci => mode_2_port, S(63) => 
                           add_in_3_63_port, S(62) => add_in_3_62_port, S(61) 
                           => add_in_3_61_port, S(60) => add_in_3_60_port, 
                           S(59) => add_in_3_59_port, S(58) => add_in_3_58_port
                           , S(57) => add_in_3_57_port, S(56) => 
                           add_in_3_56_port, S(55) => add_in_3_55_port, S(54) 
                           => add_in_3_54_port, S(53) => add_in_3_53_port, 
                           S(52) => add_in_3_52_port, S(51) => add_in_3_51_port
                           , S(50) => add_in_3_50_port, S(49) => 
                           add_in_3_49_port, S(48) => add_in_3_48_port, S(47) 
                           => add_in_3_47_port, S(46) => add_in_3_46_port, 
                           S(45) => add_in_3_45_port, S(44) => add_in_3_44_port
                           , S(43) => add_in_3_43_port, S(42) => 
                           add_in_3_42_port, S(41) => add_in_3_41_port, S(40) 
                           => add_in_3_40_port, S(39) => add_in_3_39_port, 
                           S(38) => add_in_3_38_port, S(37) => add_in_3_37_port
                           , S(36) => add_in_3_36_port, S(35) => 
                           add_in_3_35_port, S(34) => add_in_3_34_port, S(33) 
                           => add_in_3_33_port, S(32) => add_in_3_32_port, 
                           S(31) => add_in_3_31_port, S(30) => add_in_3_30_port
                           , S(29) => add_in_3_29_port, S(28) => 
                           add_in_3_28_port, S(27) => add_in_3_27_port, S(26) 
                           => add_in_3_26_port, S(25) => add_in_3_25_port, 
                           S(24) => add_in_3_24_port, S(23) => add_in_3_23_port
                           , S(22) => add_in_3_22_port, S(21) => 
                           add_in_3_21_port, S(20) => add_in_3_20_port, S(19) 
                           => add_in_3_19_port, S(18) => add_in_3_18_port, 
                           S(17) => add_in_3_17_port, S(16) => add_in_3_16_port
                           , S(15) => add_in_3_15_port, S(14) => 
                           add_in_3_14_port, S(13) => add_in_3_13_port, S(12) 
                           => add_in_3_12_port, S(11) => add_in_3_11_port, 
                           S(10) => add_in_3_10_port, S(9) => add_in_3_9_port, 
                           S(8) => add_in_3_8_port, S(7) => add_in_3_7_port, 
                           S(6) => add_in_3_6_port, S(5) => add_in_3_5_port, 
                           S(4) => add_in_3_4_port, S(3) => add_in_3_3_port, 
                           S(2) => add_in_3_2_port, S(1) => add_in_3_1_port, 
                           S(0) => add_in_3_0_port, Co => net21318);
   add_i_3 : RCA_generic_N64_12 port map( A(63) => mux_out_4_63_port, A(62) => 
                           mux_out_4_62_port, A(61) => mux_out_4_61_port, A(60)
                           => mux_out_4_60_port, A(59) => mux_out_4_59_port, 
                           A(58) => mux_out_4_58_port, A(57) => 
                           mux_out_4_57_port, A(56) => mux_out_4_56_port, A(55)
                           => mux_out_4_55_port, A(54) => mux_out_4_54_port, 
                           A(53) => mux_out_4_53_port, A(52) => 
                           mux_out_4_52_port, A(51) => mux_out_4_51_port, A(50)
                           => mux_out_4_50_port, A(49) => mux_out_4_49_port, 
                           A(48) => mux_out_4_48_port, A(47) => 
                           mux_out_4_47_port, A(46) => mux_out_4_46_port, A(45)
                           => mux_out_4_45_port, A(44) => mux_out_4_44_port, 
                           A(43) => mux_out_4_43_port, A(42) => 
                           mux_out_4_42_port, A(41) => mux_out_4_41_port, A(40)
                           => mux_out_4_40_port, A(39) => mux_out_4_39_port, 
                           A(38) => mux_out_4_38_port, A(37) => 
                           mux_out_4_37_port, A(36) => mux_out_4_36_port, A(35)
                           => mux_out_4_35_port, A(34) => mux_out_4_34_port, 
                           A(33) => mux_out_4_33_port, A(32) => 
                           mux_out_4_32_port, A(31) => mux_out_4_31_port, A(30)
                           => mux_out_4_30_port, A(29) => mux_out_4_29_port, 
                           A(28) => mux_out_4_28_port, A(27) => 
                           mux_out_4_27_port, A(26) => mux_out_4_26_port, A(25)
                           => mux_out_4_25_port, A(24) => mux_out_4_24_port, 
                           A(23) => mux_out_4_23_port, A(22) => 
                           mux_out_4_22_port, A(21) => mux_out_4_21_port, A(20)
                           => mux_out_4_20_port, A(19) => mux_out_4_19_port, 
                           A(18) => mux_out_4_18_port, A(17) => 
                           mux_out_4_17_port, A(16) => mux_out_4_16_port, A(15)
                           => mux_out_4_15_port, A(14) => mux_out_4_14_port, 
                           A(13) => mux_out_4_13_port, A(12) => 
                           mux_out_4_12_port, A(11) => mux_out_4_11_port, A(10)
                           => mux_out_4_10_port, A(9) => mux_out_4_9_port, A(8)
                           => mux_out_4_8_port, A(7) => mux_out_4_7_port, A(6) 
                           => mux_out_4_6_port, A(5) => mux_out_4_5_port, A(4) 
                           => mux_out_4_4_port, A(3) => mux_out_4_3_port, A(2) 
                           => mux_out_4_2_port, A(1) => mux_out_4_1_port, A(0) 
                           => mux_out_4_0_port, B(63) => add_in_3_63_port, 
                           B(62) => add_in_3_62_port, B(61) => add_in_3_61_port
                           , B(60) => add_in_3_60_port, B(59) => 
                           add_in_3_59_port, B(58) => add_in_3_58_port, B(57) 
                           => add_in_3_57_port, B(56) => add_in_3_56_port, 
                           B(55) => add_in_3_55_port, B(54) => add_in_3_54_port
                           , B(53) => add_in_3_53_port, B(52) => 
                           add_in_3_52_port, B(51) => add_in_3_51_port, B(50) 
                           => add_in_3_50_port, B(49) => add_in_3_49_port, 
                           B(48) => add_in_3_48_port, B(47) => add_in_3_47_port
                           , B(46) => add_in_3_46_port, B(45) => 
                           add_in_3_45_port, B(44) => add_in_3_44_port, B(43) 
                           => add_in_3_43_port, B(42) => add_in_3_42_port, 
                           B(41) => add_in_3_41_port, B(40) => add_in_3_40_port
                           , B(39) => add_in_3_39_port, B(38) => 
                           add_in_3_38_port, B(37) => add_in_3_37_port, B(36) 
                           => add_in_3_36_port, B(35) => add_in_3_35_port, 
                           B(34) => add_in_3_34_port, B(33) => add_in_3_33_port
                           , B(32) => add_in_3_32_port, B(31) => 
                           add_in_3_31_port, B(30) => add_in_3_30_port, B(29) 
                           => add_in_3_29_port, B(28) => add_in_3_28_port, 
                           B(27) => add_in_3_27_port, B(26) => add_in_3_26_port
                           , B(25) => add_in_3_25_port, B(24) => 
                           add_in_3_24_port, B(23) => add_in_3_23_port, B(22) 
                           => add_in_3_22_port, B(21) => add_in_3_21_port, 
                           B(20) => add_in_3_20_port, B(19) => add_in_3_19_port
                           , B(18) => add_in_3_18_port, B(17) => 
                           add_in_3_17_port, B(16) => add_in_3_16_port, B(15) 
                           => add_in_3_15_port, B(14) => add_in_3_14_port, 
                           B(13) => add_in_3_13_port, B(12) => add_in_3_12_port
                           , B(11) => add_in_3_11_port, B(10) => 
                           add_in_3_10_port, B(9) => add_in_3_9_port, B(8) => 
                           add_in_3_8_port, B(7) => add_in_3_7_port, B(6) => 
                           add_in_3_6_port, B(5) => add_in_3_5_port, B(4) => 
                           add_in_3_4_port, B(3) => add_in_3_3_port, B(2) => 
                           add_in_3_2_port, B(1) => add_in_3_1_port, B(0) => 
                           add_in_3_0_port, Ci => mode_3_port, S(63) => 
                           add_in_4_63_port, S(62) => add_in_4_62_port, S(61) 
                           => add_in_4_61_port, S(60) => add_in_4_60_port, 
                           S(59) => add_in_4_59_port, S(58) => add_in_4_58_port
                           , S(57) => add_in_4_57_port, S(56) => 
                           add_in_4_56_port, S(55) => add_in_4_55_port, S(54) 
                           => add_in_4_54_port, S(53) => add_in_4_53_port, 
                           S(52) => add_in_4_52_port, S(51) => add_in_4_51_port
                           , S(50) => add_in_4_50_port, S(49) => 
                           add_in_4_49_port, S(48) => add_in_4_48_port, S(47) 
                           => add_in_4_47_port, S(46) => add_in_4_46_port, 
                           S(45) => add_in_4_45_port, S(44) => add_in_4_44_port
                           , S(43) => add_in_4_43_port, S(42) => 
                           add_in_4_42_port, S(41) => add_in_4_41_port, S(40) 
                           => add_in_4_40_port, S(39) => add_in_4_39_port, 
                           S(38) => add_in_4_38_port, S(37) => add_in_4_37_port
                           , S(36) => add_in_4_36_port, S(35) => 
                           add_in_4_35_port, S(34) => add_in_4_34_port, S(33) 
                           => add_in_4_33_port, S(32) => add_in_4_32_port, 
                           S(31) => add_in_4_31_port, S(30) => add_in_4_30_port
                           , S(29) => add_in_4_29_port, S(28) => 
                           add_in_4_28_port, S(27) => add_in_4_27_port, S(26) 
                           => add_in_4_26_port, S(25) => add_in_4_25_port, 
                           S(24) => add_in_4_24_port, S(23) => add_in_4_23_port
                           , S(22) => add_in_4_22_port, S(21) => 
                           add_in_4_21_port, S(20) => add_in_4_20_port, S(19) 
                           => add_in_4_19_port, S(18) => add_in_4_18_port, 
                           S(17) => add_in_4_17_port, S(16) => add_in_4_16_port
                           , S(15) => add_in_4_15_port, S(14) => 
                           add_in_4_14_port, S(13) => add_in_4_13_port, S(12) 
                           => add_in_4_12_port, S(11) => add_in_4_11_port, 
                           S(10) => add_in_4_10_port, S(9) => add_in_4_9_port, 
                           S(8) => add_in_4_8_port, S(7) => add_in_4_7_port, 
                           S(6) => add_in_4_6_port, S(5) => add_in_4_5_port, 
                           S(4) => add_in_4_4_port, S(3) => add_in_4_3_port, 
                           S(2) => add_in_4_2_port, S(1) => add_in_4_1_port, 
                           S(0) => add_in_4_0_port, Co => net21317);
   add_i_4 : RCA_generic_N64_11 port map( A(63) => mux_out_5_63_port, A(62) => 
                           mux_out_5_62_port, A(61) => mux_out_5_61_port, A(60)
                           => mux_out_5_60_port, A(59) => mux_out_5_59_port, 
                           A(58) => mux_out_5_58_port, A(57) => 
                           mux_out_5_57_port, A(56) => mux_out_5_56_port, A(55)
                           => mux_out_5_55_port, A(54) => mux_out_5_54_port, 
                           A(53) => mux_out_5_53_port, A(52) => 
                           mux_out_5_52_port, A(51) => mux_out_5_51_port, A(50)
                           => mux_out_5_50_port, A(49) => mux_out_5_49_port, 
                           A(48) => mux_out_5_48_port, A(47) => 
                           mux_out_5_47_port, A(46) => mux_out_5_46_port, A(45)
                           => mux_out_5_45_port, A(44) => mux_out_5_44_port, 
                           A(43) => mux_out_5_43_port, A(42) => 
                           mux_out_5_42_port, A(41) => mux_out_5_41_port, A(40)
                           => mux_out_5_40_port, A(39) => mux_out_5_39_port, 
                           A(38) => mux_out_5_38_port, A(37) => 
                           mux_out_5_37_port, A(36) => mux_out_5_36_port, A(35)
                           => mux_out_5_35_port, A(34) => mux_out_5_34_port, 
                           A(33) => mux_out_5_33_port, A(32) => 
                           mux_out_5_32_port, A(31) => mux_out_5_31_port, A(30)
                           => mux_out_5_30_port, A(29) => mux_out_5_29_port, 
                           A(28) => mux_out_5_28_port, A(27) => 
                           mux_out_5_27_port, A(26) => mux_out_5_26_port, A(25)
                           => mux_out_5_25_port, A(24) => mux_out_5_24_port, 
                           A(23) => mux_out_5_23_port, A(22) => 
                           mux_out_5_22_port, A(21) => mux_out_5_21_port, A(20)
                           => mux_out_5_20_port, A(19) => mux_out_5_19_port, 
                           A(18) => mux_out_5_18_port, A(17) => 
                           mux_out_5_17_port, A(16) => mux_out_5_16_port, A(15)
                           => mux_out_5_15_port, A(14) => mux_out_5_14_port, 
                           A(13) => mux_out_5_13_port, A(12) => 
                           mux_out_5_12_port, A(11) => mux_out_5_11_port, A(10)
                           => mux_out_5_10_port, A(9) => mux_out_5_9_port, A(8)
                           => mux_out_5_8_port, A(7) => mux_out_5_7_port, A(6) 
                           => mux_out_5_6_port, A(5) => mux_out_5_5_port, A(4) 
                           => mux_out_5_4_port, A(3) => mux_out_5_3_port, A(2) 
                           => mux_out_5_2_port, A(1) => mux_out_5_1_port, A(0) 
                           => mux_out_5_0_port, B(63) => add_in_4_63_port, 
                           B(62) => add_in_4_62_port, B(61) => add_in_4_61_port
                           , B(60) => add_in_4_60_port, B(59) => 
                           add_in_4_59_port, B(58) => add_in_4_58_port, B(57) 
                           => add_in_4_57_port, B(56) => add_in_4_56_port, 
                           B(55) => add_in_4_55_port, B(54) => add_in_4_54_port
                           , B(53) => add_in_4_53_port, B(52) => 
                           add_in_4_52_port, B(51) => add_in_4_51_port, B(50) 
                           => add_in_4_50_port, B(49) => add_in_4_49_port, 
                           B(48) => add_in_4_48_port, B(47) => add_in_4_47_port
                           , B(46) => add_in_4_46_port, B(45) => 
                           add_in_4_45_port, B(44) => add_in_4_44_port, B(43) 
                           => add_in_4_43_port, B(42) => add_in_4_42_port, 
                           B(41) => add_in_4_41_port, B(40) => add_in_4_40_port
                           , B(39) => add_in_4_39_port, B(38) => 
                           add_in_4_38_port, B(37) => add_in_4_37_port, B(36) 
                           => add_in_4_36_port, B(35) => add_in_4_35_port, 
                           B(34) => add_in_4_34_port, B(33) => add_in_4_33_port
                           , B(32) => add_in_4_32_port, B(31) => 
                           add_in_4_31_port, B(30) => add_in_4_30_port, B(29) 
                           => add_in_4_29_port, B(28) => add_in_4_28_port, 
                           B(27) => add_in_4_27_port, B(26) => add_in_4_26_port
                           , B(25) => add_in_4_25_port, B(24) => 
                           add_in_4_24_port, B(23) => add_in_4_23_port, B(22) 
                           => add_in_4_22_port, B(21) => add_in_4_21_port, 
                           B(20) => add_in_4_20_port, B(19) => add_in_4_19_port
                           , B(18) => add_in_4_18_port, B(17) => 
                           add_in_4_17_port, B(16) => add_in_4_16_port, B(15) 
                           => add_in_4_15_port, B(14) => add_in_4_14_port, 
                           B(13) => add_in_4_13_port, B(12) => add_in_4_12_port
                           , B(11) => add_in_4_11_port, B(10) => 
                           add_in_4_10_port, B(9) => add_in_4_9_port, B(8) => 
                           add_in_4_8_port, B(7) => add_in_4_7_port, B(6) => 
                           add_in_4_6_port, B(5) => add_in_4_5_port, B(4) => 
                           add_in_4_4_port, B(3) => add_in_4_3_port, B(2) => 
                           add_in_4_2_port, B(1) => add_in_4_1_port, B(0) => 
                           add_in_4_0_port, Ci => mode_4_port, S(63) => 
                           add_in_5_63_port, S(62) => add_in_5_62_port, S(61) 
                           => add_in_5_61_port, S(60) => add_in_5_60_port, 
                           S(59) => add_in_5_59_port, S(58) => add_in_5_58_port
                           , S(57) => add_in_5_57_port, S(56) => 
                           add_in_5_56_port, S(55) => add_in_5_55_port, S(54) 
                           => add_in_5_54_port, S(53) => add_in_5_53_port, 
                           S(52) => add_in_5_52_port, S(51) => add_in_5_51_port
                           , S(50) => add_in_5_50_port, S(49) => 
                           add_in_5_49_port, S(48) => add_in_5_48_port, S(47) 
                           => add_in_5_47_port, S(46) => add_in_5_46_port, 
                           S(45) => add_in_5_45_port, S(44) => add_in_5_44_port
                           , S(43) => add_in_5_43_port, S(42) => 
                           add_in_5_42_port, S(41) => add_in_5_41_port, S(40) 
                           => add_in_5_40_port, S(39) => add_in_5_39_port, 
                           S(38) => add_in_5_38_port, S(37) => add_in_5_37_port
                           , S(36) => add_in_5_36_port, S(35) => 
                           add_in_5_35_port, S(34) => add_in_5_34_port, S(33) 
                           => add_in_5_33_port, S(32) => add_in_5_32_port, 
                           S(31) => add_in_5_31_port, S(30) => add_in_5_30_port
                           , S(29) => add_in_5_29_port, S(28) => 
                           add_in_5_28_port, S(27) => add_in_5_27_port, S(26) 
                           => add_in_5_26_port, S(25) => add_in_5_25_port, 
                           S(24) => add_in_5_24_port, S(23) => add_in_5_23_port
                           , S(22) => add_in_5_22_port, S(21) => 
                           add_in_5_21_port, S(20) => add_in_5_20_port, S(19) 
                           => add_in_5_19_port, S(18) => add_in_5_18_port, 
                           S(17) => add_in_5_17_port, S(16) => add_in_5_16_port
                           , S(15) => add_in_5_15_port, S(14) => 
                           add_in_5_14_port, S(13) => add_in_5_13_port, S(12) 
                           => add_in_5_12_port, S(11) => add_in_5_11_port, 
                           S(10) => add_in_5_10_port, S(9) => add_in_5_9_port, 
                           S(8) => add_in_5_8_port, S(7) => add_in_5_7_port, 
                           S(6) => add_in_5_6_port, S(5) => add_in_5_5_port, 
                           S(4) => add_in_5_4_port, S(3) => add_in_5_3_port, 
                           S(2) => add_in_5_2_port, S(1) => add_in_5_1_port, 
                           S(0) => add_in_5_0_port, Co => net21316);
   add_i_5 : RCA_generic_N64_10 port map( A(63) => mux_out_6_63_port, A(62) => 
                           mux_out_6_62_port, A(61) => mux_out_6_61_port, A(60)
                           => mux_out_6_60_port, A(59) => mux_out_6_59_port, 
                           A(58) => mux_out_6_58_port, A(57) => 
                           mux_out_6_57_port, A(56) => mux_out_6_56_port, A(55)
                           => mux_out_6_55_port, A(54) => mux_out_6_54_port, 
                           A(53) => mux_out_6_53_port, A(52) => 
                           mux_out_6_52_port, A(51) => mux_out_6_51_port, A(50)
                           => mux_out_6_50_port, A(49) => mux_out_6_49_port, 
                           A(48) => mux_out_6_48_port, A(47) => 
                           mux_out_6_47_port, A(46) => mux_out_6_46_port, A(45)
                           => mux_out_6_45_port, A(44) => mux_out_6_44_port, 
                           A(43) => mux_out_6_43_port, A(42) => 
                           mux_out_6_42_port, A(41) => mux_out_6_41_port, A(40)
                           => mux_out_6_40_port, A(39) => mux_out_6_39_port, 
                           A(38) => mux_out_6_38_port, A(37) => 
                           mux_out_6_37_port, A(36) => mux_out_6_36_port, A(35)
                           => mux_out_6_35_port, A(34) => mux_out_6_34_port, 
                           A(33) => mux_out_6_33_port, A(32) => 
                           mux_out_6_32_port, A(31) => mux_out_6_31_port, A(30)
                           => mux_out_6_30_port, A(29) => mux_out_6_29_port, 
                           A(28) => mux_out_6_28_port, A(27) => 
                           mux_out_6_27_port, A(26) => mux_out_6_26_port, A(25)
                           => mux_out_6_25_port, A(24) => mux_out_6_24_port, 
                           A(23) => mux_out_6_23_port, A(22) => 
                           mux_out_6_22_port, A(21) => mux_out_6_21_port, A(20)
                           => mux_out_6_20_port, A(19) => mux_out_6_19_port, 
                           A(18) => mux_out_6_18_port, A(17) => 
                           mux_out_6_17_port, A(16) => mux_out_6_16_port, A(15)
                           => mux_out_6_15_port, A(14) => mux_out_6_14_port, 
                           A(13) => mux_out_6_13_port, A(12) => 
                           mux_out_6_12_port, A(11) => mux_out_6_11_port, A(10)
                           => mux_out_6_10_port, A(9) => mux_out_6_9_port, A(8)
                           => mux_out_6_8_port, A(7) => mux_out_6_7_port, A(6) 
                           => mux_out_6_6_port, A(5) => mux_out_6_5_port, A(4) 
                           => mux_out_6_4_port, A(3) => mux_out_6_3_port, A(2) 
                           => mux_out_6_2_port, A(1) => mux_out_6_1_port, A(0) 
                           => mux_out_6_0_port, B(63) => add_in_5_63_port, 
                           B(62) => add_in_5_62_port, B(61) => add_in_5_61_port
                           , B(60) => add_in_5_60_port, B(59) => 
                           add_in_5_59_port, B(58) => add_in_5_58_port, B(57) 
                           => add_in_5_57_port, B(56) => add_in_5_56_port, 
                           B(55) => add_in_5_55_port, B(54) => add_in_5_54_port
                           , B(53) => add_in_5_53_port, B(52) => 
                           add_in_5_52_port, B(51) => add_in_5_51_port, B(50) 
                           => add_in_5_50_port, B(49) => add_in_5_49_port, 
                           B(48) => add_in_5_48_port, B(47) => add_in_5_47_port
                           , B(46) => add_in_5_46_port, B(45) => 
                           add_in_5_45_port, B(44) => add_in_5_44_port, B(43) 
                           => add_in_5_43_port, B(42) => add_in_5_42_port, 
                           B(41) => add_in_5_41_port, B(40) => add_in_5_40_port
                           , B(39) => add_in_5_39_port, B(38) => 
                           add_in_5_38_port, B(37) => add_in_5_37_port, B(36) 
                           => add_in_5_36_port, B(35) => add_in_5_35_port, 
                           B(34) => add_in_5_34_port, B(33) => add_in_5_33_port
                           , B(32) => add_in_5_32_port, B(31) => 
                           add_in_5_31_port, B(30) => add_in_5_30_port, B(29) 
                           => add_in_5_29_port, B(28) => add_in_5_28_port, 
                           B(27) => add_in_5_27_port, B(26) => add_in_5_26_port
                           , B(25) => add_in_5_25_port, B(24) => 
                           add_in_5_24_port, B(23) => add_in_5_23_port, B(22) 
                           => add_in_5_22_port, B(21) => add_in_5_21_port, 
                           B(20) => add_in_5_20_port, B(19) => add_in_5_19_port
                           , B(18) => add_in_5_18_port, B(17) => 
                           add_in_5_17_port, B(16) => add_in_5_16_port, B(15) 
                           => add_in_5_15_port, B(14) => add_in_5_14_port, 
                           B(13) => add_in_5_13_port, B(12) => add_in_5_12_port
                           , B(11) => add_in_5_11_port, B(10) => 
                           add_in_5_10_port, B(9) => add_in_5_9_port, B(8) => 
                           add_in_5_8_port, B(7) => add_in_5_7_port, B(6) => 
                           add_in_5_6_port, B(5) => add_in_5_5_port, B(4) => 
                           add_in_5_4_port, B(3) => add_in_5_3_port, B(2) => 
                           add_in_5_2_port, B(1) => add_in_5_1_port, B(0) => 
                           add_in_5_0_port, Ci => mode_5_port, S(63) => 
                           add_in_6_63_port, S(62) => add_in_6_62_port, S(61) 
                           => add_in_6_61_port, S(60) => add_in_6_60_port, 
                           S(59) => add_in_6_59_port, S(58) => add_in_6_58_port
                           , S(57) => add_in_6_57_port, S(56) => 
                           add_in_6_56_port, S(55) => add_in_6_55_port, S(54) 
                           => add_in_6_54_port, S(53) => add_in_6_53_port, 
                           S(52) => add_in_6_52_port, S(51) => add_in_6_51_port
                           , S(50) => add_in_6_50_port, S(49) => 
                           add_in_6_49_port, S(48) => add_in_6_48_port, S(47) 
                           => add_in_6_47_port, S(46) => add_in_6_46_port, 
                           S(45) => add_in_6_45_port, S(44) => add_in_6_44_port
                           , S(43) => add_in_6_43_port, S(42) => 
                           add_in_6_42_port, S(41) => add_in_6_41_port, S(40) 
                           => add_in_6_40_port, S(39) => add_in_6_39_port, 
                           S(38) => add_in_6_38_port, S(37) => add_in_6_37_port
                           , S(36) => add_in_6_36_port, S(35) => 
                           add_in_6_35_port, S(34) => add_in_6_34_port, S(33) 
                           => add_in_6_33_port, S(32) => add_in_6_32_port, 
                           S(31) => add_in_6_31_port, S(30) => add_in_6_30_port
                           , S(29) => add_in_6_29_port, S(28) => 
                           add_in_6_28_port, S(27) => add_in_6_27_port, S(26) 
                           => add_in_6_26_port, S(25) => add_in_6_25_port, 
                           S(24) => add_in_6_24_port, S(23) => add_in_6_23_port
                           , S(22) => add_in_6_22_port, S(21) => 
                           add_in_6_21_port, S(20) => add_in_6_20_port, S(19) 
                           => add_in_6_19_port, S(18) => add_in_6_18_port, 
                           S(17) => add_in_6_17_port, S(16) => add_in_6_16_port
                           , S(15) => add_in_6_15_port, S(14) => 
                           add_in_6_14_port, S(13) => add_in_6_13_port, S(12) 
                           => add_in_6_12_port, S(11) => add_in_6_11_port, 
                           S(10) => add_in_6_10_port, S(9) => add_in_6_9_port, 
                           S(8) => add_in_6_8_port, S(7) => add_in_6_7_port, 
                           S(6) => add_in_6_6_port, S(5) => add_in_6_5_port, 
                           S(4) => add_in_6_4_port, S(3) => add_in_6_3_port, 
                           S(2) => add_in_6_2_port, S(1) => add_in_6_1_port, 
                           S(0) => add_in_6_0_port, Co => net21315);
   add_i_6 : RCA_generic_N64_9 port map( A(63) => mux_out_7_63_port, A(62) => 
                           mux_out_7_62_port, A(61) => mux_out_7_61_port, A(60)
                           => mux_out_7_60_port, A(59) => mux_out_7_59_port, 
                           A(58) => mux_out_7_58_port, A(57) => 
                           mux_out_7_57_port, A(56) => mux_out_7_56_port, A(55)
                           => mux_out_7_55_port, A(54) => mux_out_7_54_port, 
                           A(53) => mux_out_7_53_port, A(52) => 
                           mux_out_7_52_port, A(51) => mux_out_7_51_port, A(50)
                           => mux_out_7_50_port, A(49) => mux_out_7_49_port, 
                           A(48) => mux_out_7_48_port, A(47) => 
                           mux_out_7_47_port, A(46) => mux_out_7_46_port, A(45)
                           => mux_out_7_45_port, A(44) => mux_out_7_44_port, 
                           A(43) => mux_out_7_43_port, A(42) => 
                           mux_out_7_42_port, A(41) => mux_out_7_41_port, A(40)
                           => mux_out_7_40_port, A(39) => mux_out_7_39_port, 
                           A(38) => mux_out_7_38_port, A(37) => 
                           mux_out_7_37_port, A(36) => mux_out_7_36_port, A(35)
                           => mux_out_7_35_port, A(34) => mux_out_7_34_port, 
                           A(33) => mux_out_7_33_port, A(32) => 
                           mux_out_7_32_port, A(31) => mux_out_7_31_port, A(30)
                           => mux_out_7_30_port, A(29) => mux_out_7_29_port, 
                           A(28) => mux_out_7_28_port, A(27) => 
                           mux_out_7_27_port, A(26) => mux_out_7_26_port, A(25)
                           => mux_out_7_25_port, A(24) => mux_out_7_24_port, 
                           A(23) => mux_out_7_23_port, A(22) => 
                           mux_out_7_22_port, A(21) => mux_out_7_21_port, A(20)
                           => mux_out_7_20_port, A(19) => mux_out_7_19_port, 
                           A(18) => mux_out_7_18_port, A(17) => 
                           mux_out_7_17_port, A(16) => mux_out_7_16_port, A(15)
                           => mux_out_7_15_port, A(14) => mux_out_7_14_port, 
                           A(13) => mux_out_7_13_port, A(12) => 
                           mux_out_7_12_port, A(11) => mux_out_7_11_port, A(10)
                           => mux_out_7_10_port, A(9) => mux_out_7_9_port, A(8)
                           => mux_out_7_8_port, A(7) => mux_out_7_7_port, A(6) 
                           => mux_out_7_6_port, A(5) => mux_out_7_5_port, A(4) 
                           => mux_out_7_4_port, A(3) => mux_out_7_3_port, A(2) 
                           => mux_out_7_2_port, A(1) => mux_out_7_1_port, A(0) 
                           => mux_out_7_0_port, B(63) => add_in_6_63_port, 
                           B(62) => add_in_6_62_port, B(61) => add_in_6_61_port
                           , B(60) => add_in_6_60_port, B(59) => 
                           add_in_6_59_port, B(58) => add_in_6_58_port, B(57) 
                           => add_in_6_57_port, B(56) => add_in_6_56_port, 
                           B(55) => add_in_6_55_port, B(54) => add_in_6_54_port
                           , B(53) => add_in_6_53_port, B(52) => 
                           add_in_6_52_port, B(51) => add_in_6_51_port, B(50) 
                           => add_in_6_50_port, B(49) => add_in_6_49_port, 
                           B(48) => add_in_6_48_port, B(47) => add_in_6_47_port
                           , B(46) => add_in_6_46_port, B(45) => 
                           add_in_6_45_port, B(44) => add_in_6_44_port, B(43) 
                           => add_in_6_43_port, B(42) => add_in_6_42_port, 
                           B(41) => add_in_6_41_port, B(40) => add_in_6_40_port
                           , B(39) => add_in_6_39_port, B(38) => 
                           add_in_6_38_port, B(37) => add_in_6_37_port, B(36) 
                           => add_in_6_36_port, B(35) => add_in_6_35_port, 
                           B(34) => add_in_6_34_port, B(33) => add_in_6_33_port
                           , B(32) => add_in_6_32_port, B(31) => 
                           add_in_6_31_port, B(30) => add_in_6_30_port, B(29) 
                           => add_in_6_29_port, B(28) => add_in_6_28_port, 
                           B(27) => add_in_6_27_port, B(26) => add_in_6_26_port
                           , B(25) => add_in_6_25_port, B(24) => 
                           add_in_6_24_port, B(23) => add_in_6_23_port, B(22) 
                           => add_in_6_22_port, B(21) => add_in_6_21_port, 
                           B(20) => add_in_6_20_port, B(19) => add_in_6_19_port
                           , B(18) => add_in_6_18_port, B(17) => 
                           add_in_6_17_port, B(16) => add_in_6_16_port, B(15) 
                           => add_in_6_15_port, B(14) => add_in_6_14_port, 
                           B(13) => add_in_6_13_port, B(12) => add_in_6_12_port
                           , B(11) => add_in_6_11_port, B(10) => 
                           add_in_6_10_port, B(9) => add_in_6_9_port, B(8) => 
                           add_in_6_8_port, B(7) => add_in_6_7_port, B(6) => 
                           add_in_6_6_port, B(5) => add_in_6_5_port, B(4) => 
                           add_in_6_4_port, B(3) => add_in_6_3_port, B(2) => 
                           add_in_6_2_port, B(1) => add_in_6_1_port, B(0) => 
                           add_in_6_0_port, Ci => mode_6_port, S(63) => 
                           add_in_7_63_port, S(62) => add_in_7_62_port, S(61) 
                           => add_in_7_61_port, S(60) => add_in_7_60_port, 
                           S(59) => add_in_7_59_port, S(58) => add_in_7_58_port
                           , S(57) => add_in_7_57_port, S(56) => 
                           add_in_7_56_port, S(55) => add_in_7_55_port, S(54) 
                           => add_in_7_54_port, S(53) => add_in_7_53_port, 
                           S(52) => add_in_7_52_port, S(51) => add_in_7_51_port
                           , S(50) => add_in_7_50_port, S(49) => 
                           add_in_7_49_port, S(48) => add_in_7_48_port, S(47) 
                           => add_in_7_47_port, S(46) => add_in_7_46_port, 
                           S(45) => add_in_7_45_port, S(44) => add_in_7_44_port
                           , S(43) => add_in_7_43_port, S(42) => 
                           add_in_7_42_port, S(41) => add_in_7_41_port, S(40) 
                           => add_in_7_40_port, S(39) => add_in_7_39_port, 
                           S(38) => add_in_7_38_port, S(37) => add_in_7_37_port
                           , S(36) => add_in_7_36_port, S(35) => 
                           add_in_7_35_port, S(34) => add_in_7_34_port, S(33) 
                           => add_in_7_33_port, S(32) => add_in_7_32_port, 
                           S(31) => add_in_7_31_port, S(30) => add_in_7_30_port
                           , S(29) => add_in_7_29_port, S(28) => 
                           add_in_7_28_port, S(27) => add_in_7_27_port, S(26) 
                           => add_in_7_26_port, S(25) => add_in_7_25_port, 
                           S(24) => add_in_7_24_port, S(23) => add_in_7_23_port
                           , S(22) => add_in_7_22_port, S(21) => 
                           add_in_7_21_port, S(20) => add_in_7_20_port, S(19) 
                           => add_in_7_19_port, S(18) => add_in_7_18_port, 
                           S(17) => add_in_7_17_port, S(16) => add_in_7_16_port
                           , S(15) => add_in_7_15_port, S(14) => 
                           add_in_7_14_port, S(13) => add_in_7_13_port, S(12) 
                           => add_in_7_12_port, S(11) => add_in_7_11_port, 
                           S(10) => add_in_7_10_port, S(9) => add_in_7_9_port, 
                           S(8) => add_in_7_8_port, S(7) => add_in_7_7_port, 
                           S(6) => add_in_7_6_port, S(5) => add_in_7_5_port, 
                           S(4) => add_in_7_4_port, S(3) => add_in_7_3_port, 
                           S(2) => add_in_7_2_port, S(1) => add_in_7_1_port, 
                           S(0) => add_in_7_0_port, Co => net21314);
   add_i_7 : RCA_generic_N64_8 port map( A(63) => mux_out_8_63_port, A(62) => 
                           mux_out_8_62_port, A(61) => mux_out_8_61_port, A(60)
                           => mux_out_8_60_port, A(59) => mux_out_8_59_port, 
                           A(58) => mux_out_8_58_port, A(57) => 
                           mux_out_8_57_port, A(56) => mux_out_8_56_port, A(55)
                           => mux_out_8_55_port, A(54) => mux_out_8_54_port, 
                           A(53) => mux_out_8_53_port, A(52) => 
                           mux_out_8_52_port, A(51) => mux_out_8_51_port, A(50)
                           => mux_out_8_50_port, A(49) => mux_out_8_49_port, 
                           A(48) => mux_out_8_48_port, A(47) => 
                           mux_out_8_47_port, A(46) => mux_out_8_46_port, A(45)
                           => mux_out_8_45_port, A(44) => mux_out_8_44_port, 
                           A(43) => mux_out_8_43_port, A(42) => 
                           mux_out_8_42_port, A(41) => mux_out_8_41_port, A(40)
                           => mux_out_8_40_port, A(39) => mux_out_8_39_port, 
                           A(38) => mux_out_8_38_port, A(37) => 
                           mux_out_8_37_port, A(36) => mux_out_8_36_port, A(35)
                           => mux_out_8_35_port, A(34) => mux_out_8_34_port, 
                           A(33) => mux_out_8_33_port, A(32) => 
                           mux_out_8_32_port, A(31) => mux_out_8_31_port, A(30)
                           => mux_out_8_30_port, A(29) => mux_out_8_29_port, 
                           A(28) => mux_out_8_28_port, A(27) => 
                           mux_out_8_27_port, A(26) => mux_out_8_26_port, A(25)
                           => mux_out_8_25_port, A(24) => mux_out_8_24_port, 
                           A(23) => mux_out_8_23_port, A(22) => 
                           mux_out_8_22_port, A(21) => mux_out_8_21_port, A(20)
                           => mux_out_8_20_port, A(19) => mux_out_8_19_port, 
                           A(18) => mux_out_8_18_port, A(17) => 
                           mux_out_8_17_port, A(16) => mux_out_8_16_port, A(15)
                           => mux_out_8_15_port, A(14) => mux_out_8_14_port, 
                           A(13) => mux_out_8_13_port, A(12) => 
                           mux_out_8_12_port, A(11) => mux_out_8_11_port, A(10)
                           => mux_out_8_10_port, A(9) => mux_out_8_9_port, A(8)
                           => mux_out_8_8_port, A(7) => mux_out_8_7_port, A(6) 
                           => mux_out_8_6_port, A(5) => mux_out_8_5_port, A(4) 
                           => mux_out_8_4_port, A(3) => mux_out_8_3_port, A(2) 
                           => mux_out_8_2_port, A(1) => mux_out_8_1_port, A(0) 
                           => mux_out_8_0_port, B(63) => add_in_7_63_port, 
                           B(62) => add_in_7_62_port, B(61) => add_in_7_61_port
                           , B(60) => add_in_7_60_port, B(59) => 
                           add_in_7_59_port, B(58) => add_in_7_58_port, B(57) 
                           => add_in_7_57_port, B(56) => add_in_7_56_port, 
                           B(55) => add_in_7_55_port, B(54) => add_in_7_54_port
                           , B(53) => add_in_7_53_port, B(52) => 
                           add_in_7_52_port, B(51) => add_in_7_51_port, B(50) 
                           => add_in_7_50_port, B(49) => add_in_7_49_port, 
                           B(48) => add_in_7_48_port, B(47) => add_in_7_47_port
                           , B(46) => add_in_7_46_port, B(45) => 
                           add_in_7_45_port, B(44) => add_in_7_44_port, B(43) 
                           => add_in_7_43_port, B(42) => add_in_7_42_port, 
                           B(41) => add_in_7_41_port, B(40) => add_in_7_40_port
                           , B(39) => add_in_7_39_port, B(38) => 
                           add_in_7_38_port, B(37) => add_in_7_37_port, B(36) 
                           => add_in_7_36_port, B(35) => add_in_7_35_port, 
                           B(34) => add_in_7_34_port, B(33) => add_in_7_33_port
                           , B(32) => add_in_7_32_port, B(31) => 
                           add_in_7_31_port, B(30) => add_in_7_30_port, B(29) 
                           => add_in_7_29_port, B(28) => add_in_7_28_port, 
                           B(27) => add_in_7_27_port, B(26) => add_in_7_26_port
                           , B(25) => add_in_7_25_port, B(24) => 
                           add_in_7_24_port, B(23) => add_in_7_23_port, B(22) 
                           => add_in_7_22_port, B(21) => add_in_7_21_port, 
                           B(20) => add_in_7_20_port, B(19) => add_in_7_19_port
                           , B(18) => add_in_7_18_port, B(17) => 
                           add_in_7_17_port, B(16) => add_in_7_16_port, B(15) 
                           => add_in_7_15_port, B(14) => add_in_7_14_port, 
                           B(13) => add_in_7_13_port, B(12) => add_in_7_12_port
                           , B(11) => add_in_7_11_port, B(10) => 
                           add_in_7_10_port, B(9) => add_in_7_9_port, B(8) => 
                           add_in_7_8_port, B(7) => add_in_7_7_port, B(6) => 
                           add_in_7_6_port, B(5) => add_in_7_5_port, B(4) => 
                           add_in_7_4_port, B(3) => add_in_7_3_port, B(2) => 
                           add_in_7_2_port, B(1) => add_in_7_1_port, B(0) => 
                           add_in_7_0_port, Ci => mode_7_port, S(63) => 
                           add_in_8_63_port, S(62) => add_in_8_62_port, S(61) 
                           => add_in_8_61_port, S(60) => add_in_8_60_port, 
                           S(59) => add_in_8_59_port, S(58) => add_in_8_58_port
                           , S(57) => add_in_8_57_port, S(56) => 
                           add_in_8_56_port, S(55) => add_in_8_55_port, S(54) 
                           => add_in_8_54_port, S(53) => add_in_8_53_port, 
                           S(52) => add_in_8_52_port, S(51) => add_in_8_51_port
                           , S(50) => add_in_8_50_port, S(49) => 
                           add_in_8_49_port, S(48) => add_in_8_48_port, S(47) 
                           => add_in_8_47_port, S(46) => add_in_8_46_port, 
                           S(45) => add_in_8_45_port, S(44) => add_in_8_44_port
                           , S(43) => add_in_8_43_port, S(42) => 
                           add_in_8_42_port, S(41) => add_in_8_41_port, S(40) 
                           => add_in_8_40_port, S(39) => add_in_8_39_port, 
                           S(38) => add_in_8_38_port, S(37) => add_in_8_37_port
                           , S(36) => add_in_8_36_port, S(35) => 
                           add_in_8_35_port, S(34) => add_in_8_34_port, S(33) 
                           => add_in_8_33_port, S(32) => add_in_8_32_port, 
                           S(31) => add_in_8_31_port, S(30) => add_in_8_30_port
                           , S(29) => add_in_8_29_port, S(28) => 
                           add_in_8_28_port, S(27) => add_in_8_27_port, S(26) 
                           => add_in_8_26_port, S(25) => add_in_8_25_port, 
                           S(24) => add_in_8_24_port, S(23) => add_in_8_23_port
                           , S(22) => add_in_8_22_port, S(21) => 
                           add_in_8_21_port, S(20) => add_in_8_20_port, S(19) 
                           => add_in_8_19_port, S(18) => add_in_8_18_port, 
                           S(17) => add_in_8_17_port, S(16) => add_in_8_16_port
                           , S(15) => add_in_8_15_port, S(14) => 
                           add_in_8_14_port, S(13) => add_in_8_13_port, S(12) 
                           => add_in_8_12_port, S(11) => add_in_8_11_port, 
                           S(10) => add_in_8_10_port, S(9) => add_in_8_9_port, 
                           S(8) => add_in_8_8_port, S(7) => add_in_8_7_port, 
                           S(6) => add_in_8_6_port, S(5) => add_in_8_5_port, 
                           S(4) => add_in_8_4_port, S(3) => add_in_8_3_port, 
                           S(2) => add_in_8_2_port, S(1) => add_in_8_1_port, 
                           S(0) => add_in_8_0_port, Co => net21313);
   add_i_8 : RCA_generic_N64_7 port map( A(63) => mux_out_9_63_port, A(62) => 
                           mux_out_9_62_port, A(61) => mux_out_9_61_port, A(60)
                           => mux_out_9_60_port, A(59) => mux_out_9_59_port, 
                           A(58) => mux_out_9_58_port, A(57) => 
                           mux_out_9_57_port, A(56) => mux_out_9_56_port, A(55)
                           => mux_out_9_55_port, A(54) => mux_out_9_54_port, 
                           A(53) => mux_out_9_53_port, A(52) => 
                           mux_out_9_52_port, A(51) => mux_out_9_51_port, A(50)
                           => mux_out_9_50_port, A(49) => mux_out_9_49_port, 
                           A(48) => mux_out_9_48_port, A(47) => 
                           mux_out_9_47_port, A(46) => mux_out_9_46_port, A(45)
                           => mux_out_9_45_port, A(44) => mux_out_9_44_port, 
                           A(43) => mux_out_9_43_port, A(42) => 
                           mux_out_9_42_port, A(41) => mux_out_9_41_port, A(40)
                           => mux_out_9_40_port, A(39) => mux_out_9_39_port, 
                           A(38) => mux_out_9_38_port, A(37) => 
                           mux_out_9_37_port, A(36) => mux_out_9_36_port, A(35)
                           => mux_out_9_35_port, A(34) => mux_out_9_34_port, 
                           A(33) => mux_out_9_33_port, A(32) => 
                           mux_out_9_32_port, A(31) => mux_out_9_31_port, A(30)
                           => mux_out_9_30_port, A(29) => mux_out_9_29_port, 
                           A(28) => mux_out_9_28_port, A(27) => 
                           mux_out_9_27_port, A(26) => mux_out_9_26_port, A(25)
                           => mux_out_9_25_port, A(24) => mux_out_9_24_port, 
                           A(23) => mux_out_9_23_port, A(22) => 
                           mux_out_9_22_port, A(21) => mux_out_9_21_port, A(20)
                           => mux_out_9_20_port, A(19) => mux_out_9_19_port, 
                           A(18) => mux_out_9_18_port, A(17) => 
                           mux_out_9_17_port, A(16) => mux_out_9_16_port, A(15)
                           => mux_out_9_15_port, A(14) => mux_out_9_14_port, 
                           A(13) => mux_out_9_13_port, A(12) => 
                           mux_out_9_12_port, A(11) => mux_out_9_11_port, A(10)
                           => mux_out_9_10_port, A(9) => mux_out_9_9_port, A(8)
                           => mux_out_9_8_port, A(7) => mux_out_9_7_port, A(6) 
                           => mux_out_9_6_port, A(5) => mux_out_9_5_port, A(4) 
                           => mux_out_9_4_port, A(3) => mux_out_9_3_port, A(2) 
                           => mux_out_9_2_port, A(1) => mux_out_9_1_port, A(0) 
                           => mux_out_9_0_port, B(63) => add_in_8_63_port, 
                           B(62) => add_in_8_62_port, B(61) => add_in_8_61_port
                           , B(60) => add_in_8_60_port, B(59) => 
                           add_in_8_59_port, B(58) => add_in_8_58_port, B(57) 
                           => add_in_8_57_port, B(56) => add_in_8_56_port, 
                           B(55) => add_in_8_55_port, B(54) => add_in_8_54_port
                           , B(53) => add_in_8_53_port, B(52) => 
                           add_in_8_52_port, B(51) => add_in_8_51_port, B(50) 
                           => add_in_8_50_port, B(49) => add_in_8_49_port, 
                           B(48) => add_in_8_48_port, B(47) => add_in_8_47_port
                           , B(46) => add_in_8_46_port, B(45) => 
                           add_in_8_45_port, B(44) => add_in_8_44_port, B(43) 
                           => add_in_8_43_port, B(42) => add_in_8_42_port, 
                           B(41) => add_in_8_41_port, B(40) => add_in_8_40_port
                           , B(39) => add_in_8_39_port, B(38) => 
                           add_in_8_38_port, B(37) => add_in_8_37_port, B(36) 
                           => add_in_8_36_port, B(35) => add_in_8_35_port, 
                           B(34) => add_in_8_34_port, B(33) => add_in_8_33_port
                           , B(32) => add_in_8_32_port, B(31) => 
                           add_in_8_31_port, B(30) => add_in_8_30_port, B(29) 
                           => add_in_8_29_port, B(28) => add_in_8_28_port, 
                           B(27) => add_in_8_27_port, B(26) => add_in_8_26_port
                           , B(25) => add_in_8_25_port, B(24) => 
                           add_in_8_24_port, B(23) => add_in_8_23_port, B(22) 
                           => add_in_8_22_port, B(21) => add_in_8_21_port, 
                           B(20) => add_in_8_20_port, B(19) => add_in_8_19_port
                           , B(18) => add_in_8_18_port, B(17) => 
                           add_in_8_17_port, B(16) => add_in_8_16_port, B(15) 
                           => add_in_8_15_port, B(14) => add_in_8_14_port, 
                           B(13) => add_in_8_13_port, B(12) => add_in_8_12_port
                           , B(11) => add_in_8_11_port, B(10) => 
                           add_in_8_10_port, B(9) => add_in_8_9_port, B(8) => 
                           add_in_8_8_port, B(7) => add_in_8_7_port, B(6) => 
                           add_in_8_6_port, B(5) => add_in_8_5_port, B(4) => 
                           add_in_8_4_port, B(3) => add_in_8_3_port, B(2) => 
                           add_in_8_2_port, B(1) => add_in_8_1_port, B(0) => 
                           add_in_8_0_port, Ci => mode_8_port, S(63) => 
                           add_in_9_63_port, S(62) => add_in_9_62_port, S(61) 
                           => add_in_9_61_port, S(60) => add_in_9_60_port, 
                           S(59) => add_in_9_59_port, S(58) => add_in_9_58_port
                           , S(57) => add_in_9_57_port, S(56) => 
                           add_in_9_56_port, S(55) => add_in_9_55_port, S(54) 
                           => add_in_9_54_port, S(53) => add_in_9_53_port, 
                           S(52) => add_in_9_52_port, S(51) => add_in_9_51_port
                           , S(50) => add_in_9_50_port, S(49) => 
                           add_in_9_49_port, S(48) => add_in_9_48_port, S(47) 
                           => add_in_9_47_port, S(46) => add_in_9_46_port, 
                           S(45) => add_in_9_45_port, S(44) => add_in_9_44_port
                           , S(43) => add_in_9_43_port, S(42) => 
                           add_in_9_42_port, S(41) => add_in_9_41_port, S(40) 
                           => add_in_9_40_port, S(39) => add_in_9_39_port, 
                           S(38) => add_in_9_38_port, S(37) => add_in_9_37_port
                           , S(36) => add_in_9_36_port, S(35) => 
                           add_in_9_35_port, S(34) => add_in_9_34_port, S(33) 
                           => add_in_9_33_port, S(32) => add_in_9_32_port, 
                           S(31) => add_in_9_31_port, S(30) => add_in_9_30_port
                           , S(29) => add_in_9_29_port, S(28) => 
                           add_in_9_28_port, S(27) => add_in_9_27_port, S(26) 
                           => add_in_9_26_port, S(25) => add_in_9_25_port, 
                           S(24) => add_in_9_24_port, S(23) => add_in_9_23_port
                           , S(22) => add_in_9_22_port, S(21) => 
                           add_in_9_21_port, S(20) => add_in_9_20_port, S(19) 
                           => add_in_9_19_port, S(18) => add_in_9_18_port, 
                           S(17) => add_in_9_17_port, S(16) => add_in_9_16_port
                           , S(15) => add_in_9_15_port, S(14) => 
                           add_in_9_14_port, S(13) => add_in_9_13_port, S(12) 
                           => add_in_9_12_port, S(11) => add_in_9_11_port, 
                           S(10) => add_in_9_10_port, S(9) => add_in_9_9_port, 
                           S(8) => add_in_9_8_port, S(7) => add_in_9_7_port, 
                           S(6) => add_in_9_6_port, S(5) => add_in_9_5_port, 
                           S(4) => add_in_9_4_port, S(3) => add_in_9_3_port, 
                           S(2) => add_in_9_2_port, S(1) => add_in_9_1_port, 
                           S(0) => add_in_9_0_port, Co => net21312);
   add_i_9 : RCA_generic_N64_6 port map( A(63) => mux_out_10_63_port, A(62) => 
                           mux_out_10_62_port, A(61) => mux_out_10_61_port, 
                           A(60) => mux_out_10_60_port, A(59) => 
                           mux_out_10_59_port, A(58) => mux_out_10_58_port, 
                           A(57) => mux_out_10_57_port, A(56) => 
                           mux_out_10_56_port, A(55) => mux_out_10_55_port, 
                           A(54) => mux_out_10_54_port, A(53) => 
                           mux_out_10_53_port, A(52) => mux_out_10_52_port, 
                           A(51) => mux_out_10_51_port, A(50) => 
                           mux_out_10_50_port, A(49) => mux_out_10_49_port, 
                           A(48) => mux_out_10_48_port, A(47) => 
                           mux_out_10_47_port, A(46) => mux_out_10_46_port, 
                           A(45) => mux_out_10_45_port, A(44) => 
                           mux_out_10_44_port, A(43) => mux_out_10_43_port, 
                           A(42) => mux_out_10_42_port, A(41) => 
                           mux_out_10_41_port, A(40) => mux_out_10_40_port, 
                           A(39) => mux_out_10_39_port, A(38) => 
                           mux_out_10_38_port, A(37) => mux_out_10_37_port, 
                           A(36) => mux_out_10_36_port, A(35) => 
                           mux_out_10_35_port, A(34) => mux_out_10_34_port, 
                           A(33) => mux_out_10_33_port, A(32) => 
                           mux_out_10_32_port, A(31) => mux_out_10_31_port, 
                           A(30) => mux_out_10_30_port, A(29) => 
                           mux_out_10_29_port, A(28) => mux_out_10_28_port, 
                           A(27) => mux_out_10_27_port, A(26) => 
                           mux_out_10_26_port, A(25) => mux_out_10_25_port, 
                           A(24) => mux_out_10_24_port, A(23) => 
                           mux_out_10_23_port, A(22) => mux_out_10_22_port, 
                           A(21) => mux_out_10_21_port, A(20) => 
                           mux_out_10_20_port, A(19) => mux_out_10_19_port, 
                           A(18) => mux_out_10_18_port, A(17) => 
                           mux_out_10_17_port, A(16) => mux_out_10_16_port, 
                           A(15) => mux_out_10_15_port, A(14) => 
                           mux_out_10_14_port, A(13) => mux_out_10_13_port, 
                           A(12) => mux_out_10_12_port, A(11) => 
                           mux_out_10_11_port, A(10) => mux_out_10_10_port, 
                           A(9) => mux_out_10_9_port, A(8) => mux_out_10_8_port
                           , A(7) => mux_out_10_7_port, A(6) => 
                           mux_out_10_6_port, A(5) => mux_out_10_5_port, A(4) 
                           => mux_out_10_4_port, A(3) => mux_out_10_3_port, 
                           A(2) => mux_out_10_2_port, A(1) => mux_out_10_1_port
                           , A(0) => mux_out_10_0_port, B(63) => 
                           add_in_9_63_port, B(62) => add_in_9_62_port, B(61) 
                           => add_in_9_61_port, B(60) => add_in_9_60_port, 
                           B(59) => add_in_9_59_port, B(58) => add_in_9_58_port
                           , B(57) => add_in_9_57_port, B(56) => 
                           add_in_9_56_port, B(55) => add_in_9_55_port, B(54) 
                           => add_in_9_54_port, B(53) => add_in_9_53_port, 
                           B(52) => add_in_9_52_port, B(51) => add_in_9_51_port
                           , B(50) => add_in_9_50_port, B(49) => 
                           add_in_9_49_port, B(48) => add_in_9_48_port, B(47) 
                           => add_in_9_47_port, B(46) => add_in_9_46_port, 
                           B(45) => add_in_9_45_port, B(44) => add_in_9_44_port
                           , B(43) => add_in_9_43_port, B(42) => 
                           add_in_9_42_port, B(41) => add_in_9_41_port, B(40) 
                           => add_in_9_40_port, B(39) => add_in_9_39_port, 
                           B(38) => add_in_9_38_port, B(37) => add_in_9_37_port
                           , B(36) => add_in_9_36_port, B(35) => 
                           add_in_9_35_port, B(34) => add_in_9_34_port, B(33) 
                           => add_in_9_33_port, B(32) => add_in_9_32_port, 
                           B(31) => add_in_9_31_port, B(30) => add_in_9_30_port
                           , B(29) => add_in_9_29_port, B(28) => 
                           add_in_9_28_port, B(27) => add_in_9_27_port, B(26) 
                           => add_in_9_26_port, B(25) => add_in_9_25_port, 
                           B(24) => add_in_9_24_port, B(23) => add_in_9_23_port
                           , B(22) => add_in_9_22_port, B(21) => 
                           add_in_9_21_port, B(20) => add_in_9_20_port, B(19) 
                           => add_in_9_19_port, B(18) => add_in_9_18_port, 
                           B(17) => add_in_9_17_port, B(16) => add_in_9_16_port
                           , B(15) => add_in_9_15_port, B(14) => 
                           add_in_9_14_port, B(13) => add_in_9_13_port, B(12) 
                           => add_in_9_12_port, B(11) => add_in_9_11_port, 
                           B(10) => add_in_9_10_port, B(9) => add_in_9_9_port, 
                           B(8) => add_in_9_8_port, B(7) => add_in_9_7_port, 
                           B(6) => add_in_9_6_port, B(5) => add_in_9_5_port, 
                           B(4) => add_in_9_4_port, B(3) => add_in_9_3_port, 
                           B(2) => add_in_9_2_port, B(1) => add_in_9_1_port, 
                           B(0) => add_in_9_0_port, Ci => mode_9_port, S(63) =>
                           add_in_10_63_port, S(62) => add_in_10_62_port, S(61)
                           => add_in_10_61_port, S(60) => add_in_10_60_port, 
                           S(59) => add_in_10_59_port, S(58) => 
                           add_in_10_58_port, S(57) => add_in_10_57_port, S(56)
                           => add_in_10_56_port, S(55) => add_in_10_55_port, 
                           S(54) => add_in_10_54_port, S(53) => 
                           add_in_10_53_port, S(52) => add_in_10_52_port, S(51)
                           => add_in_10_51_port, S(50) => add_in_10_50_port, 
                           S(49) => add_in_10_49_port, S(48) => 
                           add_in_10_48_port, S(47) => add_in_10_47_port, S(46)
                           => add_in_10_46_port, S(45) => add_in_10_45_port, 
                           S(44) => add_in_10_44_port, S(43) => 
                           add_in_10_43_port, S(42) => add_in_10_42_port, S(41)
                           => add_in_10_41_port, S(40) => add_in_10_40_port, 
                           S(39) => add_in_10_39_port, S(38) => 
                           add_in_10_38_port, S(37) => add_in_10_37_port, S(36)
                           => add_in_10_36_port, S(35) => add_in_10_35_port, 
                           S(34) => add_in_10_34_port, S(33) => 
                           add_in_10_33_port, S(32) => add_in_10_32_port, S(31)
                           => add_in_10_31_port, S(30) => add_in_10_30_port, 
                           S(29) => add_in_10_29_port, S(28) => 
                           add_in_10_28_port, S(27) => add_in_10_27_port, S(26)
                           => add_in_10_26_port, S(25) => add_in_10_25_port, 
                           S(24) => add_in_10_24_port, S(23) => 
                           add_in_10_23_port, S(22) => add_in_10_22_port, S(21)
                           => add_in_10_21_port, S(20) => add_in_10_20_port, 
                           S(19) => add_in_10_19_port, S(18) => 
                           add_in_10_18_port, S(17) => add_in_10_17_port, S(16)
                           => add_in_10_16_port, S(15) => add_in_10_15_port, 
                           S(14) => add_in_10_14_port, S(13) => 
                           add_in_10_13_port, S(12) => add_in_10_12_port, S(11)
                           => add_in_10_11_port, S(10) => add_in_10_10_port, 
                           S(9) => add_in_10_9_port, S(8) => add_in_10_8_port, 
                           S(7) => add_in_10_7_port, S(6) => add_in_10_6_port, 
                           S(5) => add_in_10_5_port, S(4) => add_in_10_4_port, 
                           S(3) => add_in_10_3_port, S(2) => add_in_10_2_port, 
                           S(1) => add_in_10_1_port, S(0) => add_in_10_0_port, 
                           Co => net21311);
   add_i_10 : RCA_generic_N64_5 port map( A(63) => mux_out_11_63_port, A(62) =>
                           mux_out_11_62_port, A(61) => mux_out_11_61_port, 
                           A(60) => mux_out_11_60_port, A(59) => 
                           mux_out_11_59_port, A(58) => mux_out_11_58_port, 
                           A(57) => mux_out_11_57_port, A(56) => 
                           mux_out_11_56_port, A(55) => mux_out_11_55_port, 
                           A(54) => mux_out_11_54_port, A(53) => 
                           mux_out_11_53_port, A(52) => mux_out_11_52_port, 
                           A(51) => mux_out_11_51_port, A(50) => 
                           mux_out_11_50_port, A(49) => mux_out_11_49_port, 
                           A(48) => mux_out_11_48_port, A(47) => 
                           mux_out_11_47_port, A(46) => mux_out_11_46_port, 
                           A(45) => mux_out_11_45_port, A(44) => 
                           mux_out_11_44_port, A(43) => mux_out_11_43_port, 
                           A(42) => mux_out_11_42_port, A(41) => 
                           mux_out_11_41_port, A(40) => mux_out_11_40_port, 
                           A(39) => mux_out_11_39_port, A(38) => 
                           mux_out_11_38_port, A(37) => mux_out_11_37_port, 
                           A(36) => mux_out_11_36_port, A(35) => 
                           mux_out_11_35_port, A(34) => mux_out_11_34_port, 
                           A(33) => mux_out_11_33_port, A(32) => 
                           mux_out_11_32_port, A(31) => mux_out_11_31_port, 
                           A(30) => mux_out_11_30_port, A(29) => 
                           mux_out_11_29_port, A(28) => mux_out_11_28_port, 
                           A(27) => mux_out_11_27_port, A(26) => 
                           mux_out_11_26_port, A(25) => mux_out_11_25_port, 
                           A(24) => mux_out_11_24_port, A(23) => 
                           mux_out_11_23_port, A(22) => mux_out_11_22_port, 
                           A(21) => mux_out_11_21_port, A(20) => 
                           mux_out_11_20_port, A(19) => mux_out_11_19_port, 
                           A(18) => mux_out_11_18_port, A(17) => 
                           mux_out_11_17_port, A(16) => mux_out_11_16_port, 
                           A(15) => mux_out_11_15_port, A(14) => 
                           mux_out_11_14_port, A(13) => mux_out_11_13_port, 
                           A(12) => mux_out_11_12_port, A(11) => 
                           mux_out_11_11_port, A(10) => mux_out_11_10_port, 
                           A(9) => mux_out_11_9_port, A(8) => mux_out_11_8_port
                           , A(7) => mux_out_11_7_port, A(6) => 
                           mux_out_11_6_port, A(5) => mux_out_11_5_port, A(4) 
                           => mux_out_11_4_port, A(3) => mux_out_11_3_port, 
                           A(2) => mux_out_11_2_port, A(1) => mux_out_11_1_port
                           , A(0) => mux_out_11_0_port, B(63) => 
                           add_in_10_63_port, B(62) => add_in_10_62_port, B(61)
                           => add_in_10_61_port, B(60) => add_in_10_60_port, 
                           B(59) => add_in_10_59_port, B(58) => 
                           add_in_10_58_port, B(57) => add_in_10_57_port, B(56)
                           => add_in_10_56_port, B(55) => add_in_10_55_port, 
                           B(54) => add_in_10_54_port, B(53) => 
                           add_in_10_53_port, B(52) => add_in_10_52_port, B(51)
                           => add_in_10_51_port, B(50) => add_in_10_50_port, 
                           B(49) => add_in_10_49_port, B(48) => 
                           add_in_10_48_port, B(47) => add_in_10_47_port, B(46)
                           => add_in_10_46_port, B(45) => add_in_10_45_port, 
                           B(44) => add_in_10_44_port, B(43) => 
                           add_in_10_43_port, B(42) => add_in_10_42_port, B(41)
                           => add_in_10_41_port, B(40) => add_in_10_40_port, 
                           B(39) => add_in_10_39_port, B(38) => 
                           add_in_10_38_port, B(37) => add_in_10_37_port, B(36)
                           => add_in_10_36_port, B(35) => add_in_10_35_port, 
                           B(34) => add_in_10_34_port, B(33) => 
                           add_in_10_33_port, B(32) => add_in_10_32_port, B(31)
                           => add_in_10_31_port, B(30) => add_in_10_30_port, 
                           B(29) => add_in_10_29_port, B(28) => 
                           add_in_10_28_port, B(27) => add_in_10_27_port, B(26)
                           => add_in_10_26_port, B(25) => add_in_10_25_port, 
                           B(24) => add_in_10_24_port, B(23) => 
                           add_in_10_23_port, B(22) => add_in_10_22_port, B(21)
                           => add_in_10_21_port, B(20) => add_in_10_20_port, 
                           B(19) => add_in_10_19_port, B(18) => 
                           add_in_10_18_port, B(17) => add_in_10_17_port, B(16)
                           => add_in_10_16_port, B(15) => add_in_10_15_port, 
                           B(14) => add_in_10_14_port, B(13) => 
                           add_in_10_13_port, B(12) => add_in_10_12_port, B(11)
                           => add_in_10_11_port, B(10) => add_in_10_10_port, 
                           B(9) => add_in_10_9_port, B(8) => add_in_10_8_port, 
                           B(7) => add_in_10_7_port, B(6) => add_in_10_6_port, 
                           B(5) => add_in_10_5_port, B(4) => add_in_10_4_port, 
                           B(3) => add_in_10_3_port, B(2) => add_in_10_2_port, 
                           B(1) => add_in_10_1_port, B(0) => add_in_10_0_port, 
                           Ci => mode_10_port, S(63) => add_in_11_63_port, 
                           S(62) => add_in_11_62_port, S(61) => 
                           add_in_11_61_port, S(60) => add_in_11_60_port, S(59)
                           => add_in_11_59_port, S(58) => add_in_11_58_port, 
                           S(57) => add_in_11_57_port, S(56) => 
                           add_in_11_56_port, S(55) => add_in_11_55_port, S(54)
                           => add_in_11_54_port, S(53) => add_in_11_53_port, 
                           S(52) => add_in_11_52_port, S(51) => 
                           add_in_11_51_port, S(50) => add_in_11_50_port, S(49)
                           => add_in_11_49_port, S(48) => add_in_11_48_port, 
                           S(47) => add_in_11_47_port, S(46) => 
                           add_in_11_46_port, S(45) => add_in_11_45_port, S(44)
                           => add_in_11_44_port, S(43) => add_in_11_43_port, 
                           S(42) => add_in_11_42_port, S(41) => 
                           add_in_11_41_port, S(40) => add_in_11_40_port, S(39)
                           => add_in_11_39_port, S(38) => add_in_11_38_port, 
                           S(37) => add_in_11_37_port, S(36) => 
                           add_in_11_36_port, S(35) => add_in_11_35_port, S(34)
                           => add_in_11_34_port, S(33) => add_in_11_33_port, 
                           S(32) => add_in_11_32_port, S(31) => 
                           add_in_11_31_port, S(30) => add_in_11_30_port, S(29)
                           => add_in_11_29_port, S(28) => add_in_11_28_port, 
                           S(27) => add_in_11_27_port, S(26) => 
                           add_in_11_26_port, S(25) => add_in_11_25_port, S(24)
                           => add_in_11_24_port, S(23) => add_in_11_23_port, 
                           S(22) => add_in_11_22_port, S(21) => 
                           add_in_11_21_port, S(20) => add_in_11_20_port, S(19)
                           => add_in_11_19_port, S(18) => add_in_11_18_port, 
                           S(17) => add_in_11_17_port, S(16) => 
                           add_in_11_16_port, S(15) => add_in_11_15_port, S(14)
                           => add_in_11_14_port, S(13) => add_in_11_13_port, 
                           S(12) => add_in_11_12_port, S(11) => 
                           add_in_11_11_port, S(10) => add_in_11_10_port, S(9) 
                           => add_in_11_9_port, S(8) => add_in_11_8_port, S(7) 
                           => add_in_11_7_port, S(6) => add_in_11_6_port, S(5) 
                           => add_in_11_5_port, S(4) => add_in_11_4_port, S(3) 
                           => add_in_11_3_port, S(2) => add_in_11_2_port, S(1) 
                           => add_in_11_1_port, S(0) => add_in_11_0_port, Co =>
                           net21310);
   add_i_11 : RCA_generic_N64_4 port map( A(63) => mux_out_12_63_port, A(62) =>
                           mux_out_12_62_port, A(61) => mux_out_12_61_port, 
                           A(60) => mux_out_12_60_port, A(59) => 
                           mux_out_12_59_port, A(58) => mux_out_12_58_port, 
                           A(57) => mux_out_12_57_port, A(56) => 
                           mux_out_12_56_port, A(55) => mux_out_12_55_port, 
                           A(54) => mux_out_12_54_port, A(53) => 
                           mux_out_12_53_port, A(52) => mux_out_12_52_port, 
                           A(51) => mux_out_12_51_port, A(50) => 
                           mux_out_12_50_port, A(49) => mux_out_12_49_port, 
                           A(48) => mux_out_12_48_port, A(47) => 
                           mux_out_12_47_port, A(46) => mux_out_12_46_port, 
                           A(45) => mux_out_12_45_port, A(44) => 
                           mux_out_12_44_port, A(43) => mux_out_12_43_port, 
                           A(42) => mux_out_12_42_port, A(41) => 
                           mux_out_12_41_port, A(40) => mux_out_12_40_port, 
                           A(39) => mux_out_12_39_port, A(38) => 
                           mux_out_12_38_port, A(37) => mux_out_12_37_port, 
                           A(36) => mux_out_12_36_port, A(35) => 
                           mux_out_12_35_port, A(34) => mux_out_12_34_port, 
                           A(33) => mux_out_12_33_port, A(32) => 
                           mux_out_12_32_port, A(31) => mux_out_12_31_port, 
                           A(30) => mux_out_12_30_port, A(29) => 
                           mux_out_12_29_port, A(28) => mux_out_12_28_port, 
                           A(27) => mux_out_12_27_port, A(26) => 
                           mux_out_12_26_port, A(25) => mux_out_12_25_port, 
                           A(24) => mux_out_12_24_port, A(23) => 
                           mux_out_12_23_port, A(22) => mux_out_12_22_port, 
                           A(21) => mux_out_12_21_port, A(20) => 
                           mux_out_12_20_port, A(19) => mux_out_12_19_port, 
                           A(18) => mux_out_12_18_port, A(17) => 
                           mux_out_12_17_port, A(16) => mux_out_12_16_port, 
                           A(15) => mux_out_12_15_port, A(14) => 
                           mux_out_12_14_port, A(13) => mux_out_12_13_port, 
                           A(12) => mux_out_12_12_port, A(11) => 
                           mux_out_12_11_port, A(10) => mux_out_12_10_port, 
                           A(9) => mux_out_12_9_port, A(8) => mux_out_12_8_port
                           , A(7) => mux_out_12_7_port, A(6) => 
                           mux_out_12_6_port, A(5) => mux_out_12_5_port, A(4) 
                           => mux_out_12_4_port, A(3) => mux_out_12_3_port, 
                           A(2) => mux_out_12_2_port, A(1) => mux_out_12_1_port
                           , A(0) => mux_out_12_0_port, B(63) => 
                           add_in_11_63_port, B(62) => add_in_11_62_port, B(61)
                           => add_in_11_61_port, B(60) => add_in_11_60_port, 
                           B(59) => add_in_11_59_port, B(58) => 
                           add_in_11_58_port, B(57) => add_in_11_57_port, B(56)
                           => add_in_11_56_port, B(55) => add_in_11_55_port, 
                           B(54) => add_in_11_54_port, B(53) => 
                           add_in_11_53_port, B(52) => add_in_11_52_port, B(51)
                           => add_in_11_51_port, B(50) => add_in_11_50_port, 
                           B(49) => add_in_11_49_port, B(48) => 
                           add_in_11_48_port, B(47) => add_in_11_47_port, B(46)
                           => add_in_11_46_port, B(45) => add_in_11_45_port, 
                           B(44) => add_in_11_44_port, B(43) => 
                           add_in_11_43_port, B(42) => add_in_11_42_port, B(41)
                           => add_in_11_41_port, B(40) => add_in_11_40_port, 
                           B(39) => add_in_11_39_port, B(38) => 
                           add_in_11_38_port, B(37) => add_in_11_37_port, B(36)
                           => add_in_11_36_port, B(35) => add_in_11_35_port, 
                           B(34) => add_in_11_34_port, B(33) => 
                           add_in_11_33_port, B(32) => add_in_11_32_port, B(31)
                           => add_in_11_31_port, B(30) => add_in_11_30_port, 
                           B(29) => add_in_11_29_port, B(28) => 
                           add_in_11_28_port, B(27) => add_in_11_27_port, B(26)
                           => add_in_11_26_port, B(25) => add_in_11_25_port, 
                           B(24) => add_in_11_24_port, B(23) => 
                           add_in_11_23_port, B(22) => add_in_11_22_port, B(21)
                           => add_in_11_21_port, B(20) => add_in_11_20_port, 
                           B(19) => add_in_11_19_port, B(18) => 
                           add_in_11_18_port, B(17) => add_in_11_17_port, B(16)
                           => add_in_11_16_port, B(15) => add_in_11_15_port, 
                           B(14) => add_in_11_14_port, B(13) => 
                           add_in_11_13_port, B(12) => add_in_11_12_port, B(11)
                           => add_in_11_11_port, B(10) => add_in_11_10_port, 
                           B(9) => add_in_11_9_port, B(8) => add_in_11_8_port, 
                           B(7) => add_in_11_7_port, B(6) => add_in_11_6_port, 
                           B(5) => add_in_11_5_port, B(4) => add_in_11_4_port, 
                           B(3) => add_in_11_3_port, B(2) => add_in_11_2_port, 
                           B(1) => add_in_11_1_port, B(0) => add_in_11_0_port, 
                           Ci => mode_11_port, S(63) => add_in_12_63_port, 
                           S(62) => add_in_12_62_port, S(61) => 
                           add_in_12_61_port, S(60) => add_in_12_60_port, S(59)
                           => add_in_12_59_port, S(58) => add_in_12_58_port, 
                           S(57) => add_in_12_57_port, S(56) => 
                           add_in_12_56_port, S(55) => add_in_12_55_port, S(54)
                           => add_in_12_54_port, S(53) => add_in_12_53_port, 
                           S(52) => add_in_12_52_port, S(51) => 
                           add_in_12_51_port, S(50) => add_in_12_50_port, S(49)
                           => add_in_12_49_port, S(48) => add_in_12_48_port, 
                           S(47) => add_in_12_47_port, S(46) => 
                           add_in_12_46_port, S(45) => add_in_12_45_port, S(44)
                           => add_in_12_44_port, S(43) => add_in_12_43_port, 
                           S(42) => add_in_12_42_port, S(41) => 
                           add_in_12_41_port, S(40) => add_in_12_40_port, S(39)
                           => add_in_12_39_port, S(38) => add_in_12_38_port, 
                           S(37) => add_in_12_37_port, S(36) => 
                           add_in_12_36_port, S(35) => add_in_12_35_port, S(34)
                           => add_in_12_34_port, S(33) => add_in_12_33_port, 
                           S(32) => add_in_12_32_port, S(31) => 
                           add_in_12_31_port, S(30) => add_in_12_30_port, S(29)
                           => add_in_12_29_port, S(28) => add_in_12_28_port, 
                           S(27) => add_in_12_27_port, S(26) => 
                           add_in_12_26_port, S(25) => add_in_12_25_port, S(24)
                           => add_in_12_24_port, S(23) => add_in_12_23_port, 
                           S(22) => add_in_12_22_port, S(21) => 
                           add_in_12_21_port, S(20) => add_in_12_20_port, S(19)
                           => add_in_12_19_port, S(18) => add_in_12_18_port, 
                           S(17) => add_in_12_17_port, S(16) => 
                           add_in_12_16_port, S(15) => add_in_12_15_port, S(14)
                           => add_in_12_14_port, S(13) => add_in_12_13_port, 
                           S(12) => add_in_12_12_port, S(11) => 
                           add_in_12_11_port, S(10) => add_in_12_10_port, S(9) 
                           => add_in_12_9_port, S(8) => add_in_12_8_port, S(7) 
                           => add_in_12_7_port, S(6) => add_in_12_6_port, S(5) 
                           => add_in_12_5_port, S(4) => add_in_12_4_port, S(3) 
                           => add_in_12_3_port, S(2) => add_in_12_2_port, S(1) 
                           => add_in_12_1_port, S(0) => add_in_12_0_port, Co =>
                           net21309);
   add_i_12 : RCA_generic_N64_3 port map( A(63) => mux_out_13_63_port, A(62) =>
                           mux_out_13_62_port, A(61) => mux_out_13_61_port, 
                           A(60) => mux_out_13_60_port, A(59) => 
                           mux_out_13_59_port, A(58) => mux_out_13_58_port, 
                           A(57) => mux_out_13_57_port, A(56) => 
                           mux_out_13_56_port, A(55) => mux_out_13_55_port, 
                           A(54) => mux_out_13_54_port, A(53) => 
                           mux_out_13_53_port, A(52) => mux_out_13_52_port, 
                           A(51) => mux_out_13_51_port, A(50) => 
                           mux_out_13_50_port, A(49) => mux_out_13_49_port, 
                           A(48) => mux_out_13_48_port, A(47) => 
                           mux_out_13_47_port, A(46) => mux_out_13_46_port, 
                           A(45) => mux_out_13_45_port, A(44) => 
                           mux_out_13_44_port, A(43) => mux_out_13_43_port, 
                           A(42) => mux_out_13_42_port, A(41) => 
                           mux_out_13_41_port, A(40) => mux_out_13_40_port, 
                           A(39) => mux_out_13_39_port, A(38) => 
                           mux_out_13_38_port, A(37) => mux_out_13_37_port, 
                           A(36) => mux_out_13_36_port, A(35) => 
                           mux_out_13_35_port, A(34) => mux_out_13_34_port, 
                           A(33) => mux_out_13_33_port, A(32) => 
                           mux_out_13_32_port, A(31) => mux_out_13_31_port, 
                           A(30) => mux_out_13_30_port, A(29) => 
                           mux_out_13_29_port, A(28) => mux_out_13_28_port, 
                           A(27) => mux_out_13_27_port, A(26) => 
                           mux_out_13_26_port, A(25) => mux_out_13_25_port, 
                           A(24) => mux_out_13_24_port, A(23) => 
                           mux_out_13_23_port, A(22) => mux_out_13_22_port, 
                           A(21) => mux_out_13_21_port, A(20) => 
                           mux_out_13_20_port, A(19) => mux_out_13_19_port, 
                           A(18) => mux_out_13_18_port, A(17) => 
                           mux_out_13_17_port, A(16) => mux_out_13_16_port, 
                           A(15) => mux_out_13_15_port, A(14) => 
                           mux_out_13_14_port, A(13) => mux_out_13_13_port, 
                           A(12) => mux_out_13_12_port, A(11) => 
                           mux_out_13_11_port, A(10) => mux_out_13_10_port, 
                           A(9) => mux_out_13_9_port, A(8) => mux_out_13_8_port
                           , A(7) => mux_out_13_7_port, A(6) => 
                           mux_out_13_6_port, A(5) => mux_out_13_5_port, A(4) 
                           => mux_out_13_4_port, A(3) => mux_out_13_3_port, 
                           A(2) => mux_out_13_2_port, A(1) => mux_out_13_1_port
                           , A(0) => mux_out_13_0_port, B(63) => 
                           add_in_12_63_port, B(62) => add_in_12_62_port, B(61)
                           => add_in_12_61_port, B(60) => add_in_12_60_port, 
                           B(59) => add_in_12_59_port, B(58) => 
                           add_in_12_58_port, B(57) => add_in_12_57_port, B(56)
                           => add_in_12_56_port, B(55) => add_in_12_55_port, 
                           B(54) => add_in_12_54_port, B(53) => 
                           add_in_12_53_port, B(52) => add_in_12_52_port, B(51)
                           => add_in_12_51_port, B(50) => add_in_12_50_port, 
                           B(49) => add_in_12_49_port, B(48) => 
                           add_in_12_48_port, B(47) => add_in_12_47_port, B(46)
                           => add_in_12_46_port, B(45) => add_in_12_45_port, 
                           B(44) => add_in_12_44_port, B(43) => 
                           add_in_12_43_port, B(42) => add_in_12_42_port, B(41)
                           => add_in_12_41_port, B(40) => add_in_12_40_port, 
                           B(39) => add_in_12_39_port, B(38) => 
                           add_in_12_38_port, B(37) => add_in_12_37_port, B(36)
                           => add_in_12_36_port, B(35) => add_in_12_35_port, 
                           B(34) => add_in_12_34_port, B(33) => 
                           add_in_12_33_port, B(32) => add_in_12_32_port, B(31)
                           => add_in_12_31_port, B(30) => add_in_12_30_port, 
                           B(29) => add_in_12_29_port, B(28) => 
                           add_in_12_28_port, B(27) => add_in_12_27_port, B(26)
                           => add_in_12_26_port, B(25) => add_in_12_25_port, 
                           B(24) => add_in_12_24_port, B(23) => 
                           add_in_12_23_port, B(22) => add_in_12_22_port, B(21)
                           => add_in_12_21_port, B(20) => add_in_12_20_port, 
                           B(19) => add_in_12_19_port, B(18) => 
                           add_in_12_18_port, B(17) => add_in_12_17_port, B(16)
                           => add_in_12_16_port, B(15) => add_in_12_15_port, 
                           B(14) => add_in_12_14_port, B(13) => 
                           add_in_12_13_port, B(12) => add_in_12_12_port, B(11)
                           => add_in_12_11_port, B(10) => add_in_12_10_port, 
                           B(9) => add_in_12_9_port, B(8) => add_in_12_8_port, 
                           B(7) => add_in_12_7_port, B(6) => add_in_12_6_port, 
                           B(5) => add_in_12_5_port, B(4) => add_in_12_4_port, 
                           B(3) => add_in_12_3_port, B(2) => add_in_12_2_port, 
                           B(1) => add_in_12_1_port, B(0) => add_in_12_0_port, 
                           Ci => mode_12_port, S(63) => add_in_13_63_port, 
                           S(62) => add_in_13_62_port, S(61) => 
                           add_in_13_61_port, S(60) => add_in_13_60_port, S(59)
                           => add_in_13_59_port, S(58) => add_in_13_58_port, 
                           S(57) => add_in_13_57_port, S(56) => 
                           add_in_13_56_port, S(55) => add_in_13_55_port, S(54)
                           => add_in_13_54_port, S(53) => add_in_13_53_port, 
                           S(52) => add_in_13_52_port, S(51) => 
                           add_in_13_51_port, S(50) => add_in_13_50_port, S(49)
                           => add_in_13_49_port, S(48) => add_in_13_48_port, 
                           S(47) => add_in_13_47_port, S(46) => 
                           add_in_13_46_port, S(45) => add_in_13_45_port, S(44)
                           => add_in_13_44_port, S(43) => add_in_13_43_port, 
                           S(42) => add_in_13_42_port, S(41) => 
                           add_in_13_41_port, S(40) => add_in_13_40_port, S(39)
                           => add_in_13_39_port, S(38) => add_in_13_38_port, 
                           S(37) => add_in_13_37_port, S(36) => 
                           add_in_13_36_port, S(35) => add_in_13_35_port, S(34)
                           => add_in_13_34_port, S(33) => add_in_13_33_port, 
                           S(32) => add_in_13_32_port, S(31) => 
                           add_in_13_31_port, S(30) => add_in_13_30_port, S(29)
                           => add_in_13_29_port, S(28) => add_in_13_28_port, 
                           S(27) => add_in_13_27_port, S(26) => 
                           add_in_13_26_port, S(25) => add_in_13_25_port, S(24)
                           => add_in_13_24_port, S(23) => add_in_13_23_port, 
                           S(22) => add_in_13_22_port, S(21) => 
                           add_in_13_21_port, S(20) => add_in_13_20_port, S(19)
                           => add_in_13_19_port, S(18) => add_in_13_18_port, 
                           S(17) => add_in_13_17_port, S(16) => 
                           add_in_13_16_port, S(15) => add_in_13_15_port, S(14)
                           => add_in_13_14_port, S(13) => add_in_13_13_port, 
                           S(12) => add_in_13_12_port, S(11) => 
                           add_in_13_11_port, S(10) => add_in_13_10_port, S(9) 
                           => add_in_13_9_port, S(8) => add_in_13_8_port, S(7) 
                           => add_in_13_7_port, S(6) => add_in_13_6_port, S(5) 
                           => add_in_13_5_port, S(4) => add_in_13_4_port, S(3) 
                           => add_in_13_3_port, S(2) => add_in_13_2_port, S(1) 
                           => add_in_13_1_port, S(0) => add_in_13_0_port, Co =>
                           net21308);
   add_i_13 : RCA_generic_N64_2 port map( A(63) => mux_out_14_63_port, A(62) =>
                           mux_out_14_62_port, A(61) => mux_out_14_61_port, 
                           A(60) => mux_out_14_60_port, A(59) => 
                           mux_out_14_59_port, A(58) => mux_out_14_58_port, 
                           A(57) => mux_out_14_57_port, A(56) => 
                           mux_out_14_56_port, A(55) => mux_out_14_55_port, 
                           A(54) => mux_out_14_54_port, A(53) => 
                           mux_out_14_53_port, A(52) => mux_out_14_52_port, 
                           A(51) => mux_out_14_51_port, A(50) => 
                           mux_out_14_50_port, A(49) => mux_out_14_49_port, 
                           A(48) => mux_out_14_48_port, A(47) => 
                           mux_out_14_47_port, A(46) => mux_out_14_46_port, 
                           A(45) => mux_out_14_45_port, A(44) => 
                           mux_out_14_44_port, A(43) => mux_out_14_43_port, 
                           A(42) => mux_out_14_42_port, A(41) => 
                           mux_out_14_41_port, A(40) => mux_out_14_40_port, 
                           A(39) => mux_out_14_39_port, A(38) => 
                           mux_out_14_38_port, A(37) => mux_out_14_37_port, 
                           A(36) => mux_out_14_36_port, A(35) => 
                           mux_out_14_35_port, A(34) => mux_out_14_34_port, 
                           A(33) => mux_out_14_33_port, A(32) => 
                           mux_out_14_32_port, A(31) => mux_out_14_31_port, 
                           A(30) => mux_out_14_30_port, A(29) => 
                           mux_out_14_29_port, A(28) => mux_out_14_28_port, 
                           A(27) => mux_out_14_27_port, A(26) => 
                           mux_out_14_26_port, A(25) => mux_out_14_25_port, 
                           A(24) => mux_out_14_24_port, A(23) => 
                           mux_out_14_23_port, A(22) => mux_out_14_22_port, 
                           A(21) => mux_out_14_21_port, A(20) => 
                           mux_out_14_20_port, A(19) => mux_out_14_19_port, 
                           A(18) => mux_out_14_18_port, A(17) => 
                           mux_out_14_17_port, A(16) => mux_out_14_16_port, 
                           A(15) => mux_out_14_15_port, A(14) => 
                           mux_out_14_14_port, A(13) => mux_out_14_13_port, 
                           A(12) => mux_out_14_12_port, A(11) => 
                           mux_out_14_11_port, A(10) => mux_out_14_10_port, 
                           A(9) => mux_out_14_9_port, A(8) => mux_out_14_8_port
                           , A(7) => mux_out_14_7_port, A(6) => 
                           mux_out_14_6_port, A(5) => mux_out_14_5_port, A(4) 
                           => mux_out_14_4_port, A(3) => mux_out_14_3_port, 
                           A(2) => mux_out_14_2_port, A(1) => mux_out_14_1_port
                           , A(0) => mux_out_14_0_port, B(63) => 
                           add_in_13_63_port, B(62) => add_in_13_62_port, B(61)
                           => add_in_13_61_port, B(60) => add_in_13_60_port, 
                           B(59) => add_in_13_59_port, B(58) => 
                           add_in_13_58_port, B(57) => add_in_13_57_port, B(56)
                           => add_in_13_56_port, B(55) => add_in_13_55_port, 
                           B(54) => add_in_13_54_port, B(53) => 
                           add_in_13_53_port, B(52) => add_in_13_52_port, B(51)
                           => add_in_13_51_port, B(50) => add_in_13_50_port, 
                           B(49) => add_in_13_49_port, B(48) => 
                           add_in_13_48_port, B(47) => add_in_13_47_port, B(46)
                           => add_in_13_46_port, B(45) => add_in_13_45_port, 
                           B(44) => add_in_13_44_port, B(43) => 
                           add_in_13_43_port, B(42) => add_in_13_42_port, B(41)
                           => add_in_13_41_port, B(40) => add_in_13_40_port, 
                           B(39) => add_in_13_39_port, B(38) => 
                           add_in_13_38_port, B(37) => add_in_13_37_port, B(36)
                           => add_in_13_36_port, B(35) => add_in_13_35_port, 
                           B(34) => add_in_13_34_port, B(33) => 
                           add_in_13_33_port, B(32) => add_in_13_32_port, B(31)
                           => add_in_13_31_port, B(30) => add_in_13_30_port, 
                           B(29) => add_in_13_29_port, B(28) => 
                           add_in_13_28_port, B(27) => add_in_13_27_port, B(26)
                           => add_in_13_26_port, B(25) => add_in_13_25_port, 
                           B(24) => add_in_13_24_port, B(23) => 
                           add_in_13_23_port, B(22) => add_in_13_22_port, B(21)
                           => add_in_13_21_port, B(20) => add_in_13_20_port, 
                           B(19) => add_in_13_19_port, B(18) => 
                           add_in_13_18_port, B(17) => add_in_13_17_port, B(16)
                           => add_in_13_16_port, B(15) => add_in_13_15_port, 
                           B(14) => add_in_13_14_port, B(13) => 
                           add_in_13_13_port, B(12) => add_in_13_12_port, B(11)
                           => add_in_13_11_port, B(10) => add_in_13_10_port, 
                           B(9) => add_in_13_9_port, B(8) => add_in_13_8_port, 
                           B(7) => add_in_13_7_port, B(6) => add_in_13_6_port, 
                           B(5) => add_in_13_5_port, B(4) => add_in_13_4_port, 
                           B(3) => add_in_13_3_port, B(2) => add_in_13_2_port, 
                           B(1) => add_in_13_1_port, B(0) => add_in_13_0_port, 
                           Ci => mode_13_port, S(63) => add_in_14_63_port, 
                           S(62) => add_in_14_62_port, S(61) => 
                           add_in_14_61_port, S(60) => add_in_14_60_port, S(59)
                           => add_in_14_59_port, S(58) => add_in_14_58_port, 
                           S(57) => add_in_14_57_port, S(56) => 
                           add_in_14_56_port, S(55) => add_in_14_55_port, S(54)
                           => add_in_14_54_port, S(53) => add_in_14_53_port, 
                           S(52) => add_in_14_52_port, S(51) => 
                           add_in_14_51_port, S(50) => add_in_14_50_port, S(49)
                           => add_in_14_49_port, S(48) => add_in_14_48_port, 
                           S(47) => add_in_14_47_port, S(46) => 
                           add_in_14_46_port, S(45) => add_in_14_45_port, S(44)
                           => add_in_14_44_port, S(43) => add_in_14_43_port, 
                           S(42) => add_in_14_42_port, S(41) => 
                           add_in_14_41_port, S(40) => add_in_14_40_port, S(39)
                           => add_in_14_39_port, S(38) => add_in_14_38_port, 
                           S(37) => add_in_14_37_port, S(36) => 
                           add_in_14_36_port, S(35) => add_in_14_35_port, S(34)
                           => add_in_14_34_port, S(33) => add_in_14_33_port, 
                           S(32) => add_in_14_32_port, S(31) => 
                           add_in_14_31_port, S(30) => add_in_14_30_port, S(29)
                           => add_in_14_29_port, S(28) => add_in_14_28_port, 
                           S(27) => add_in_14_27_port, S(26) => 
                           add_in_14_26_port, S(25) => add_in_14_25_port, S(24)
                           => add_in_14_24_port, S(23) => add_in_14_23_port, 
                           S(22) => add_in_14_22_port, S(21) => 
                           add_in_14_21_port, S(20) => add_in_14_20_port, S(19)
                           => add_in_14_19_port, S(18) => add_in_14_18_port, 
                           S(17) => add_in_14_17_port, S(16) => 
                           add_in_14_16_port, S(15) => add_in_14_15_port, S(14)
                           => add_in_14_14_port, S(13) => add_in_14_13_port, 
                           S(12) => add_in_14_12_port, S(11) => 
                           add_in_14_11_port, S(10) => add_in_14_10_port, S(9) 
                           => add_in_14_9_port, S(8) => add_in_14_8_port, S(7) 
                           => add_in_14_7_port, S(6) => add_in_14_6_port, S(5) 
                           => add_in_14_5_port, S(4) => add_in_14_4_port, S(3) 
                           => add_in_14_3_port, S(2) => add_in_14_2_port, S(1) 
                           => add_in_14_1_port, S(0) => add_in_14_0_port, Co =>
                           net21307);
   add_i_14 : RCA_generic_N64_1 port map( A(63) => mux_out_15_63_port, A(62) =>
                           mux_out_15_62_port, A(61) => mux_out_15_61_port, 
                           A(60) => mux_out_15_60_port, A(59) => 
                           mux_out_15_59_port, A(58) => mux_out_15_58_port, 
                           A(57) => mux_out_15_57_port, A(56) => 
                           mux_out_15_56_port, A(55) => mux_out_15_55_port, 
                           A(54) => mux_out_15_54_port, A(53) => 
                           mux_out_15_53_port, A(52) => mux_out_15_52_port, 
                           A(51) => mux_out_15_51_port, A(50) => 
                           mux_out_15_50_port, A(49) => mux_out_15_49_port, 
                           A(48) => mux_out_15_48_port, A(47) => 
                           mux_out_15_47_port, A(46) => mux_out_15_46_port, 
                           A(45) => mux_out_15_45_port, A(44) => 
                           mux_out_15_44_port, A(43) => mux_out_15_43_port, 
                           A(42) => mux_out_15_42_port, A(41) => 
                           mux_out_15_41_port, A(40) => mux_out_15_40_port, 
                           A(39) => mux_out_15_39_port, A(38) => 
                           mux_out_15_38_port, A(37) => mux_out_15_37_port, 
                           A(36) => mux_out_15_36_port, A(35) => 
                           mux_out_15_35_port, A(34) => mux_out_15_34_port, 
                           A(33) => mux_out_15_33_port, A(32) => 
                           mux_out_15_32_port, A(31) => mux_out_15_31_port, 
                           A(30) => mux_out_15_30_port, A(29) => 
                           mux_out_15_29_port, A(28) => mux_out_15_28_port, 
                           A(27) => mux_out_15_27_port, A(26) => 
                           mux_out_15_26_port, A(25) => mux_out_15_25_port, 
                           A(24) => mux_out_15_24_port, A(23) => 
                           mux_out_15_23_port, A(22) => mux_out_15_22_port, 
                           A(21) => mux_out_15_21_port, A(20) => 
                           mux_out_15_20_port, A(19) => mux_out_15_19_port, 
                           A(18) => mux_out_15_18_port, A(17) => 
                           mux_out_15_17_port, A(16) => mux_out_15_16_port, 
                           A(15) => mux_out_15_15_port, A(14) => 
                           mux_out_15_14_port, A(13) => mux_out_15_13_port, 
                           A(12) => mux_out_15_12_port, A(11) => 
                           mux_out_15_11_port, A(10) => mux_out_15_10_port, 
                           A(9) => mux_out_15_9_port, A(8) => mux_out_15_8_port
                           , A(7) => mux_out_15_7_port, A(6) => 
                           mux_out_15_6_port, A(5) => mux_out_15_5_port, A(4) 
                           => mux_out_15_4_port, A(3) => mux_out_15_3_port, 
                           A(2) => mux_out_15_2_port, A(1) => mux_out_15_1_port
                           , A(0) => mux_out_15_0_port, B(63) => 
                           add_in_14_63_port, B(62) => add_in_14_62_port, B(61)
                           => add_in_14_61_port, B(60) => add_in_14_60_port, 
                           B(59) => add_in_14_59_port, B(58) => 
                           add_in_14_58_port, B(57) => add_in_14_57_port, B(56)
                           => add_in_14_56_port, B(55) => add_in_14_55_port, 
                           B(54) => add_in_14_54_port, B(53) => 
                           add_in_14_53_port, B(52) => add_in_14_52_port, B(51)
                           => add_in_14_51_port, B(50) => add_in_14_50_port, 
                           B(49) => add_in_14_49_port, B(48) => 
                           add_in_14_48_port, B(47) => add_in_14_47_port, B(46)
                           => add_in_14_46_port, B(45) => add_in_14_45_port, 
                           B(44) => add_in_14_44_port, B(43) => 
                           add_in_14_43_port, B(42) => add_in_14_42_port, B(41)
                           => add_in_14_41_port, B(40) => add_in_14_40_port, 
                           B(39) => add_in_14_39_port, B(38) => 
                           add_in_14_38_port, B(37) => add_in_14_37_port, B(36)
                           => add_in_14_36_port, B(35) => add_in_14_35_port, 
                           B(34) => add_in_14_34_port, B(33) => 
                           add_in_14_33_port, B(32) => add_in_14_32_port, B(31)
                           => add_in_14_31_port, B(30) => add_in_14_30_port, 
                           B(29) => add_in_14_29_port, B(28) => 
                           add_in_14_28_port, B(27) => add_in_14_27_port, B(26)
                           => add_in_14_26_port, B(25) => add_in_14_25_port, 
                           B(24) => add_in_14_24_port, B(23) => 
                           add_in_14_23_port, B(22) => add_in_14_22_port, B(21)
                           => add_in_14_21_port, B(20) => add_in_14_20_port, 
                           B(19) => add_in_14_19_port, B(18) => 
                           add_in_14_18_port, B(17) => add_in_14_17_port, B(16)
                           => add_in_14_16_port, B(15) => add_in_14_15_port, 
                           B(14) => add_in_14_14_port, B(13) => 
                           add_in_14_13_port, B(12) => add_in_14_12_port, B(11)
                           => add_in_14_11_port, B(10) => add_in_14_10_port, 
                           B(9) => add_in_14_9_port, B(8) => add_in_14_8_port, 
                           B(7) => add_in_14_7_port, B(6) => add_in_14_6_port, 
                           B(5) => add_in_14_5_port, B(4) => add_in_14_4_port, 
                           B(3) => add_in_14_3_port, B(2) => add_in_14_2_port, 
                           B(1) => add_in_14_1_port, B(0) => add_in_14_0_port, 
                           Ci => mode_14_port, S(63) => add_in_15_63_port, 
                           S(62) => add_in_15_62_port, S(61) => 
                           add_in_15_61_port, S(60) => add_in_15_60_port, S(59)
                           => add_in_15_59_port, S(58) => add_in_15_58_port, 
                           S(57) => add_in_15_57_port, S(56) => 
                           add_in_15_56_port, S(55) => add_in_15_55_port, S(54)
                           => add_in_15_54_port, S(53) => add_in_15_53_port, 
                           S(52) => add_in_15_52_port, S(51) => 
                           add_in_15_51_port, S(50) => add_in_15_50_port, S(49)
                           => add_in_15_49_port, S(48) => add_in_15_48_port, 
                           S(47) => add_in_15_47_port, S(46) => 
                           add_in_15_46_port, S(45) => add_in_15_45_port, S(44)
                           => add_in_15_44_port, S(43) => add_in_15_43_port, 
                           S(42) => add_in_15_42_port, S(41) => 
                           add_in_15_41_port, S(40) => add_in_15_40_port, S(39)
                           => add_in_15_39_port, S(38) => add_in_15_38_port, 
                           S(37) => add_in_15_37_port, S(36) => 
                           add_in_15_36_port, S(35) => add_in_15_35_port, S(34)
                           => add_in_15_34_port, S(33) => add_in_15_33_port, 
                           S(32) => add_in_15_32_port, S(31) => 
                           add_in_15_31_port, S(30) => add_in_15_30_port, S(29)
                           => add_in_15_29_port, S(28) => add_in_15_28_port, 
                           S(27) => add_in_15_27_port, S(26) => 
                           add_in_15_26_port, S(25) => add_in_15_25_port, S(24)
                           => add_in_15_24_port, S(23) => add_in_15_23_port, 
                           S(22) => add_in_15_22_port, S(21) => 
                           add_in_15_21_port, S(20) => add_in_15_20_port, S(19)
                           => add_in_15_19_port, S(18) => add_in_15_18_port, 
                           S(17) => add_in_15_17_port, S(16) => 
                           add_in_15_16_port, S(15) => add_in_15_15_port, S(14)
                           => add_in_15_14_port, S(13) => add_in_15_13_port, 
                           S(12) => add_in_15_12_port, S(11) => 
                           add_in_15_11_port, S(10) => add_in_15_10_port, S(9) 
                           => add_in_15_9_port, S(8) => add_in_15_8_port, S(7) 
                           => add_in_15_7_port, S(6) => add_in_15_6_port, S(5) 
                           => add_in_15_5_port, S(4) => add_in_15_4_port, S(3) 
                           => add_in_15_3_port, S(2) => add_in_15_2_port, S(1) 
                           => add_in_15_1_port, S(0) => add_in_15_0_port, Co =>
                           net21306);
   add_128 : BOOTHMUL_N32_DW01_add_0 port map( A(63) => add_in_15_63_port, 
                           A(62) => add_in_15_62_port, A(61) => 
                           add_in_15_61_port, A(60) => add_in_15_60_port, A(59)
                           => add_in_15_59_port, A(58) => add_in_15_58_port, 
                           A(57) => add_in_15_57_port, A(56) => 
                           add_in_15_56_port, A(55) => add_in_15_55_port, A(54)
                           => add_in_15_54_port, A(53) => add_in_15_53_port, 
                           A(52) => add_in_15_52_port, A(51) => 
                           add_in_15_51_port, A(50) => add_in_15_50_port, A(49)
                           => add_in_15_49_port, A(48) => add_in_15_48_port, 
                           A(47) => add_in_15_47_port, A(46) => 
                           add_in_15_46_port, A(45) => add_in_15_45_port, A(44)
                           => add_in_15_44_port, A(43) => add_in_15_43_port, 
                           A(42) => add_in_15_42_port, A(41) => 
                           add_in_15_41_port, A(40) => add_in_15_40_port, A(39)
                           => add_in_15_39_port, A(38) => add_in_15_38_port, 
                           A(37) => add_in_15_37_port, A(36) => 
                           add_in_15_36_port, A(35) => add_in_15_35_port, A(34)
                           => add_in_15_34_port, A(33) => add_in_15_33_port, 
                           A(32) => add_in_15_32_port, A(31) => 
                           add_in_15_31_port, A(30) => add_in_15_30_port, A(29)
                           => add_in_15_29_port, A(28) => add_in_15_28_port, 
                           A(27) => add_in_15_27_port, A(26) => 
                           add_in_15_26_port, A(25) => add_in_15_25_port, A(24)
                           => add_in_15_24_port, A(23) => add_in_15_23_port, 
                           A(22) => add_in_15_22_port, A(21) => 
                           add_in_15_21_port, A(20) => add_in_15_20_port, A(19)
                           => add_in_15_19_port, A(18) => add_in_15_18_port, 
                           A(17) => add_in_15_17_port, A(16) => 
                           add_in_15_16_port, A(15) => add_in_15_15_port, A(14)
                           => add_in_15_14_port, A(13) => add_in_15_13_port, 
                           A(12) => add_in_15_12_port, A(11) => 
                           add_in_15_11_port, A(10) => add_in_15_10_port, A(9) 
                           => add_in_15_9_port, A(8) => add_in_15_8_port, A(7) 
                           => add_in_15_7_port, A(6) => add_in_15_6_port, A(5) 
                           => add_in_15_5_port, A(4) => add_in_15_4_port, A(3) 
                           => add_in_15_3_port, A(2) => add_in_15_2_port, A(1) 
                           => add_in_15_1_port, A(0) => add_in_15_0_port, B(63)
                           => n696, B(62) => n696, B(61) => n696, B(60) => n696
                           , B(59) => n696, B(58) => n696, B(57) => n696, B(56)
                           => n696, B(55) => n696, B(54) => n696, B(53) => n696
                           , B(52) => n696, B(51) => n696, B(50) => n696, B(49)
                           => n696, B(48) => n696, B(47) => n696, B(46) => n696
                           , B(45) => n696, B(44) => n696, B(43) => n696, B(42)
                           => n696, B(41) => n696, B(40) => n696, B(39) => n696
                           , B(38) => n696, B(37) => n696, B(36) => n696, B(35)
                           => n696, B(34) => n696, B(33) => n696, B(32) => n696
                           , B(31) => n696, B(30) => n696, B(29) => n696, B(28)
                           => n696, B(27) => n696, B(26) => n696, B(25) => n696
                           , B(24) => n696, B(23) => n696, B(22) => n696, B(21)
                           => n696, B(20) => n696, B(19) => n696, B(18) => n696
                           , B(17) => n696, B(16) => n696, B(15) => n696, B(14)
                           => n696, B(13) => n696, B(12) => n696, B(11) => n696
                           , B(10) => n696, B(9) => n696, B(8) => n696, B(7) =>
                           n696, B(6) => n696, B(5) => n696, B(4) => n696, B(3)
                           => n696, B(2) => n696, B(1) => n696, B(0) => 
                           mode_15_port, CI => n696, SUM(63) => P(63), SUM(62) 
                           => P(62), SUM(61) => P(61), SUM(60) => P(60), 
                           SUM(59) => P(59), SUM(58) => P(58), SUM(57) => P(57)
                           , SUM(56) => P(56), SUM(55) => P(55), SUM(54) => 
                           P(54), SUM(53) => P(53), SUM(52) => P(52), SUM(51) 
                           => P(51), SUM(50) => P(50), SUM(49) => P(49), 
                           SUM(48) => P(48), SUM(47) => P(47), SUM(46) => P(46)
                           , SUM(45) => P(45), SUM(44) => P(44), SUM(43) => 
                           P(43), SUM(42) => P(42), SUM(41) => P(41), SUM(40) 
                           => P(40), SUM(39) => P(39), SUM(38) => P(38), 
                           SUM(37) => P(37), SUM(36) => P(36), SUM(35) => P(35)
                           , SUM(34) => P(34), SUM(33) => P(33), SUM(32) => 
                           P(32), SUM(31) => P(31), SUM(30) => P(30), SUM(29) 
                           => P(29), SUM(28) => P(28), SUM(27) => P(27), 
                           SUM(26) => P(26), SUM(25) => P(25), SUM(24) => P(24)
                           , SUM(23) => P(23), SUM(22) => P(22), SUM(21) => 
                           P(21), SUM(20) => P(20), SUM(19) => P(19), SUM(18) 
                           => P(18), SUM(17) => P(17), SUM(16) => P(16), 
                           SUM(15) => P(15), SUM(14) => P(14), SUM(13) => P(13)
                           , SUM(12) => P(12), SUM(11) => P(11), SUM(10) => 
                           P(10), SUM(9) => P(9), SUM(8) => P(8), SUM(7) => 
                           P(7), SUM(6) => P(6), SUM(5) => P(5), SUM(4) => P(4)
                           , SUM(3) => P(3), SUM(2) => P(2), SUM(1) => P(1), 
                           SUM(0) => P(0), CO => net165111);
   U130 : BUF_X1 port map( A => n596, Z => n589);
   U131 : CLKBUF_X1 port map( A => n619, Z => n521);
   U132 : CLKBUF_X1 port map( A => n622, Z => n513);
   U133 : CLKBUF_X1 port map( A => n623, Z => n509);
   U134 : CLKBUF_X1 port map( A => n598, Z => n585);
   U135 : BUF_X1 port map( A => n596, Z => n591);
   U136 : BUF_X1 port map( A => n596, Z => n590);
   U137 : CLKBUF_X1 port map( A => n595, Z => n594);
   U138 : CLKBUF_X1 port map( A => n610, Z => n549);
   U139 : CLKBUF_X1 port map( A => n613, Z => n540);
   U140 : CLKBUF_X1 port map( A => n612, Z => n543);
   U141 : CLKBUF_X1 port map( A => n615, Z => n533);
   U142 : CLKBUF_X1 port map( A => n614, Z => n537);
   U143 : CLKBUF_X1 port map( A => n616, Z => n530);
   U144 : CLKBUF_X1 port map( A => n609, Z => n552);
   U145 : CLKBUF_X1 port map( A => n605, Z => n564);
   U146 : CLKBUF_X1 port map( A => n624, Z => n623);
   U147 : CLKBUF_X1 port map( A => n632, Z => n597);
   U148 : CLKBUF_X1 port map( A => n625, Z => n620);
   U149 : CLKBUF_X1 port map( A => n627, Z => n612);
   U150 : CLKBUF_X1 port map( A => n629, Z => n606);
   U151 : BUF_X1 port map( A => n403, Z => n402);
   U152 : CLKBUF_X1 port map( A => n635, Z => n625);
   U153 : CLKBUF_X1 port map( A => n634, Z => n632);
   U154 : CLKBUF_X1 port map( A => n635, Z => n626);
   U155 : INV_X1 port map( A => n592, ZN => n654);
   U156 : INV_X1 port map( A => n594, ZN => n637);
   U157 : INV_X1 port map( A => n591, ZN => n661);
   U158 : INV_X1 port map( A => n589, ZN => n674);
   U159 : INV_X1 port map( A => n594, ZN => n640);
   U160 : INV_X1 port map( A => n594, ZN => n639);
   U161 : INV_X1 port map( A => n594, ZN => n638);
   U162 : INV_X1 port map( A => n588, ZN => n680);
   U163 : INV_X1 port map( A => n593, ZN => n647);
   U164 : INV_X1 port map( A => n590, ZN => n668);
   U165 : BUF_X2 port map( A => n595, Z => n592);
   U166 : BUF_X1 port map( A => n597, Z => n588);
   U167 : BUF_X1 port map( A => n600, Z => n578);
   U168 : BUF_X1 port map( A => n618, Z => n525);
   U169 : BUF_X1 port map( A => n599, Z => n580);
   U170 : BUF_X1 port map( A => n620, Z => n517);
   U171 : BUF_X1 port map( A => n598, Z => n583);
   U172 : BUF_X1 port map( A => n622, Z => n512);
   U173 : CLKBUF_X1 port map( A => n600, Z => n579);
   U174 : BUF_X1 port map( A => n623, Z => n508);
   U175 : CLKBUF_X1 port map( A => n598, Z => n584);
   U176 : BUF_X1 port map( A => n619, Z => n520);
   U177 : BUF_X1 port map( A => n621, Z => n516);
   U178 : BUF_X1 port map( A => n617, Z => n528);
   U179 : BUF_X1 port map( A => n618, Z => n524);
   U180 : CLKBUF_X1 port map( A => n595, Z => n593);
   U181 : BUF_X1 port map( A => n611, Z => n546);
   U182 : CLKBUF_X1 port map( A => n617, Z => n526);
   U183 : BUF_X1 port map( A => n614, Z => n536);
   U184 : CLKBUF_X1 port map( A => n615, Z => n534);
   U185 : BUF_X1 port map( A => n613, Z => n539);
   U186 : BUF_X1 port map( A => n616, Z => n529);
   U187 : CLKBUF_X1 port map( A => n619, Z => n522);
   U188 : CLKBUF_X1 port map( A => n620, Z => n518);
   U189 : BUF_X1 port map( A => n610, Z => n548);
   U190 : CLKBUF_X1 port map( A => n621, Z => n514);
   U191 : BUF_X1 port map( A => n611, Z => n545);
   U192 : CLKBUF_X1 port map( A => n599, Z => n581);
   U193 : CLKBUF_X1 port map( A => n623, Z => n510);
   U194 : BUF_X1 port map( A => n612, Z => n542);
   U195 : BUF_X1 port map( A => n615, Z => n532);
   U196 : CLKBUF_X1 port map( A => n617, Z => n527);
   U197 : CLKBUF_X1 port map( A => n618, Z => n523);
   U198 : CLKBUF_X1 port map( A => n597, Z => n586);
   U199 : CLKBUF_X1 port map( A => n616, Z => n531);
   U200 : CLKBUF_X1 port map( A => n620, Z => n519);
   U201 : BUF_X1 port map( A => n614, Z => n535);
   U202 : CLKBUF_X1 port map( A => n621, Z => n515);
   U203 : CLKBUF_X1 port map( A => n599, Z => n582);
   U204 : CLKBUF_X1 port map( A => n622, Z => n511);
   U205 : CLKBUF_X1 port map( A => n597, Z => n587);
   U206 : BUF_X1 port map( A => n607, Z => n557);
   U207 : BUF_X1 port map( A => n606, Z => n559);
   U208 : BUF_X1 port map( A => n604, Z => n567);
   U209 : BUF_X1 port map( A => n605, Z => n563);
   U210 : CLKBUF_X1 port map( A => n605, Z => n562);
   U211 : BUF_X1 port map( A => n608, Z => n554);
   U212 : CLKBUF_X1 port map( A => n608, Z => n555);
   U213 : CLKBUF_X1 port map( A => n606, Z => n561);
   U214 : CLKBUF_X1 port map( A => n606, Z => n560);
   U215 : BUF_X1 port map( A => n604, Z => n565);
   U216 : CLKBUF_X1 port map( A => n610, Z => n547);
   U217 : CLKBUF_X1 port map( A => n609, Z => n550);
   U218 : CLKBUF_X1 port map( A => n611, Z => n544);
   U219 : CLKBUF_X1 port map( A => n607, Z => n558);
   U220 : CLKBUF_X1 port map( A => n608, Z => n553);
   U221 : BUF_X1 port map( A => n609, Z => n551);
   U222 : CLKBUF_X1 port map( A => n612, Z => n541);
   U223 : CLKBUF_X1 port map( A => n607, Z => n556);
   U224 : CLKBUF_X1 port map( A => n613, Z => n538);
   U225 : CLKBUF_X1 port map( A => n604, Z => n566);
   U226 : BUF_X1 port map( A => n603, Z => n570);
   U227 : BUF_X1 port map( A => n602, Z => n571);
   U228 : BUF_X1 port map( A => n603, Z => n568);
   U229 : CLKBUF_X1 port map( A => n602, Z => n573);
   U230 : CLKBUF_X1 port map( A => n603, Z => n569);
   U231 : BUF_X1 port map( A => n601, Z => n574);
   U232 : CLKBUF_X1 port map( A => n602, Z => n572);
   U233 : BUF_X1 port map( A => n601, Z => n575);
   U234 : CLKBUF_X1 port map( A => n601, Z => n576);
   U235 : CLKBUF_X1 port map( A => n600, Z => n577);
   U236 : INV_X1 port map( A => n202, ZN => n205);
   U237 : INV_X1 port map( A => n212, ZN => n215);
   U238 : INV_X1 port map( A => n222, ZN => n225);
   U239 : INV_X1 port map( A => n232, ZN => n235);
   U240 : INV_X1 port map( A => n242, ZN => n245);
   U241 : INV_X1 port map( A => n252, ZN => n255);
   U242 : INV_X1 port map( A => n262, ZN => n265);
   U243 : INV_X1 port map( A => n272, ZN => n275);
   U244 : INV_X1 port map( A => n282, ZN => n285);
   U245 : INV_X1 port map( A => n292, ZN => n295);
   U246 : INV_X1 port map( A => n302, ZN => n305);
   U247 : INV_X1 port map( A => n312, ZN => n315);
   U248 : INV_X1 port map( A => n322, ZN => n325);
   U249 : INV_X1 port map( A => n332, ZN => n335);
   U250 : INV_X1 port map( A => n202, ZN => n206);
   U251 : INV_X1 port map( A => n212, ZN => n216);
   U252 : INV_X1 port map( A => n222, ZN => n226);
   U253 : INV_X1 port map( A => n232, ZN => n236);
   U254 : INV_X1 port map( A => n242, ZN => n246);
   U255 : INV_X1 port map( A => n252, ZN => n256);
   U256 : INV_X1 port map( A => n262, ZN => n266);
   U257 : INV_X1 port map( A => n272, ZN => n276);
   U258 : INV_X1 port map( A => n282, ZN => n286);
   U259 : INV_X1 port map( A => n292, ZN => n296);
   U260 : INV_X1 port map( A => n302, ZN => n306);
   U261 : INV_X1 port map( A => n312, ZN => n316);
   U262 : INV_X1 port map( A => n322, ZN => n326);
   U263 : INV_X1 port map( A => n452, ZN => n455);
   U264 : INV_X1 port map( A => n472, ZN => n475);
   U265 : INV_X1 port map( A => n462, ZN => n465);
   U266 : INV_X1 port map( A => n432, ZN => n435);
   U267 : INV_X1 port map( A => n492, ZN => n495);
   U268 : INV_X1 port map( A => n482, ZN => n485);
   U269 : INV_X1 port map( A => n442, ZN => n445);
   U270 : INV_X1 port map( A => n412, ZN => n415);
   U271 : INV_X1 port map( A => n422, ZN => n425);
   U272 : INV_X1 port map( A => n402, ZN => n405);
   U273 : INV_X1 port map( A => n342, ZN => n345);
   U274 : INV_X1 port map( A => n352, ZN => n355);
   U275 : INV_X1 port map( A => n362, ZN => n365);
   U276 : INV_X1 port map( A => n372, ZN => n375);
   U277 : INV_X1 port map( A => n382, ZN => n385);
   U278 : INV_X1 port map( A => n392, ZN => n395);
   U279 : INV_X1 port map( A => n472, ZN => n476);
   U280 : INV_X1 port map( A => n462, ZN => n466);
   U281 : INV_X1 port map( A => n452, ZN => n456);
   U282 : INV_X1 port map( A => n442, ZN => n446);
   U283 : INV_X1 port map( A => n432, ZN => n436);
   U284 : INV_X1 port map( A => n422, ZN => n426);
   U285 : INV_X1 port map( A => n412, ZN => n416);
   U286 : INV_X1 port map( A => n402, ZN => n406);
   U287 : INV_X1 port map( A => n332, ZN => n336);
   U288 : INV_X1 port map( A => n342, ZN => n346);
   U289 : INV_X1 port map( A => n352, ZN => n356);
   U290 : INV_X1 port map( A => n362, ZN => n366);
   U291 : INV_X1 port map( A => n372, ZN => n376);
   U292 : INV_X1 port map( A => n382, ZN => n386);
   U293 : INV_X1 port map( A => n392, ZN => n396);
   U294 : INV_X1 port map( A => n502, ZN => n505);
   U295 : INV_X1 port map( A => n502, ZN => n506);
   U296 : INV_X1 port map( A => n482, ZN => n486);
   U297 : INV_X1 port map( A => n492, ZN => n496);
   U298 : BUF_X1 port map( A => n631, Z => n600);
   U299 : BUF_X1 port map( A => n626, Z => n617);
   U300 : BUF_X1 port map( A => n625, Z => n619);
   U301 : BUF_X1 port map( A => n632, Z => n598);
   U302 : CLKBUF_X1 port map( A => n625, Z => n618);
   U303 : CLKBUF_X1 port map( A => n632, Z => n599);
   U304 : CLKBUF_X1 port map( A => n624, Z => n621);
   U305 : BUF_X1 port map( A => n624, Z => n622);
   U306 : BUF_X1 port map( A => n633, Z => n595);
   U307 : CLKBUF_X1 port map( A => n633, Z => n596);
   U308 : BUF_X1 port map( A => n628, Z => n610);
   U309 : CLKBUF_X1 port map( A => n628, Z => n611);
   U310 : CLKBUF_X1 port map( A => n627, Z => n613);
   U311 : CLKBUF_X1 port map( A => n626, Z => n615);
   U312 : BUF_X1 port map( A => n627, Z => n614);
   U313 : CLKBUF_X1 port map( A => n626, Z => n616);
   U314 : BUF_X1 port map( A => n630, Z => n605);
   U315 : CLKBUF_X1 port map( A => n630, Z => n604);
   U316 : CLKBUF_X1 port map( A => n629, Z => n607);
   U317 : BUF_X1 port map( A => n629, Z => n608);
   U318 : CLKBUF_X1 port map( A => n628, Z => n609);
   U319 : CLKBUF_X1 port map( A => n630, Z => n603);
   U320 : CLKBUF_X1 port map( A => n631, Z => n602);
   U321 : CLKBUF_X1 port map( A => n631, Z => n601);
   U322 : BUF_X2 port map( A => n203, Z => n202);
   U323 : BUF_X2 port map( A => n213, Z => n212);
   U324 : BUF_X1 port map( A => n223, Z => n222);
   U325 : BUF_X1 port map( A => n233, Z => n232);
   U326 : BUF_X1 port map( A => n243, Z => n242);
   U327 : BUF_X1 port map( A => n253, Z => n252);
   U328 : BUF_X1 port map( A => n263, Z => n262);
   U329 : BUF_X1 port map( A => n273, Z => n272);
   U330 : BUF_X1 port map( A => n283, Z => n282);
   U331 : BUF_X1 port map( A => n293, Z => n292);
   U332 : BUF_X1 port map( A => n303, Z => n302);
   U333 : BUF_X1 port map( A => n313, Z => n312);
   U334 : BUF_X1 port map( A => n323, Z => n322);
   U335 : BUF_X1 port map( A => n333, Z => n332);
   U336 : BUF_X1 port map( A => n204, Z => n198);
   U337 : BUF_X1 port map( A => n214, Z => n208);
   U338 : BUF_X1 port map( A => n224, Z => n218);
   U339 : BUF_X1 port map( A => n234, Z => n228);
   U340 : BUF_X1 port map( A => n244, Z => n238);
   U341 : BUF_X1 port map( A => n254, Z => n248);
   U342 : BUF_X1 port map( A => n264, Z => n258);
   U343 : BUF_X1 port map( A => n274, Z => n268);
   U344 : BUF_X1 port map( A => n284, Z => n278);
   U345 : BUF_X1 port map( A => n294, Z => n288);
   U346 : BUF_X2 port map( A => n453, Z => n452);
   U347 : BUF_X2 port map( A => n493, Z => n492);
   U348 : BUF_X2 port map( A => n473, Z => n472);
   U349 : BUF_X2 port map( A => n463, Z => n462);
   U350 : BUF_X2 port map( A => n483, Z => n482);
   U351 : BUF_X2 port map( A => n433, Z => n432);
   U352 : BUF_X2 port map( A => n443, Z => n442);
   U353 : BUF_X2 port map( A => n413, Z => n412);
   U354 : BUF_X2 port map( A => n423, Z => n422);
   U355 : BUF_X1 port map( A => n343, Z => n342);
   U356 : BUF_X1 port map( A => n353, Z => n352);
   U357 : BUF_X1 port map( A => n363, Z => n362);
   U358 : BUF_X1 port map( A => n373, Z => n372);
   U359 : BUF_X1 port map( A => n383, Z => n382);
   U360 : BUF_X1 port map( A => n393, Z => n392);
   U361 : BUF_X1 port map( A => n304, Z => n298);
   U362 : BUF_X1 port map( A => n314, Z => n308);
   U363 : BUF_X1 port map( A => n324, Z => n318);
   U364 : CLKBUF_X1 port map( A => n204, Z => n199);
   U365 : BUF_X1 port map( A => n334, Z => n328);
   U366 : BUF_X1 port map( A => n344, Z => n338);
   U367 : CLKBUF_X1 port map( A => n214, Z => n209);
   U368 : BUF_X1 port map( A => n354, Z => n348);
   U369 : CLKBUF_X1 port map( A => n224, Z => n219);
   U370 : BUF_X1 port map( A => n364, Z => n358);
   U371 : CLKBUF_X1 port map( A => n234, Z => n229);
   U372 : BUF_X1 port map( A => n374, Z => n368);
   U373 : CLKBUF_X1 port map( A => n244, Z => n239);
   U374 : BUF_X1 port map( A => n384, Z => n378);
   U375 : CLKBUF_X1 port map( A => n254, Z => n249);
   U376 : BUF_X1 port map( A => n394, Z => n388);
   U377 : CLKBUF_X1 port map( A => n264, Z => n259);
   U378 : BUF_X1 port map( A => n404, Z => n398);
   U379 : CLKBUF_X1 port map( A => n274, Z => n269);
   U380 : BUF_X1 port map( A => n414, Z => n408);
   U381 : CLKBUF_X1 port map( A => n284, Z => n279);
   U382 : BUF_X1 port map( A => n424, Z => n418);
   U383 : CLKBUF_X1 port map( A => n294, Z => n289);
   U384 : BUF_X1 port map( A => n434, Z => n428);
   U385 : CLKBUF_X1 port map( A => n304, Z => n299);
   U386 : BUF_X1 port map( A => n444, Z => n438);
   U387 : CLKBUF_X1 port map( A => n314, Z => n309);
   U388 : BUF_X1 port map( A => n454, Z => n448);
   U389 : BUF_X2 port map( A => n503, Z => n502);
   U390 : CLKBUF_X1 port map( A => n203, Z => n200);
   U391 : CLKBUF_X1 port map( A => n213, Z => n210);
   U392 : CLKBUF_X1 port map( A => n223, Z => n220);
   U393 : CLKBUF_X1 port map( A => n233, Z => n230);
   U394 : CLKBUF_X1 port map( A => n243, Z => n240);
   U395 : CLKBUF_X1 port map( A => n253, Z => n250);
   U396 : CLKBUF_X1 port map( A => n263, Z => n260);
   U397 : CLKBUF_X1 port map( A => n273, Z => n270);
   U398 : CLKBUF_X1 port map( A => n283, Z => n280);
   U399 : CLKBUF_X1 port map( A => n293, Z => n290);
   U400 : CLKBUF_X1 port map( A => n324, Z => n319);
   U401 : BUF_X1 port map( A => n464, Z => n458);
   U402 : CLKBUF_X1 port map( A => n334, Z => n329);
   U403 : BUF_X1 port map( A => n474, Z => n468);
   U404 : BUF_X1 port map( A => n484, Z => n478);
   U405 : CLKBUF_X1 port map( A => n344, Z => n339);
   U406 : BUF_X1 port map( A => n494, Z => n488);
   U407 : CLKBUF_X1 port map( A => n354, Z => n349);
   U408 : CLKBUF_X1 port map( A => n364, Z => n359);
   U409 : BUF_X1 port map( A => n504, Z => n498);
   U410 : CLKBUF_X1 port map( A => n374, Z => n369);
   U411 : CLKBUF_X1 port map( A => n384, Z => n379);
   U412 : CLKBUF_X1 port map( A => n474, Z => n469);
   U413 : CLKBUF_X1 port map( A => n394, Z => n389);
   U414 : CLKBUF_X1 port map( A => n404, Z => n399);
   U415 : CLKBUF_X1 port map( A => n414, Z => n409);
   U416 : CLKBUF_X1 port map( A => n424, Z => n419);
   U417 : CLKBUF_X1 port map( A => n434, Z => n429);
   U418 : CLKBUF_X1 port map( A => n464, Z => n459);
   U419 : CLKBUF_X1 port map( A => n444, Z => n439);
   U420 : CLKBUF_X1 port map( A => n454, Z => n449);
   U421 : CLKBUF_X1 port map( A => n634, Z => n631);
   U422 : BUF_X1 port map( A => n635, Z => n624);
   U423 : BUF_X1 port map( A => n634, Z => n633);
   U424 : CLKBUF_X1 port map( A => n443, Z => n440);
   U425 : CLKBUF_X1 port map( A => n433, Z => n430);
   U426 : CLKBUF_X1 port map( A => n423, Z => n420);
   U427 : CLKBUF_X1 port map( A => n303, Z => n300);
   U428 : CLKBUF_X1 port map( A => n313, Z => n310);
   U429 : CLKBUF_X1 port map( A => n323, Z => n320);
   U430 : CLKBUF_X1 port map( A => n333, Z => n330);
   U431 : CLKBUF_X1 port map( A => n203, Z => n201);
   U432 : CLKBUF_X1 port map( A => n343, Z => n340);
   U433 : CLKBUF_X1 port map( A => n213, Z => n211);
   U434 : CLKBUF_X1 port map( A => n353, Z => n350);
   U435 : CLKBUF_X1 port map( A => n223, Z => n221);
   U436 : CLKBUF_X1 port map( A => n363, Z => n360);
   U437 : CLKBUF_X1 port map( A => n233, Z => n231);
   U438 : CLKBUF_X1 port map( A => n373, Z => n370);
   U439 : CLKBUF_X1 port map( A => n413, Z => n410);
   U440 : CLKBUF_X1 port map( A => n243, Z => n241);
   U441 : CLKBUF_X1 port map( A => n383, Z => n380);
   U442 : CLKBUF_X1 port map( A => n253, Z => n251);
   U443 : CLKBUF_X1 port map( A => n393, Z => n390);
   U444 : CLKBUF_X1 port map( A => n263, Z => n261);
   U445 : CLKBUF_X1 port map( A => n403, Z => n400);
   U446 : CLKBUF_X1 port map( A => n273, Z => n271);
   U447 : CLKBUF_X1 port map( A => n283, Z => n281);
   U448 : CLKBUF_X1 port map( A => n293, Z => n291);
   U449 : CLKBUF_X1 port map( A => n303, Z => n301);
   U450 : CLKBUF_X1 port map( A => n504, Z => n499);
   U451 : CLKBUF_X1 port map( A => n494, Z => n489);
   U452 : CLKBUF_X1 port map( A => n484, Z => n479);
   U453 : CLKBUF_X1 port map( A => n635, Z => n628);
   U454 : CLKBUF_X1 port map( A => n635, Z => n627);
   U455 : CLKBUF_X1 port map( A => n503, Z => n500);
   U456 : CLKBUF_X1 port map( A => n463, Z => n461);
   U457 : CLKBUF_X1 port map( A => n453, Z => n451);
   U458 : CLKBUF_X1 port map( A => n493, Z => n490);
   U459 : CLKBUF_X1 port map( A => n443, Z => n441);
   U460 : CLKBUF_X1 port map( A => n483, Z => n480);
   U461 : CLKBUF_X1 port map( A => n433, Z => n431);
   U462 : CLKBUF_X1 port map( A => n473, Z => n470);
   U463 : CLKBUF_X1 port map( A => n423, Z => n421);
   U464 : CLKBUF_X1 port map( A => n463, Z => n460);
   U465 : CLKBUF_X1 port map( A => n453, Z => n450);
   U466 : CLKBUF_X1 port map( A => n413, Z => n411);
   U467 : CLKBUF_X1 port map( A => n403, Z => n401);
   U468 : CLKBUF_X1 port map( A => n393, Z => n391);
   U469 : CLKBUF_X1 port map( A => n313, Z => n311);
   U470 : CLKBUF_X1 port map( A => n323, Z => n321);
   U471 : CLKBUF_X1 port map( A => n333, Z => n331);
   U472 : CLKBUF_X1 port map( A => n343, Z => n341);
   U473 : CLKBUF_X1 port map( A => n353, Z => n351);
   U474 : CLKBUF_X1 port map( A => n363, Z => n361);
   U475 : CLKBUF_X1 port map( A => n373, Z => n371);
   U476 : CLKBUF_X1 port map( A => n383, Z => n381);
   U477 : CLKBUF_X1 port map( A => n634, Z => n630);
   U478 : CLKBUF_X1 port map( A => n634, Z => n629);
   U479 : CLKBUF_X1 port map( A => n473, Z => n471);
   U480 : CLKBUF_X1 port map( A => n483, Z => n481);
   U481 : CLKBUF_X1 port map( A => n493, Z => n491);
   U482 : CLKBUF_X1 port map( A => n503, Z => n501);
   U483 : BUF_X1 port map( A => A(0), Z => n203);
   U484 : BUF_X1 port map( A => A(1), Z => n213);
   U485 : BUF_X1 port map( A => A(2), Z => n223);
   U486 : BUF_X1 port map( A => A(3), Z => n233);
   U487 : BUF_X1 port map( A => A(4), Z => n243);
   U488 : BUF_X1 port map( A => A(5), Z => n253);
   U489 : BUF_X1 port map( A => A(6), Z => n263);
   U490 : BUF_X1 port map( A => A(7), Z => n273);
   U491 : BUF_X1 port map( A => A(8), Z => n283);
   U492 : BUF_X1 port map( A => A(9), Z => n293);
   U493 : BUF_X1 port map( A => A(10), Z => n303);
   U494 : BUF_X1 port map( A => A(11), Z => n313);
   U495 : BUF_X1 port map( A => A(12), Z => n323);
   U496 : BUF_X1 port map( A => A(13), Z => n333);
   U497 : BUF_X1 port map( A => A(0), Z => n204);
   U498 : BUF_X1 port map( A => A(1), Z => n214);
   U499 : BUF_X1 port map( A => A(2), Z => n224);
   U500 : BUF_X1 port map( A => A(3), Z => n234);
   U501 : BUF_X1 port map( A => A(4), Z => n244);
   U502 : BUF_X1 port map( A => A(5), Z => n254);
   U503 : BUF_X1 port map( A => A(6), Z => n264);
   U504 : BUF_X1 port map( A => A(7), Z => n274);
   U505 : BUF_X1 port map( A => A(8), Z => n284);
   U506 : BUF_X1 port map( A => A(9), Z => n294);
   U507 : BUF_X1 port map( A => A(29), Z => n493);
   U508 : BUF_X1 port map( A => A(27), Z => n473);
   U509 : BUF_X1 port map( A => A(28), Z => n483);
   U510 : BUF_X1 port map( A => A(25), Z => n453);
   U511 : BUF_X1 port map( A => A(26), Z => n463);
   U512 : BUF_X1 port map( A => A(23), Z => n433);
   U513 : BUF_X1 port map( A => A(24), Z => n443);
   U514 : BUF_X1 port map( A => A(22), Z => n423);
   U515 : BUF_X1 port map( A => A(21), Z => n413);
   U516 : BUF_X1 port map( A => A(20), Z => n403);
   U517 : BUF_X1 port map( A => A(14), Z => n343);
   U518 : BUF_X1 port map( A => A(15), Z => n353);
   U519 : BUF_X1 port map( A => A(16), Z => n363);
   U520 : BUF_X1 port map( A => A(17), Z => n373);
   U521 : BUF_X1 port map( A => A(19), Z => n393);
   U522 : BUF_X1 port map( A => A(18), Z => n383);
   U523 : BUF_X1 port map( A => A(10), Z => n304);
   U524 : BUF_X1 port map( A => A(11), Z => n314);
   U525 : BUF_X1 port map( A => A(12), Z => n324);
   U526 : BUF_X1 port map( A => A(13), Z => n334);
   U527 : BUF_X1 port map( A => A(14), Z => n344);
   U528 : BUF_X1 port map( A => A(15), Z => n354);
   U529 : BUF_X1 port map( A => A(16), Z => n364);
   U530 : BUF_X1 port map( A => A(17), Z => n374);
   U531 : BUF_X1 port map( A => A(18), Z => n384);
   U532 : BUF_X1 port map( A => A(19), Z => n394);
   U533 : BUF_X1 port map( A => A(20), Z => n404);
   U534 : BUF_X1 port map( A => A(21), Z => n414);
   U535 : BUF_X1 port map( A => A(22), Z => n424);
   U536 : BUF_X1 port map( A => A(23), Z => n434);
   U537 : BUF_X1 port map( A => A(24), Z => n444);
   U538 : BUF_X1 port map( A => A(25), Z => n454);
   U539 : BUF_X1 port map( A => A(30), Z => n503);
   U540 : BUF_X2 port map( A => A(31), Z => n634);
   U541 : BUF_X1 port map( A => A(31), Z => n635);
   U542 : BUF_X1 port map( A => A(30), Z => n504);
   U543 : BUF_X1 port map( A => A(29), Z => n494);
   U544 : BUF_X1 port map( A => A(28), Z => n484);
   U545 : BUF_X1 port map( A => A(27), Z => n474);
   U546 : BUF_X1 port map( A => A(26), Z => n464);
   U547 : INV_X1 port map( A => n202, ZN => n207);
   U548 : INV_X1 port map( A => n212, ZN => n217);
   U549 : INV_X1 port map( A => n222, ZN => n227);
   U550 : INV_X1 port map( A => n232, ZN => n237);
   U551 : INV_X1 port map( A => n242, ZN => n247);
   U552 : INV_X1 port map( A => n252, ZN => n257);
   U553 : INV_X1 port map( A => n262, ZN => n267);
   U554 : INV_X1 port map( A => n272, ZN => n277);
   U555 : INV_X1 port map( A => n282, ZN => n287);
   U556 : INV_X1 port map( A => n292, ZN => n297);
   U557 : INV_X1 port map( A => n302, ZN => n307);
   U558 : INV_X1 port map( A => n312, ZN => n317);
   U559 : INV_X1 port map( A => n322, ZN => n327);
   U560 : INV_X1 port map( A => n332, ZN => n337);
   U561 : INV_X1 port map( A => n342, ZN => n347);
   U562 : INV_X1 port map( A => n352, ZN => n357);
   U563 : INV_X1 port map( A => n362, ZN => n367);
   U564 : INV_X1 port map( A => n372, ZN => n377);
   U565 : INV_X1 port map( A => n382, ZN => n387);
   U566 : INV_X1 port map( A => n392, ZN => n397);
   U567 : INV_X1 port map( A => n402, ZN => n407);
   U568 : INV_X1 port map( A => n412, ZN => n417);
   U569 : INV_X1 port map( A => n422, ZN => n427);
   U570 : INV_X1 port map( A => n432, ZN => n437);
   U571 : INV_X1 port map( A => n442, ZN => n447);
   U572 : INV_X1 port map( A => n452, ZN => n457);
   U573 : INV_X1 port map( A => n462, ZN => n467);
   U574 : INV_X1 port map( A => n472, ZN => n477);
   U575 : INV_X1 port map( A => n482, ZN => n487);
   U576 : INV_X1 port map( A => n492, ZN => n497);
   U577 : INV_X1 port map( A => n502, ZN => n507);
   U578 : INV_X1 port map( A => n594, ZN => n636);
   U579 : INV_X1 port map( A => n593, ZN => n641);
   U580 : INV_X1 port map( A => n593, ZN => n642);
   U581 : INV_X1 port map( A => n593, ZN => n643);
   U582 : INV_X1 port map( A => n593, ZN => n644);
   U583 : INV_X1 port map( A => n593, ZN => n645);
   U584 : INV_X1 port map( A => n593, ZN => n646);
   U585 : INV_X1 port map( A => n592, ZN => n648);
   U586 : INV_X1 port map( A => n592, ZN => n649);
   U587 : INV_X1 port map( A => n592, ZN => n650);
   U588 : INV_X1 port map( A => n592, ZN => n651);
   U589 : INV_X1 port map( A => n592, ZN => n652);
   U590 : INV_X1 port map( A => n592, ZN => n653);
   U591 : INV_X1 port map( A => n591, ZN => n655);
   U592 : INV_X1 port map( A => n591, ZN => n656);
   U593 : INV_X1 port map( A => n591, ZN => n657);
   U594 : INV_X1 port map( A => n591, ZN => n658);
   U595 : INV_X1 port map( A => n591, ZN => n659);
   U596 : INV_X1 port map( A => n591, ZN => n660);
   U597 : INV_X1 port map( A => n590, ZN => n662);
   U598 : INV_X1 port map( A => n590, ZN => n663);
   U599 : INV_X1 port map( A => n590, ZN => n664);
   U600 : INV_X1 port map( A => n590, ZN => n665);
   U601 : INV_X1 port map( A => n590, ZN => n666);
   U602 : INV_X1 port map( A => n590, ZN => n667);
   U603 : INV_X1 port map( A => n589, ZN => n669);
   U604 : INV_X1 port map( A => n589, ZN => n670);
   U605 : INV_X1 port map( A => n589, ZN => n671);
   U606 : INV_X1 port map( A => n589, ZN => n672);
   U607 : INV_X1 port map( A => n589, ZN => n673);
   U608 : INV_X1 port map( A => n588, ZN => n675);
   U609 : INV_X1 port map( A => n588, ZN => n676);
   U610 : INV_X1 port map( A => n588, ZN => n677);
   U611 : INV_X1 port map( A => n588, ZN => n678);
   U612 : INV_X1 port map( A => n588, ZN => n679);
   U613 : INV_X1 port map( A => B(29), ZN => n681);
   U614 : AOI21_X1 port map( B1 => B(28), B2 => B(27), A => n681, ZN => 
                           mode_14_port);
   U615 : INV_X1 port map( A => B(27), ZN => n682);
   U616 : AOI21_X1 port map( B1 => B(26), B2 => B(25), A => n682, ZN => 
                           mode_13_port);
   U617 : INV_X1 port map( A => B(25), ZN => n683);
   U618 : AOI21_X1 port map( B1 => B(24), B2 => B(23), A => n683, ZN => 
                           mode_12_port);
   U619 : INV_X1 port map( A => B(23), ZN => n684);
   U620 : AOI21_X1 port map( B1 => B(22), B2 => B(21), A => n684, ZN => 
                           mode_11_port);
   U621 : INV_X1 port map( A => B(21), ZN => n685);
   U622 : AOI21_X1 port map( B1 => B(20), B2 => B(19), A => n685, ZN => 
                           mode_10_port);
   U623 : INV_X1 port map( A => B(19), ZN => n686);
   U624 : AOI21_X1 port map( B1 => B(18), B2 => B(17), A => n686, ZN => 
                           mode_9_port);
   U625 : INV_X1 port map( A => B(17), ZN => n687);
   U626 : AOI21_X1 port map( B1 => B(16), B2 => B(15), A => n687, ZN => 
                           mode_8_port);
   U627 : INV_X1 port map( A => B(15), ZN => n688);
   U628 : AOI21_X1 port map( B1 => B(14), B2 => B(13), A => n688, ZN => 
                           mode_7_port);
   U629 : INV_X1 port map( A => B(13), ZN => n689);
   U630 : AOI21_X1 port map( B1 => B(12), B2 => B(11), A => n689, ZN => 
                           mode_6_port);
   U631 : INV_X1 port map( A => B(11), ZN => n690);
   U632 : AOI21_X1 port map( B1 => B(10), B2 => B(9), A => n690, ZN => 
                           mode_5_port);
   U633 : INV_X1 port map( A => B(9), ZN => n691);
   U634 : AOI21_X1 port map( B1 => B(8), B2 => B(7), A => n691, ZN => 
                           mode_4_port);
   U635 : INV_X1 port map( A => B(7), ZN => n692);
   U636 : AOI21_X1 port map( B1 => B(6), B2 => B(5), A => n692, ZN => 
                           mode_3_port);
   U637 : INV_X1 port map( A => B(5), ZN => n693);
   U638 : AOI21_X1 port map( B1 => B(4), B2 => B(3), A => n693, ZN => 
                           mode_2_port);
   U639 : INV_X1 port map( A => B(3), ZN => n694);
   U640 : AOI21_X1 port map( B1 => B(2), B2 => B(1), A => n694, ZN => 
                           mode_1_port);
   U641 : INV_X1 port map( A => B(31), ZN => n695);
   U642 : AOI21_X1 port map( B1 => B(30), B2 => B(29), A => n695, ZN => 
                           mode_15_port);
   n696 <= '0';

end SYN_STRUCTURAL;
