
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4.all;

entity register_file_reg_size64_file_size4_1 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_reg_size64_file_size4_1;

architecture SYN_BEHAVIORAL of register_file_reg_size64_file_size4_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n415, n1200, n1202, n1204, n1310, n1311, n1312, n1313, n1314, n1315
      , n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n871, n872, 
      n873, n875, n876, n936, n938, n939, n975, n978, n979, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176 : std_logic
      ;

begin
   
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => n174,
                           QN => n2028);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => n175,
                           QN => n2027);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => n176,
                           QN => n2026);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => n177,
                           QN => n2025);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => n178,
                           QN => n2024);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => n179,
                           QN => n2023);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => n180,
                           QN => n2022);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => n181,
                           QN => n2021);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => n182,
                           QN => n2020);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => n183, 
                           QN => n2019);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => n184, 
                           QN => n2018);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => n185, 
                           QN => n2017);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => n186, 
                           QN => n2016);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => n187, 
                           QN => n2015);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => n188, 
                           QN => n2014);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => n189, 
                           QN => n2013);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => n190, 
                           QN => n2012);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => n191, 
                           QN => n2011);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => n192, 
                           QN => n2010);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => n65, 
                           QN => n2063);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => n66, 
                           QN => n2062);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n67, 
                           QN => n2061);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => n68, 
                           QN => n2060);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => n69, 
                           QN => n2059);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => n70, 
                           QN => n2058);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => n71, 
                           QN => n2057);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => n72, 
                           QN => n2056);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => n73, 
                           QN => n2055);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => n74, 
                           QN => n2054);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => n75, 
                           QN => n2053);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => n76, 
                           QN => n2052);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => n77, 
                           QN => n2051);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => n78, 
                           QN => n2050);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => n79, 
                           QN => n2049);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => n80, 
                           QN => n2048);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => n81, 
                           QN => n2047);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => n82, 
                           QN => n2046);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => n83, 
                           QN => n2045);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => n84, 
                           QN => n2044);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => n85, 
                           QN => n2043);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => n86, 
                           QN => n2042);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => n87, 
                           QN => n2041);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => n88, 
                           QN => n2040);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => n89, 
                           QN => n2039);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => n90, 
                           QN => n2038);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => n91, 
                           QN => n2037);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => n92, 
                           QN => n2036);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => n93, 
                           QN => n2035);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => n94, 
                           QN => n2034);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => n95, 
                           QN => n2033);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => n96, 
                           QN => n2032);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => n97, 
                           QN => n2031);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => n98, 
                           QN => n2030);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => n99, 
                           QN => n2029);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => n2, 
                           QN => n2009);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => n3, 
                           QN => n2008);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => n4, 
                           QN => n2007);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => n5, 
                           QN => n2006);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => n6, 
                           QN => n2005);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => n7, 
                           QN => n2004);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => n8, 
                           QN => n2003);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => n9, 
                           QN => n2002);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => n13, 
                           QN => n2001);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => n14, 
                           QN => n2000);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => n15, 
                           QN => n1999);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => n16, 
                           QN => n1998);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => n17, 
                           QN => n1997);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => n18, 
                           QN => n1996);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => n19, 
                           QN => n1995);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => n20, 
                           QN => n1994);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => n21, 
                           QN => n1993);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => n22, 
                           QN => n1992);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => n23, 
                           QN => n1991);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => n24, 
                           QN => n1990);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => n25, 
                           QN => n1989);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => n26, 
                           QN => n1988);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n27, 
                           QN => n1987);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => n28, 
                           QN => n1986);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n29, 
                           QN => n1985);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => n30, 
                           QN => n1984);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n31, 
                           QN => n1983);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => n32, 
                           QN => n1982);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n33, 
                           QN => n1981);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => n34, 
                           QN => n1980);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n35, 
                           QN => n1979);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => n36, 
                           QN => n1978);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => n37, 
                           QN => n1977);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => n38, 
                           QN => n1976);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => n39, 
                           QN => n1975);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => n40, 
                           QN => n1974);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => n41, 
                           QN => n1973);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => n42, 
                           QN => n1972);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => n43, 
                           QN => n1971);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => n44, 
                           QN => n1970);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => n45, 
                           QN => n1969);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => n46, 
                           QN => n1968);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => n47, 
                           QN => n1967);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => n48, 
                           QN => n1966);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => n49, 
                           QN => n1965);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => n50, 
                           QN => n1964);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => n51, 
                           QN => n1963);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => n52, 
                           QN => n1962);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => n53, 
                           QN => n1961);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => n54, 
                           QN => n1960);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n55, 
                           QN => n1959);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => n56, 
                           QN => n1958);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n57, 
                           QN => n1957);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => n58, 
                           QN => n1956);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n59, 
                           QN => n1955);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => n60, 
                           QN => n1954);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n61, 
                           QN => n1953);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => n62, 
                           QN => n1952);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n63, 
                           QN => n1951);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => n64, 
                           QN => n1950);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n999,
                           QN => n728);
   OUT2_reg_63_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => OUT2(63), QN
                           => n1822);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n1000
                           , QN => n725);
   OUT2_reg_62_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => OUT2(62), QN
                           => n1823);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n1001
                           , QN => n722);
   OUT2_reg_61_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => OUT2(61), QN
                           => n1824);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n1002
                           , QN => n719);
   OUT2_reg_60_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => OUT2(60), QN
                           => n1825);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n1003
                           , QN => n716);
   OUT2_reg_59_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => OUT2(59), QN
                           => n1826);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n1004
                           , QN => n713);
   OUT2_reg_58_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => OUT2(58), QN
                           => n1827);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n1005
                           , QN => n710);
   OUT2_reg_57_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => OUT2(57), QN
                           => n1828);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n1006
                           , QN => n707);
   OUT2_reg_56_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => OUT2(56), QN
                           => n1829);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n1007
                           , QN => n704);
   OUT2_reg_55_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => OUT2(55), QN
                           => n1830);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n1008
                           , QN => n700);
   OUT2_reg_54_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => OUT2(54), QN
                           => n1831);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n1009
                           , QN => n696);
   OUT2_reg_53_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => OUT2(53), QN
                           => n1832);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n1010
                           , QN => n692);
   OUT2_reg_52_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => OUT2(52), QN
                           => n1833);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n1011
                           , QN => n689);
   OUT2_reg_51_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => OUT2(51), QN
                           => n1834);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n1012
                           , QN => n686);
   OUT2_reg_50_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => OUT2(50), QN
                           => n1835);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n1013
                           , QN => n683);
   OUT2_reg_49_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => OUT2(49), QN
                           => n1836);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n1014
                           , QN => n680);
   OUT2_reg_48_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => OUT2(48), QN
                           => n1837);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n1015
                           , QN => n677);
   OUT2_reg_47_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => OUT2(47), QN
                           => n1838);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n1016
                           , QN => n674);
   OUT2_reg_46_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => OUT2(46), QN
                           => n1839);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n1017
                           , QN => n671);
   OUT2_reg_45_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => OUT2(45), QN
                           => n1840);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n1018
                           , QN => n668);
   OUT2_reg_44_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => OUT2(44), QN
                           => n1841);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n1019
                           , QN => n665);
   OUT2_reg_43_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => OUT2(43), QN
                           => n1842);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n1020
                           , QN => n662);
   OUT2_reg_42_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => OUT2(42), QN
                           => n1843);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n1021
                           , QN => n659);
   OUT2_reg_41_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => OUT2(41), QN
                           => n1844);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n1022
                           , QN => n656);
   OUT2_reg_40_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => OUT2(40), QN
                           => n1845);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n1023
                           , QN => n653);
   OUT2_reg_39_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => OUT2(39), QN
                           => n1846);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n1024
                           , QN => n650);
   OUT2_reg_38_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => OUT2(38), QN
                           => n1847);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n1025
                           , QN => n647);
   OUT2_reg_37_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => OUT2(37), QN
                           => n1848);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n1026
                           , QN => n644);
   OUT2_reg_36_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => OUT2(36), QN
                           => n1849);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n1027
                           , QN => n641);
   OUT2_reg_35_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => OUT2(35), QN
                           => n1850);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n1028
                           , QN => n638);
   OUT2_reg_34_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => OUT2(34), QN
                           => n1851);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n1029
                           , QN => n635);
   OUT2_reg_33_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => OUT2(33), QN
                           => n1852);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n1030
                           , QN => n632);
   OUT2_reg_32_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => OUT2(32), QN
                           => n1853);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n1031
                           , QN => n629);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => OUT2(31), QN
                           => n1854);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n1032
                           , QN => n626);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => OUT2(30), QN
                           => n1855);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n1033
                           , QN => n623);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => OUT2(29), QN
                           => n1856);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n1034
                           , QN => n619);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => OUT2(28), QN
                           => n1857);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n1035
                           , QN => n615);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => OUT2(27), QN
                           => n1858);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n1036
                           , QN => n611);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => OUT2(26), QN
                           => n1859);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n1037
                           , QN => n607);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => OUT2(25), QN
                           => n1860);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n1038
                           , QN => n603);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => OUT2(24), QN
                           => n1861);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n1039
                           , QN => n599);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => OUT2(23), QN
                           => n1862);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n1040
                           , QN => n595);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => OUT2(22), QN
                           => n1863);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n1041
                           , QN => n591);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => OUT2(21), QN
                           => n1864);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n1042
                           , QN => n587);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => OUT2(20), QN
                           => n1865);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n1043
                           , QN => n583);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => OUT2(19), QN
                           => n1866);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n1044
                           , QN => n580);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => OUT2(18), QN
                           => n1867);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n1045
                           , QN => n577);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => OUT2(17), QN
                           => n1868);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n1046
                           , QN => n574);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => OUT2(16), QN
                           => n1869);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n1047
                           , QN => n571);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => OUT2(15), QN
                           => n1870);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n1048
                           , QN => n568);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => OUT2(14), QN
                           => n1871);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n1049
                           , QN => n565);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => OUT2(13), QN
                           => n1872);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n1050
                           , QN => n562);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => OUT2(12), QN
                           => n1873);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n1051
                           , QN => n559);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => OUT2(11), QN
                           => n1874);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n1052
                           , QN => n556);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => OUT2(10), QN
                           => n1875);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n1053,
                           QN => n553);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => OUT2(9), QN 
                           => n1876);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => n1054,
                           QN => n550);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => OUT2(8), QN 
                           => n1877);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => n1055,
                           QN => n547);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => OUT2(7), QN 
                           => n1878);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => n1056,
                           QN => n544);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => OUT2(6), QN 
                           => n1879);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => n1057,
                           QN => n541);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => OUT2(5), QN 
                           => n1880);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => n1058,
                           QN => n538);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => OUT2(4), QN 
                           => n1881);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => n1059,
                           QN => n535);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => OUT2(3), QN 
                           => n1882);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n1060,
                           QN => n532);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => OUT2(2), QN 
                           => n1883);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n1061,
                           QN => n529);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => OUT2(1), QN 
                           => n1884);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n1062,
                           QN => n522);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => OUT2(0), QN 
                           => n1885);
   OUT1_reg_63_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => OUT1(63), QN
                           => n1886);
   OUT1_reg_62_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => OUT1(62), QN
                           => n1887);
   OUT1_reg_61_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => OUT1(61), QN
                           => n1888);
   OUT1_reg_60_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => OUT1(60), QN
                           => n1889);
   OUT1_reg_59_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => OUT1(59), QN
                           => n1890);
   OUT1_reg_58_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => OUT1(58), QN
                           => n1891);
   OUT1_reg_57_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => OUT1(57), QN
                           => n1892);
   OUT1_reg_56_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => OUT1(56), QN
                           => n1893);
   OUT1_reg_55_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => OUT1(55), QN
                           => n1894);
   OUT1_reg_54_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => OUT1(54), QN
                           => n1895);
   OUT1_reg_53_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => OUT1(53), QN
                           => n1896);
   OUT1_reg_52_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => OUT1(52), QN
                           => n1897);
   OUT1_reg_51_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => OUT1(51), QN
                           => n1898);
   OUT1_reg_50_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => OUT1(50), QN
                           => n1899);
   OUT1_reg_49_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => OUT1(49), QN
                           => n1900);
   OUT1_reg_48_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => OUT1(48), QN
                           => n1901);
   OUT1_reg_47_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => OUT1(47), QN
                           => n1902);
   OUT1_reg_46_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => OUT1(46), QN
                           => n1903);
   OUT1_reg_45_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => OUT1(45), QN
                           => n1904);
   OUT1_reg_44_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => OUT1(44), QN
                           => n1905);
   OUT1_reg_43_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => OUT1(43), QN
                           => n1906);
   OUT1_reg_42_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => OUT1(42), QN
                           => n1907);
   OUT1_reg_41_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => OUT1(41), QN
                           => n1908);
   OUT1_reg_40_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => OUT1(40), QN
                           => n1909);
   OUT1_reg_39_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => OUT1(39), QN
                           => n1910);
   OUT1_reg_38_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => OUT1(38), QN
                           => n1911);
   OUT1_reg_37_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => OUT1(37), QN
                           => n1912);
   OUT1_reg_36_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => OUT1(36), QN
                           => n1913);
   OUT1_reg_35_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => OUT1(35), QN
                           => n1914);
   OUT1_reg_34_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => OUT1(34), QN
                           => n1915);
   OUT1_reg_33_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => OUT1(33), QN
                           => n1916);
   OUT1_reg_32_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => OUT1(32), QN
                           => n1917);
   OUT1_reg_31_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => OUT1(31), QN
                           => n1918);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => OUT1(30), QN
                           => n1919);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => OUT1(29), QN
                           => n1920);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => OUT1(28), QN
                           => n1921);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => OUT1(27), QN
                           => n1922);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => OUT1(26), QN
                           => n1923);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => OUT1(25), QN
                           => n1924);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => OUT1(24), QN
                           => n1925);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => OUT1(23), QN
                           => n1926);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => OUT1(22), QN
                           => n1927);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => OUT1(21), QN
                           => n1928);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => OUT1(20), QN
                           => n1929);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => OUT1(19), QN
                           => n1930);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => OUT1(18), QN
                           => n1931);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => OUT1(17), QN
                           => n1932);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => OUT1(16), QN
                           => n1933);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => OUT1(15), QN
                           => n1934);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => OUT1(14), QN
                           => n1935);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => OUT1(13), QN
                           => n1936);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => OUT1(12), QN
                           => n1937);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => OUT1(11), QN
                           => n1938);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => OUT1(10), QN
                           => n1939);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => OUT1(9), QN 
                           => n1940);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => OUT1(8), QN 
                           => n1941);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => OUT1(7), QN 
                           => n1942);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => OUT1(6), QN 
                           => n1943);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => OUT1(5), QN 
                           => n1944);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => OUT1(4), QN 
                           => n1945);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => OUT1(3), QN 
                           => n1946);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => OUT1(2), QN 
                           => n1947);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => OUT1(1), QN 
                           => n1948);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => OUT1(0), QN 
                           => n1949);
   U859 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n2164, A3 => ADD_RD1(1), 
                           ZN => n521);
   U860 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n2135, A3 => ADD_RD2(1), 
                           ZN => n735);
   U861 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n873, A3 => ADD_WR(1), ZN 
                           => n872);
   U862 : NAND3_X1 port map( A1 => n873, A2 => n2175, A3 => ADD_WR(1), ZN => 
                           n936);
   U863 : NAND3_X1 port map( A1 => n873, A2 => n2176, A3 => ADD_WR(0), ZN => 
                           n975);
   U864 : NAND3_X1 port map( A1 => n2175, A2 => n2176, A3 => n873, ZN => n998);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => n537, 
                           QN => n1818);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => n534, 
                           QN => n1819);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => n531, 
                           QN => n1820);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => n528, 
                           QN => n1821);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => n730,
                           QN => n415);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => n702,
                           QN => n1200);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => n698,
                           QN => n1202);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => n694,
                           QN => n1204);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => n622,
                           QN => n1793);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => n618,
                           QN => n1794);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => n614,
                           QN => n1795);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => n610,
                           QN => n1796);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => n606,
                           QN => n1797);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => n602,
                           QN => n1798);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => n598,
                           QN => n1799);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => n594,
                           QN => n1800);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => n590,
                           QN => n1801);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => n586,
                           QN => n1802);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => n582,
                           QN => n1803);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => n579,
                           QN => n1804);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => n576,
                           QN => n1805);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => n573,
                           QN => n1806);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => n570,
                           QN => n1807);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => n567,
                           QN => n1808);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => n564,
                           QN => n1809);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => n561,
                           QN => n1810);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => n558,
                           QN => n1811);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => n555, 
                           QN => n1812);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => n552, 
                           QN => n1813);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => n549, 
                           QN => n1814);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => n546, 
                           QN => n1815);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => n543, 
                           QN => n1816);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => n540, 
                           QN => n1817);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => n731,
                           QN => n1694);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => n727,
                           QN => n1695);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => n724,
                           QN => n1696);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => n721,
                           QN => n1697);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => n718,
                           QN => n1698);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => n715,
                           QN => n1699);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => n712,
                           QN => n1700);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => n709,
                           QN => n1701);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => n706,
                           QN => n1702);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => n703,
                           QN => n1703);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => n699,
                           QN => n1704);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => n695,
                           QN => n1705);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => n691,
                           QN => n1706);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => n688,
                           QN => n1707);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => n685,
                           QN => n1708);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => n682,
                           QN => n1709);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => n679,
                           QN => n1710);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => n676,
                           QN => n1711);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => n673,
                           QN => n1712);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => n670,
                           QN => n1713);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => n667,
                           QN => n1714);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => n664,
                           QN => n1715);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => n661,
                           QN => n1716);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => n658,
                           QN => n1717);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => n655,
                           QN => n1718);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => n652,
                           QN => n1719);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => n649,
                           QN => n1720);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => n646,
                           QN => n1721);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => n643,
                           QN => n1722);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => n640,
                           QN => n1723);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => n637,
                           QN => n1724);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => n634,
                           QN => n1725);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => n631,
                           QN => n1726);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => n628,
                           QN => n1727);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n625,
                           QN => n1728);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => n621,
                           QN => n1729);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => n617,
                           QN => n1730);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => n613,
                           QN => n1731);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => n609,
                           QN => n1732);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => n605,
                           QN => n1733);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => n601,
                           QN => n1734);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => n597,
                           QN => n1735);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => n593,
                           QN => n1736);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => n589,
                           QN => n1737);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => n585,
                           QN => n1738);
   U3 : BUF_X1 port map( A => n521, Z => n2167);
   U4 : BUF_X1 port map( A => n521, Z => n2166);
   U5 : BUF_X1 port map( A => n521, Z => n2165);
   U6 : BUF_X1 port map( A => n735, Z => n2139);
   U7 : BUF_X1 port map( A => n735, Z => n2138);
   U8 : BUF_X1 port map( A => n735, Z => n2137);
   U9 : BUF_X1 port map( A => n735, Z => n2136);
   U10 : BUF_X1 port map( A => n521, Z => n2169);
   U11 : BUF_X1 port map( A => n521, Z => n2168);
   U12 : BUF_X1 port map( A => n735, Z => n2140);
   U13 : BUF_X1 port map( A => n526, Z => n2151);
   U14 : BUF_X1 port map( A => n526, Z => n2152);
   U15 : BUF_X1 port map( A => n527, Z => n2144);
   U16 : BUF_X1 port map( A => n527, Z => n2146);
   U17 : BUF_X1 port map( A => n527, Z => n2145);
   U18 : BUF_X1 port map( A => n523, Z => n2159);
   U19 : BUF_X1 port map( A => n523, Z => n2160);
   U20 : BUF_X1 port map( A => n523, Z => n2161);
   U21 : BUF_X1 port map( A => n523, Z => n2162);
   U22 : BUF_X1 port map( A => n523, Z => n2163);
   U23 : BUF_X1 port map( A => n736, Z => n2130);
   U24 : BUF_X1 port map( A => n736, Z => n2131);
   U25 : BUF_X1 port map( A => n736, Z => n2132);
   U26 : BUF_X1 port map( A => n736, Z => n2133);
   U27 : BUF_X1 port map( A => n736, Z => n2134);
   U28 : BUF_X1 port map( A => n525, Z => n2154);
   U29 : BUF_X1 port map( A => n525, Z => n2155);
   U30 : BUF_X1 port map( A => n525, Z => n2156);
   U31 : BUF_X1 port map( A => n525, Z => n2157);
   U32 : BUF_X1 port map( A => n738, Z => n2128);
   U33 : BUF_X1 port map( A => n738, Z => n2127);
   U34 : BUF_X1 port map( A => n738, Z => n2126);
   U35 : BUF_X1 port map( A => n738, Z => n2125);
   U36 : BUF_X1 port map( A => n738, Z => n2124);
   U37 : BUF_X1 port map( A => n742, Z => n2104);
   U38 : BUF_X1 port map( A => n742, Z => n2103);
   U39 : BUF_X1 port map( A => n742, Z => n2102);
   U40 : BUF_X1 port map( A => n742, Z => n2101);
   U41 : BUF_X1 port map( A => n739, Z => n2122);
   U42 : BUF_X1 port map( A => n739, Z => n2121);
   U43 : BUF_X1 port map( A => n739, Z => n2120);
   U44 : BUF_X1 port map( A => n739, Z => n2119);
   U45 : BUF_X1 port map( A => n739, Z => n2118);
   U46 : BUF_X1 port map( A => n740, Z => n2116);
   U47 : BUF_X1 port map( A => n740, Z => n2115);
   U48 : BUF_X1 port map( A => n740, Z => n2114);
   U49 : BUF_X1 port map( A => n740, Z => n2113);
   U50 : BUF_X1 port map( A => n740, Z => n2112);
   U51 : BUF_X1 port map( A => n741, Z => n2106);
   U52 : BUF_X1 port map( A => n875, Z => n2094);
   U53 : BUF_X1 port map( A => n938, Z => n2082);
   U54 : BUF_X1 port map( A => n978, Z => n2070);
   U55 : BUF_X1 port map( A => n741, Z => n2110);
   U56 : BUF_X1 port map( A => n741, Z => n2109);
   U57 : BUF_X1 port map( A => n741, Z => n2108);
   U58 : BUF_X1 port map( A => n741, Z => n2107);
   U59 : BUF_X1 port map( A => n875, Z => n2098);
   U60 : BUF_X1 port map( A => n875, Z => n2097);
   U61 : BUF_X1 port map( A => n875, Z => n2096);
   U62 : BUF_X1 port map( A => n875, Z => n2095);
   U63 : BUF_X1 port map( A => n938, Z => n2086);
   U64 : BUF_X1 port map( A => n938, Z => n2085);
   U65 : BUF_X1 port map( A => n938, Z => n2084);
   U66 : BUF_X1 port map( A => n938, Z => n2083);
   U67 : BUF_X1 port map( A => n978, Z => n2074);
   U68 : BUF_X1 port map( A => n978, Z => n2073);
   U69 : BUF_X1 port map( A => n978, Z => n2072);
   U70 : BUF_X1 port map( A => n978, Z => n2071);
   U71 : BUF_X1 port map( A => n526, Z => n2148);
   U72 : BUF_X1 port map( A => n526, Z => n2150);
   U73 : BUF_X1 port map( A => n876, Z => n2092);
   U74 : BUF_X1 port map( A => n876, Z => n2091);
   U75 : BUF_X1 port map( A => n876, Z => n2090);
   U76 : BUF_X1 port map( A => n876, Z => n2089);
   U77 : BUF_X1 port map( A => n876, Z => n2088);
   U78 : BUF_X1 port map( A => n939, Z => n2080);
   U79 : BUF_X1 port map( A => n939, Z => n2079);
   U80 : BUF_X1 port map( A => n939, Z => n2078);
   U81 : BUF_X1 port map( A => n939, Z => n2077);
   U82 : BUF_X1 port map( A => n939, Z => n2076);
   U83 : BUF_X1 port map( A => n979, Z => n2068);
   U84 : BUF_X1 port map( A => n979, Z => n2067);
   U85 : BUF_X1 port map( A => n979, Z => n2066);
   U86 : BUF_X1 port map( A => n979, Z => n2065);
   U87 : BUF_X1 port map( A => n979, Z => n2064);
   U88 : BUF_X1 port map( A => n527, Z => n2143);
   U89 : BUF_X1 port map( A => n527, Z => n2142);
   U90 : BUF_X1 port map( A => n526, Z => n2149);
   U91 : BUF_X1 port map( A => n525, Z => n2153);
   U92 : BUF_X1 port map( A => n742, Z => n2100);
   U93 : NAND2_X1 port map( A1 => n734, A2 => n872, ZN => n741);
   U94 : NAND2_X1 port map( A1 => n734, A2 => n936, ZN => n875);
   U95 : NAND2_X1 port map( A1 => n734, A2 => n2094, ZN => n876);
   U96 : NAND2_X1 port map( A1 => n734, A2 => n975, ZN => n938);
   U97 : NAND2_X1 port map( A1 => n734, A2 => n2082, ZN => n939);
   U98 : NAND2_X1 port map( A1 => n734, A2 => n998, ZN => n978);
   U99 : NAND2_X1 port map( A1 => n734, A2 => n2070, ZN => n979);
   U100 : OAI22_X1 port map( A1 => n538, A2 => n2111, B1 => n2104, B2 => n751, 
                           ZN => n1620);
   U101 : OAI22_X1 port map( A1 => n541, A2 => n2110, B1 => n2104, B2 => n753, 
                           ZN => n1618);
   U102 : OAI22_X1 port map( A1 => n544, A2 => n2110, B1 => n2104, B2 => n755, 
                           ZN => n1616);
   U103 : OAI22_X1 port map( A1 => n547, A2 => n2110, B1 => n2104, B2 => n757, 
                           ZN => n1614);
   U104 : OAI22_X1 port map( A1 => n550, A2 => n2110, B1 => n2104, B2 => n759, 
                           ZN => n1612);
   U105 : OAI22_X1 port map( A1 => n553, A2 => n2110, B1 => n2104, B2 => n761, 
                           ZN => n1610);
   U106 : OAI22_X1 port map( A1 => n556, A2 => n2110, B1 => n2104, B2 => n763, 
                           ZN => n1608);
   U107 : OAI22_X1 port map( A1 => n559, A2 => n2110, B1 => n2104, B2 => n765, 
                           ZN => n1606);
   U108 : OAI22_X1 port map( A1 => n562, A2 => n2110, B1 => n2104, B2 => n767, 
                           ZN => n1604);
   U109 : OAI22_X1 port map( A1 => n565, A2 => n2110, B1 => n2104, B2 => n769, 
                           ZN => n1602);
   U110 : OAI22_X1 port map( A1 => n568, A2 => n2110, B1 => n2104, B2 => n771, 
                           ZN => n1600);
   U111 : OAI22_X1 port map( A1 => n571, A2 => n2110, B1 => n2104, B2 => n773, 
                           ZN => n1598);
   U112 : OAI22_X1 port map( A1 => n574, A2 => n2110, B1 => n2103, B2 => n775, 
                           ZN => n1596);
   U113 : OAI22_X1 port map( A1 => n577, A2 => n2109, B1 => n2103, B2 => n777, 
                           ZN => n1594);
   U114 : OAI22_X1 port map( A1 => n580, A2 => n2109, B1 => n2103, B2 => n779, 
                           ZN => n1592);
   U115 : OAI22_X1 port map( A1 => n583, A2 => n2109, B1 => n2103, B2 => n781, 
                           ZN => n1590);
   U116 : OAI22_X1 port map( A1 => n587, A2 => n2109, B1 => n2103, B2 => n783, 
                           ZN => n1588);
   U117 : OAI22_X1 port map( A1 => n591, A2 => n2109, B1 => n2103, B2 => n785, 
                           ZN => n1586);
   U118 : OAI22_X1 port map( A1 => n595, A2 => n2109, B1 => n2103, B2 => n787, 
                           ZN => n1584);
   U119 : OAI22_X1 port map( A1 => n599, A2 => n2109, B1 => n2103, B2 => n789, 
                           ZN => n1582);
   U120 : OAI22_X1 port map( A1 => n603, A2 => n2109, B1 => n2103, B2 => n791, 
                           ZN => n1580);
   U121 : OAI22_X1 port map( A1 => n607, A2 => n2109, B1 => n2103, B2 => n793, 
                           ZN => n1578);
   U122 : OAI22_X1 port map( A1 => n611, A2 => n2109, B1 => n2103, B2 => n795, 
                           ZN => n1576);
   U123 : OAI22_X1 port map( A1 => n615, A2 => n2109, B1 => n2103, B2 => n797, 
                           ZN => n1574);
   U124 : OAI22_X1 port map( A1 => n619, A2 => n2109, B1 => n2102, B2 => n799, 
                           ZN => n1572);
   U125 : OAI22_X1 port map( A1 => n623, A2 => n2108, B1 => n2102, B2 => n801, 
                           ZN => n1570);
   U126 : OAI22_X1 port map( A1 => n626, A2 => n2108, B1 => n2102, B2 => n803, 
                           ZN => n1568);
   U127 : OAI22_X1 port map( A1 => n629, A2 => n2108, B1 => n2102, B2 => n805, 
                           ZN => n1566);
   U128 : OAI22_X1 port map( A1 => n632, A2 => n2108, B1 => n2102, B2 => n807, 
                           ZN => n1564);
   U129 : OAI22_X1 port map( A1 => n635, A2 => n2108, B1 => n2102, B2 => n809, 
                           ZN => n1562);
   U130 : OAI22_X1 port map( A1 => n638, A2 => n2108, B1 => n2102, B2 => n811, 
                           ZN => n1560);
   U131 : OAI22_X1 port map( A1 => n641, A2 => n2108, B1 => n2102, B2 => n813, 
                           ZN => n1558);
   U132 : OAI22_X1 port map( A1 => n644, A2 => n2108, B1 => n2102, B2 => n815, 
                           ZN => n1556);
   U133 : OAI22_X1 port map( A1 => n647, A2 => n2108, B1 => n2102, B2 => n817, 
                           ZN => n1554);
   U134 : OAI22_X1 port map( A1 => n650, A2 => n2108, B1 => n2102, B2 => n819, 
                           ZN => n1552);
   U135 : OAI22_X1 port map( A1 => n653, A2 => n2108, B1 => n2102, B2 => n821, 
                           ZN => n1550);
   U136 : OAI22_X1 port map( A1 => n656, A2 => n2108, B1 => n2101, B2 => n823, 
                           ZN => n1548);
   U137 : OAI22_X1 port map( A1 => n659, A2 => n2107, B1 => n2101, B2 => n825, 
                           ZN => n1546);
   U138 : OAI22_X1 port map( A1 => n662, A2 => n2107, B1 => n2101, B2 => n827, 
                           ZN => n1544);
   U139 : OAI22_X1 port map( A1 => n665, A2 => n2107, B1 => n2101, B2 => n829, 
                           ZN => n1542);
   U140 : OAI22_X1 port map( A1 => n668, A2 => n2107, B1 => n2101, B2 => n831, 
                           ZN => n1540);
   U141 : OAI22_X1 port map( A1 => n671, A2 => n2107, B1 => n2101, B2 => n833, 
                           ZN => n1538);
   U142 : OAI22_X1 port map( A1 => n674, A2 => n2107, B1 => n2101, B2 => n835, 
                           ZN => n1536);
   U143 : OAI22_X1 port map( A1 => n677, A2 => n2107, B1 => n2101, B2 => n837, 
                           ZN => n1534);
   U144 : OAI22_X1 port map( A1 => n680, A2 => n2107, B1 => n2101, B2 => n839, 
                           ZN => n1532);
   U145 : OAI22_X1 port map( A1 => n683, A2 => n2107, B1 => n2101, B2 => n841, 
                           ZN => n1530);
   U146 : OAI22_X1 port map( A1 => n686, A2 => n2107, B1 => n2101, B2 => n843, 
                           ZN => n1528);
   U147 : OAI22_X1 port map( A1 => n689, A2 => n2107, B1 => n2101, B2 => n845, 
                           ZN => n1526);
   U148 : OAI22_X1 port map( A1 => n522, A2 => n2111, B1 => n2105, B2 => n743, 
                           ZN => n1628);
   U149 : OAI22_X1 port map( A1 => n529, A2 => n2111, B1 => n2105, B2 => n745, 
                           ZN => n1626);
   U150 : OAI22_X1 port map( A1 => n532, A2 => n2111, B1 => n2105, B2 => n747, 
                           ZN => n1624);
   U151 : OAI22_X1 port map( A1 => n535, A2 => n2111, B1 => n2105, B2 => n749, 
                           ZN => n1622);
   U152 : OAI22_X1 port map( A1 => n692, A2 => n2107, B1 => n2100, B2 => n847, 
                           ZN => n1524);
   U153 : OAI22_X1 port map( A1 => n696, A2 => n2106, B1 => n2100, B2 => n849, 
                           ZN => n1522);
   U154 : OAI22_X1 port map( A1 => n700, A2 => n2106, B1 => n2100, B2 => n851, 
                           ZN => n1520);
   U155 : OAI22_X1 port map( A1 => n704, A2 => n2106, B1 => n2100, B2 => n853, 
                           ZN => n1518);
   U156 : OAI22_X1 port map( A1 => n707, A2 => n2106, B1 => n2100, B2 => n855, 
                           ZN => n1516);
   U157 : OAI22_X1 port map( A1 => n710, A2 => n2106, B1 => n2100, B2 => n857, 
                           ZN => n1514);
   U158 : OAI22_X1 port map( A1 => n713, A2 => n2106, B1 => n2100, B2 => n859, 
                           ZN => n1512);
   U159 : OAI22_X1 port map( A1 => n716, A2 => n2106, B1 => n2100, B2 => n861, 
                           ZN => n1510);
   U160 : OAI22_X1 port map( A1 => n719, A2 => n2106, B1 => n2100, B2 => n863, 
                           ZN => n1508);
   U161 : OAI22_X1 port map( A1 => n722, A2 => n2106, B1 => n2100, B2 => n865, 
                           ZN => n1506);
   U162 : OAI22_X1 port map( A1 => n725, A2 => n2106, B1 => n2100, B2 => n867, 
                           ZN => n1504);
   U163 : OAI22_X1 port map( A1 => n728, A2 => n2106, B1 => n2100, B2 => n871, 
                           ZN => n1502);
   U164 : AND3_X1 port map( A1 => n2173, A2 => n2174, A3 => n2164, ZN => n526);
   U165 : AND3_X1 port map( A1 => n2164, A2 => n2174, A3 => ADD_RD1(0), ZN => 
                           n527);
   U166 : AND3_X1 port map( A1 => n2164, A2 => n2173, A3 => ADD_RD1(1), ZN => 
                           n525);
   U167 : NAND2_X1 port map( A1 => n734, A2 => n2106, ZN => n742);
   U168 : AND3_X1 port map( A1 => n2135, A2 => n2172, A3 => ADD_RD2(0), ZN => 
                           n740);
   U169 : AND3_X1 port map( A1 => n2135, A2 => n2171, A3 => ADD_RD2(1), ZN => 
                           n738);
   U170 : AND3_X1 port map( A1 => n2171, A2 => n2172, A3 => n2135, ZN => n739);
   U171 : AND2_X1 port map( A1 => RD1, A2 => n734, ZN => n523);
   U172 : AND2_X1 port map( A1 => RD2, A2 => n734, ZN => n736);
   U173 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n873);
   U174 : OAI221_X1 port map( B1 => n2169, B2 => n562, C1 => n1937, C2 => n2160
                           , A => n563, ZN => n1681);
   U175 : AOI222_X1 port map( A1 => n52, A2 => n2153, B1 => n180, B2 => n2149, 
                           C1 => n2146, C2 => n564, ZN => n563);
   U176 : OAI221_X1 port map( B1 => n2169, B2 => n565, C1 => n1936, C2 => n2160
                           , A => n566, ZN => n1680);
   U177 : AOI222_X1 port map( A1 => n51, A2 => n2154, B1 => n179, B2 => n2149, 
                           C1 => n2146, C2 => n567, ZN => n566);
   U178 : OAI221_X1 port map( B1 => n2169, B2 => n568, C1 => n1935, C2 => n2160
                           , A => n569, ZN => n1679);
   U179 : AOI222_X1 port map( A1 => n50, A2 => n2154, B1 => n178, B2 => n2149, 
                           C1 => n2146, C2 => n570, ZN => n569);
   U180 : OAI221_X1 port map( B1 => n2169, B2 => n571, C1 => n1934, C2 => n2161
                           , A => n572, ZN => n1678);
   U181 : AOI222_X1 port map( A1 => n49, A2 => n2154, B1 => n177, B2 => n2149, 
                           C1 => n2145, C2 => n573, ZN => n572);
   U182 : OAI221_X1 port map( B1 => n2168, B2 => n574, C1 => n1933, C2 => n2160
                           , A => n575, ZN => n1677);
   U183 : AOI222_X1 port map( A1 => n48, A2 => n2154, B1 => n176, B2 => n2149, 
                           C1 => n2145, C2 => n576, ZN => n575);
   U184 : OAI221_X1 port map( B1 => n2168, B2 => n577, C1 => n1932, C2 => n2160
                           , A => n578, ZN => n1676);
   U185 : AOI222_X1 port map( A1 => n47, A2 => n2154, B1 => n175, B2 => n2149, 
                           C1 => n2145, C2 => n579, ZN => n578);
   U186 : OAI221_X1 port map( B1 => n2168, B2 => n580, C1 => n1931, C2 => n2160
                           , A => n581, ZN => n1675);
   U187 : AOI222_X1 port map( A1 => n46, A2 => n2154, B1 => n174, B2 => n2149, 
                           C1 => n2145, C2 => n582, ZN => n581);
   U188 : OAI221_X1 port map( B1 => n538, B2 => n2140, C1 => n1881, C2 => n2130
                           , A => n750, ZN => n1621);
   U189 : AOI222_X1 port map( A1 => n2128, A2 => n60, B1 => n2122, B2 => n188, 
                           C1 => n2116, C2 => n540, ZN => n750);
   U190 : OAI221_X1 port map( B1 => n541, B2 => n2140, C1 => n1880, C2 => n2130
                           , A => n752, ZN => n1619);
   U191 : AOI222_X1 port map( A1 => n2128, A2 => n59, B1 => n2122, B2 => n187, 
                           C1 => n2116, C2 => n543, ZN => n752);
   U192 : OAI221_X1 port map( B1 => n544, B2 => n2140, C1 => n1879, C2 => n2130
                           , A => n754, ZN => n1617);
   U193 : AOI222_X1 port map( A1 => n2128, A2 => n58, B1 => n2122, B2 => n186, 
                           C1 => n2116, C2 => n546, ZN => n754);
   U194 : OAI221_X1 port map( B1 => n547, B2 => n2140, C1 => n1878, C2 => n2130
                           , A => n756, ZN => n1615);
   U195 : AOI222_X1 port map( A1 => n2128, A2 => n57, B1 => n2122, B2 => n185, 
                           C1 => n2116, C2 => n549, ZN => n756);
   U196 : OAI221_X1 port map( B1 => n550, B2 => n2140, C1 => n1877, C2 => n2130
                           , A => n758, ZN => n1613);
   U197 : AOI222_X1 port map( A1 => n2128, A2 => n56, B1 => n2122, B2 => n184, 
                           C1 => n2116, C2 => n552, ZN => n758);
   U198 : OAI221_X1 port map( B1 => n553, B2 => n2140, C1 => n1876, C2 => n2130
                           , A => n760, ZN => n1611);
   U199 : AOI222_X1 port map( A1 => n2128, A2 => n55, B1 => n2122, B2 => n183, 
                           C1 => n2116, C2 => n555, ZN => n760);
   U200 : OAI221_X1 port map( B1 => n556, B2 => n2140, C1 => n1875, C2 => n2130
                           , A => n762, ZN => n1609);
   U201 : AOI222_X1 port map( A1 => n2128, A2 => n54, B1 => n2122, B2 => n182, 
                           C1 => n2116, C2 => n558, ZN => n762);
   U202 : OAI221_X1 port map( B1 => n559, B2 => n2140, C1 => n1874, C2 => n2130
                           , A => n764, ZN => n1607);
   U203 : AOI222_X1 port map( A1 => n2128, A2 => n53, B1 => n2122, B2 => n181, 
                           C1 => n2116, C2 => n561, ZN => n764);
   U204 : OAI221_X1 port map( B1 => n562, B2 => n2140, C1 => n1873, C2 => n2131
                           , A => n766, ZN => n1605);
   U205 : AOI222_X1 port map( A1 => n2128, A2 => n52, B1 => n2122, B2 => n180, 
                           C1 => n2116, C2 => n564, ZN => n766);
   U206 : OAI221_X1 port map( B1 => n565, B2 => n2140, C1 => n1872, C2 => n2131
                           , A => n768, ZN => n1603);
   U207 : AOI222_X1 port map( A1 => n2128, A2 => n51, B1 => n2122, B2 => n179, 
                           C1 => n2116, C2 => n567, ZN => n768);
   U208 : OAI221_X1 port map( B1 => n568, B2 => n2140, C1 => n1871, C2 => n2131
                           , A => n770, ZN => n1601);
   U209 : AOI222_X1 port map( A1 => n2128, A2 => n50, B1 => n2122, B2 => n178, 
                           C1 => n2116, C2 => n570, ZN => n770);
   U210 : OAI221_X1 port map( B1 => n571, B2 => n2140, C1 => n1870, C2 => n2132
                           , A => n772, ZN => n1599);
   U211 : AOI222_X1 port map( A1 => n2128, A2 => n49, B1 => n2122, B2 => n177, 
                           C1 => n2116, C2 => n573, ZN => n772);
   U212 : OAI221_X1 port map( B1 => n574, B2 => n2139, C1 => n1869, C2 => n2131
                           , A => n774, ZN => n1597);
   U213 : AOI222_X1 port map( A1 => n2127, A2 => n48, B1 => n2121, B2 => n176, 
                           C1 => n2115, C2 => n576, ZN => n774);
   U214 : OAI221_X1 port map( B1 => n577, B2 => n2139, C1 => n1868, C2 => n2131
                           , A => n776, ZN => n1595);
   U215 : AOI222_X1 port map( A1 => n2127, A2 => n47, B1 => n2121, B2 => n175, 
                           C1 => n2115, C2 => n579, ZN => n776);
   U216 : OAI221_X1 port map( B1 => n580, B2 => n2139, C1 => n1867, C2 => n2131
                           , A => n778, ZN => n1593);
   U217 : AOI222_X1 port map( A1 => n2127, A2 => n46, B1 => n2121, B2 => n174, 
                           C1 => n2115, C2 => n582, ZN => n778);
   U218 : OAI221_X1 port map( B1 => n2166, B2 => n656, C1 => n1909, C2 => n2162
                           , A => n657, ZN => n1653);
   U219 : AOI222_X1 port map( A1 => n24, A2 => n2156, B1 => n2151, B2 => n658, 
                           C1 => n88, C2 => n2143, ZN => n657);
   U220 : OAI221_X1 port map( B1 => n2166, B2 => n659, C1 => n1908, C2 => n2162
                           , A => n660, ZN => n1652);
   U221 : AOI222_X1 port map( A1 => n23, A2 => n2156, B1 => n2151, B2 => n661, 
                           C1 => n87, C2 => n2143, ZN => n660);
   U222 : OAI221_X1 port map( B1 => n2166, B2 => n662, C1 => n1907, C2 => n2162
                           , A => n663, ZN => n1651);
   U223 : AOI222_X1 port map( A1 => n22, A2 => n2156, B1 => n2151, B2 => n664, 
                           C1 => n86, C2 => n2143, ZN => n663);
   U224 : OAI221_X1 port map( B1 => n2166, B2 => n665, C1 => n1906, C2 => n2162
                           , A => n666, ZN => n1650);
   U225 : AOI222_X1 port map( A1 => n21, A2 => n2156, B1 => n2151, B2 => n667, 
                           C1 => n85, C2 => n2143, ZN => n666);
   U226 : OAI221_X1 port map( B1 => n2166, B2 => n668, C1 => n1905, C2 => n2162
                           , A => n669, ZN => n1649);
   U227 : AOI222_X1 port map( A1 => n20, A2 => n2156, B1 => n2151, B2 => n670, 
                           C1 => n84, C2 => n2143, ZN => n669);
   U228 : OAI221_X1 port map( B1 => n2166, B2 => n671, C1 => n1904, C2 => n2162
                           , A => n672, ZN => n1648);
   U229 : AOI222_X1 port map( A1 => n19, A2 => n2156, B1 => n2151, B2 => n673, 
                           C1 => n83, C2 => n2143, ZN => n672);
   U230 : OAI221_X1 port map( B1 => n2166, B2 => n674, C1 => n1903, C2 => n2162
                           , A => n675, ZN => n1647);
   U231 : AOI222_X1 port map( A1 => n18, A2 => n2156, B1 => n2151, B2 => n676, 
                           C1 => n82, C2 => n2143, ZN => n675);
   U232 : OAI221_X1 port map( B1 => n2166, B2 => n677, C1 => n1902, C2 => n2162
                           , A => n678, ZN => n1646);
   U233 : AOI222_X1 port map( A1 => n17, A2 => n2156, B1 => n2151, B2 => n679, 
                           C1 => n81, C2 => n2143, ZN => n678);
   U234 : OAI221_X1 port map( B1 => n2166, B2 => n680, C1 => n1901, C2 => n2163
                           , A => n681, ZN => n1645);
   U235 : AOI222_X1 port map( A1 => n16, A2 => n2157, B1 => n2151, B2 => n682, 
                           C1 => n80, C2 => n2143, ZN => n681);
   U236 : OAI221_X1 port map( B1 => n2166, B2 => n683, C1 => n1900, C2 => n2163
                           , A => n684, ZN => n1644);
   U237 : AOI222_X1 port map( A1 => n15, A2 => n2157, B1 => n2151, B2 => n685, 
                           C1 => n79, C2 => n2143, ZN => n684);
   U238 : OAI221_X1 port map( B1 => n2166, B2 => n686, C1 => n1899, C2 => n2163
                           , A => n687, ZN => n1643);
   U239 : AOI222_X1 port map( A1 => n14, A2 => n2157, B1 => n2152, B2 => n688, 
                           C1 => n78, C2 => n2143, ZN => n687);
   U240 : OAI221_X1 port map( B1 => n2166, B2 => n689, C1 => n1898, C2 => n2163
                           , A => n690, ZN => n1642);
   U241 : AOI222_X1 port map( A1 => n13, A2 => n2157, B1 => n2152, B2 => n691, 
                           C1 => n77, C2 => n2143, ZN => n690);
   U242 : OAI221_X1 port map( B1 => n2165, B2 => n692, C1 => n1897, C2 => n2163
                           , A => n693, ZN => n1641);
   U243 : AOI222_X1 port map( A1 => n2158, A2 => n694, B1 => n2152, B2 => n695,
                           C1 => n76, C2 => n2142, ZN => n693);
   U244 : OAI221_X1 port map( B1 => n2165, B2 => n696, C1 => n1896, C2 => n2163
                           , A => n697, ZN => n1640);
   U245 : AOI222_X1 port map( A1 => n2158, A2 => n698, B1 => n2152, B2 => n699,
                           C1 => n75, C2 => n2142, ZN => n697);
   U246 : OAI221_X1 port map( B1 => n2165, B2 => n700, C1 => n1895, C2 => n2163
                           , A => n701, ZN => n1639);
   U247 : AOI222_X1 port map( A1 => n2158, A2 => n702, B1 => n2152, B2 => n703,
                           C1 => n74, C2 => n2142, ZN => n701);
   U248 : OAI221_X1 port map( B1 => n2165, B2 => n704, C1 => n1894, C2 => n2163
                           , A => n705, ZN => n1638);
   U249 : AOI222_X1 port map( A1 => n9, A2 => n2157, B1 => n2152, B2 => n706, 
                           C1 => n73, C2 => n2142, ZN => n705);
   U250 : OAI221_X1 port map( B1 => n2165, B2 => n707, C1 => n1893, C2 => n2163
                           , A => n708, ZN => n1637);
   U251 : AOI222_X1 port map( A1 => n8, A2 => n2157, B1 => n2152, B2 => n709, 
                           C1 => n72, C2 => n2142, ZN => n708);
   U252 : OAI221_X1 port map( B1 => n2165, B2 => n710, C1 => n1892, C2 => n2163
                           , A => n711, ZN => n1636);
   U253 : AOI222_X1 port map( A1 => n7, A2 => n2157, B1 => n2152, B2 => n712, 
                           C1 => n71, C2 => n2142, ZN => n711);
   U254 : OAI221_X1 port map( B1 => n2165, B2 => n713, C1 => n1891, C2 => n2163
                           , A => n714, ZN => n1635);
   U255 : AOI222_X1 port map( A1 => n6, A2 => n2157, B1 => n2152, B2 => n715, 
                           C1 => n70, C2 => n2142, ZN => n714);
   U256 : OAI221_X1 port map( B1 => n2165, B2 => n719, C1 => n1889, C2 => n2163
                           , A => n720, ZN => n1633);
   U257 : AOI222_X1 port map( A1 => n4, A2 => n2157, B1 => n2152, B2 => n721, 
                           C1 => n68, C2 => n2142, ZN => n720);
   U258 : OAI221_X1 port map( B1 => n2165, B2 => n728, C1 => n1886, C2 => n2164
                           , A => n729, ZN => n1630);
   U259 : AOI222_X1 port map( A1 => n2158, A2 => n730, B1 => n2148, B2 => n731,
                           C1 => n65, C2 => n2142, ZN => n729);
   U260 : OAI221_X1 port map( B1 => n623, B2 => n2138, C1 => n1856, C2 => n2132
                           , A => n800, ZN => n1571);
   U261 : AOI222_X1 port map( A1 => n2126, A2 => n35, B1 => n2120, B2 => n625, 
                           C1 => n2114, C2 => n99, ZN => n800);
   U262 : OAI221_X1 port map( B1 => n626, B2 => n2138, C1 => n1855, C2 => n2132
                           , A => n802, ZN => n1569);
   U263 : AOI222_X1 port map( A1 => n2126, A2 => n34, B1 => n2120, B2 => n628, 
                           C1 => n2114, C2 => n98, ZN => n802);
   U264 : OAI221_X1 port map( B1 => n629, B2 => n2138, C1 => n1854, C2 => n2132
                           , A => n804, ZN => n1567);
   U265 : AOI222_X1 port map( A1 => n2126, A2 => n33, B1 => n2120, B2 => n631, 
                           C1 => n2114, C2 => n97, ZN => n804);
   U266 : OAI221_X1 port map( B1 => n632, B2 => n2138, C1 => n1853, C2 => n2132
                           , A => n806, ZN => n1565);
   U267 : AOI222_X1 port map( A1 => n2126, A2 => n32, B1 => n2120, B2 => n634, 
                           C1 => n2114, C2 => n96, ZN => n806);
   U268 : OAI221_X1 port map( B1 => n635, B2 => n2138, C1 => n1852, C2 => n2132
                           , A => n808, ZN => n1563);
   U269 : AOI222_X1 port map( A1 => n2126, A2 => n31, B1 => n2120, B2 => n637, 
                           C1 => n2114, C2 => n95, ZN => n808);
   U270 : OAI221_X1 port map( B1 => n638, B2 => n2138, C1 => n1851, C2 => n2132
                           , A => n810, ZN => n1561);
   U271 : AOI222_X1 port map( A1 => n2126, A2 => n30, B1 => n2120, B2 => n640, 
                           C1 => n2114, C2 => n94, ZN => n810);
   U272 : OAI221_X1 port map( B1 => n641, B2 => n2138, C1 => n1850, C2 => n2132
                           , A => n812, ZN => n1559);
   U273 : AOI222_X1 port map( A1 => n2126, A2 => n29, B1 => n2120, B2 => n643, 
                           C1 => n2114, C2 => n93, ZN => n812);
   U274 : OAI221_X1 port map( B1 => n644, B2 => n2138, C1 => n1849, C2 => n2133
                           , A => n814, ZN => n1557);
   U275 : AOI222_X1 port map( A1 => n2126, A2 => n28, B1 => n2120, B2 => n646, 
                           C1 => n2114, C2 => n92, ZN => n814);
   U276 : OAI221_X1 port map( B1 => n647, B2 => n2138, C1 => n1848, C2 => n2133
                           , A => n816, ZN => n1555);
   U277 : AOI222_X1 port map( A1 => n2126, A2 => n27, B1 => n2120, B2 => n649, 
                           C1 => n2114, C2 => n91, ZN => n816);
   U278 : OAI221_X1 port map( B1 => n650, B2 => n2138, C1 => n1847, C2 => n2133
                           , A => n818, ZN => n1553);
   U279 : AOI222_X1 port map( A1 => n2126, A2 => n26, B1 => n2120, B2 => n652, 
                           C1 => n2114, C2 => n90, ZN => n818);
   U280 : OAI221_X1 port map( B1 => n653, B2 => n2138, C1 => n1846, C2 => n2133
                           , A => n820, ZN => n1551);
   U281 : AOI222_X1 port map( A1 => n2126, A2 => n25, B1 => n2120, B2 => n655, 
                           C1 => n2114, C2 => n89, ZN => n820);
   U282 : OAI221_X1 port map( B1 => n656, B2 => n2137, C1 => n1845, C2 => n2133
                           , A => n822, ZN => n1549);
   U283 : AOI222_X1 port map( A1 => n2125, A2 => n24, B1 => n2119, B2 => n658, 
                           C1 => n2113, C2 => n88, ZN => n822);
   U284 : OAI221_X1 port map( B1 => n659, B2 => n2137, C1 => n1844, C2 => n2133
                           , A => n824, ZN => n1547);
   U285 : AOI222_X1 port map( A1 => n2125, A2 => n23, B1 => n2119, B2 => n661, 
                           C1 => n2113, C2 => n87, ZN => n824);
   U286 : OAI221_X1 port map( B1 => n662, B2 => n2137, C1 => n1843, C2 => n2133
                           , A => n826, ZN => n1545);
   U287 : AOI222_X1 port map( A1 => n2125, A2 => n22, B1 => n2119, B2 => n664, 
                           C1 => n2113, C2 => n86, ZN => n826);
   U288 : OAI221_X1 port map( B1 => n665, B2 => n2137, C1 => n1842, C2 => n2133
                           , A => n828, ZN => n1543);
   U289 : AOI222_X1 port map( A1 => n2125, A2 => n21, B1 => n2119, B2 => n667, 
                           C1 => n2113, C2 => n85, ZN => n828);
   U290 : OAI221_X1 port map( B1 => n668, B2 => n2137, C1 => n1841, C2 => n2133
                           , A => n830, ZN => n1541);
   U291 : AOI222_X1 port map( A1 => n2125, A2 => n20, B1 => n2119, B2 => n670, 
                           C1 => n2113, C2 => n84, ZN => n830);
   U292 : OAI221_X1 port map( B1 => n671, B2 => n2137, C1 => n1840, C2 => n2133
                           , A => n832, ZN => n1539);
   U293 : AOI222_X1 port map( A1 => n2125, A2 => n19, B1 => n2119, B2 => n673, 
                           C1 => n2113, C2 => n83, ZN => n832);
   U294 : OAI221_X1 port map( B1 => n674, B2 => n2137, C1 => n1839, C2 => n2133
                           , A => n834, ZN => n1537);
   U295 : AOI222_X1 port map( A1 => n2125, A2 => n18, B1 => n2119, B2 => n676, 
                           C1 => n2113, C2 => n82, ZN => n834);
   U296 : OAI221_X1 port map( B1 => n677, B2 => n2137, C1 => n1838, C2 => n2133
                           , A => n836, ZN => n1535);
   U297 : AOI222_X1 port map( A1 => n2125, A2 => n17, B1 => n2119, B2 => n679, 
                           C1 => n2113, C2 => n81, ZN => n836);
   U298 : OAI221_X1 port map( B1 => n680, B2 => n2137, C1 => n1837, C2 => n2134
                           , A => n838, ZN => n1533);
   U299 : AOI222_X1 port map( A1 => n2125, A2 => n16, B1 => n2119, B2 => n682, 
                           C1 => n2113, C2 => n80, ZN => n838);
   U300 : OAI221_X1 port map( B1 => n683, B2 => n2137, C1 => n1836, C2 => n2134
                           , A => n840, ZN => n1531);
   U301 : AOI222_X1 port map( A1 => n2125, A2 => n15, B1 => n2119, B2 => n685, 
                           C1 => n2113, C2 => n79, ZN => n840);
   U302 : OAI221_X1 port map( B1 => n686, B2 => n2137, C1 => n1835, C2 => n2134
                           , A => n842, ZN => n1529);
   U303 : AOI222_X1 port map( A1 => n2125, A2 => n14, B1 => n2119, B2 => n688, 
                           C1 => n2113, C2 => n78, ZN => n842);
   U304 : OAI221_X1 port map( B1 => n689, B2 => n2137, C1 => n1834, C2 => n2134
                           , A => n844, ZN => n1527);
   U305 : AOI222_X1 port map( A1 => n2125, A2 => n13, B1 => n2119, B2 => n691, 
                           C1 => n2113, C2 => n77, ZN => n844);
   U306 : OAI221_X1 port map( B1 => n692, B2 => n2136, C1 => n1833, C2 => n2134
                           , A => n846, ZN => n1525);
   U307 : AOI222_X1 port map( A1 => n2124, A2 => n694, B1 => n2118, B2 => n695,
                           C1 => n2112, C2 => n76, ZN => n846);
   U308 : OAI221_X1 port map( B1 => n696, B2 => n2136, C1 => n1832, C2 => n2134
                           , A => n848, ZN => n1523);
   U309 : AOI222_X1 port map( A1 => n2124, A2 => n698, B1 => n2118, B2 => n699,
                           C1 => n2112, C2 => n75, ZN => n848);
   U310 : OAI221_X1 port map( B1 => n700, B2 => n2136, C1 => n1831, C2 => n2134
                           , A => n850, ZN => n1521);
   U311 : AOI222_X1 port map( A1 => n2124, A2 => n702, B1 => n2118, B2 => n703,
                           C1 => n2112, C2 => n74, ZN => n850);
   U312 : OAI221_X1 port map( B1 => n704, B2 => n2136, C1 => n1830, C2 => n2134
                           , A => n852, ZN => n1519);
   U313 : AOI222_X1 port map( A1 => n2124, A2 => n9, B1 => n2118, B2 => n706, 
                           C1 => n2112, C2 => n73, ZN => n852);
   U314 : OAI221_X1 port map( B1 => n707, B2 => n2136, C1 => n1829, C2 => n2134
                           , A => n854, ZN => n1517);
   U315 : AOI222_X1 port map( A1 => n2124, A2 => n8, B1 => n2118, B2 => n709, 
                           C1 => n2112, C2 => n72, ZN => n854);
   U316 : OAI221_X1 port map( B1 => n710, B2 => n2136, C1 => n1828, C2 => n2134
                           , A => n856, ZN => n1515);
   U317 : AOI222_X1 port map( A1 => n2124, A2 => n7, B1 => n2118, B2 => n712, 
                           C1 => n2112, C2 => n71, ZN => n856);
   U318 : OAI221_X1 port map( B1 => n713, B2 => n2136, C1 => n1827, C2 => n2134
                           , A => n858, ZN => n1513);
   U319 : AOI222_X1 port map( A1 => n2124, A2 => n6, B1 => n2118, B2 => n715, 
                           C1 => n2112, C2 => n70, ZN => n858);
   U320 : OAI221_X1 port map( B1 => n716, B2 => n2136, C1 => n1826, C2 => n2135
                           , A => n860, ZN => n1511);
   U321 : AOI222_X1 port map( A1 => n2124, A2 => n5, B1 => n2118, B2 => n718, 
                           C1 => n2112, C2 => n69, ZN => n860);
   U322 : OAI221_X1 port map( B1 => n719, B2 => n2136, C1 => n1825, C2 => n2134
                           , A => n862, ZN => n1509);
   U323 : AOI222_X1 port map( A1 => n2124, A2 => n4, B1 => n2118, B2 => n721, 
                           C1 => n2112, C2 => n68, ZN => n862);
   U324 : OAI221_X1 port map( B1 => n722, B2 => n2136, C1 => n1824, C2 => n2135
                           , A => n864, ZN => n1507);
   U325 : AOI222_X1 port map( A1 => n2124, A2 => n3, B1 => n2118, B2 => n724, 
                           C1 => n2112, C2 => n67, ZN => n864);
   U326 : OAI221_X1 port map( B1 => n725, B2 => n2136, C1 => n1823, C2 => n2135
                           , A => n866, ZN => n1505);
   U327 : AOI222_X1 port map( A1 => n2124, A2 => n2, B1 => n2118, B2 => n727, 
                           C1 => n2112, C2 => n66, ZN => n866);
   U328 : OAI221_X1 port map( B1 => n728, B2 => n2136, C1 => n1822, C2 => n2135
                           , A => n868, ZN => n1503);
   U329 : AOI222_X1 port map( A1 => n2124, A2 => n730, B1 => n2118, B2 => n731,
                           C1 => n2112, C2 => n65, ZN => n868);
   U330 : INV_X1 port map( A => RESET, ZN => n734);
   U331 : OAI221_X1 port map( B1 => n2170, B2 => n522, C1 => n1949, C2 => n2159
                           , A => n524, ZN => n1693);
   U332 : AOI222_X1 port map( A1 => n64, A2 => n2155, B1 => n192, B2 => n2148, 
                           C1 => n2147, C2 => n528, ZN => n524);
   U333 : OAI221_X1 port map( B1 => n2170, B2 => n529, C1 => n1948, C2 => n2159
                           , A => n530, ZN => n1692);
   U334 : AOI222_X1 port map( A1 => n63, A2 => n2153, B1 => n191, B2 => n2148, 
                           C1 => n2147, C2 => n531, ZN => n530);
   U335 : OAI221_X1 port map( B1 => n2170, B2 => n532, C1 => n1947, C2 => n2159
                           , A => n533, ZN => n1691);
   U336 : AOI222_X1 port map( A1 => n62, A2 => n2153, B1 => n190, B2 => n2148, 
                           C1 => n2146, C2 => n534, ZN => n533);
   U337 : OAI221_X1 port map( B1 => n2170, B2 => n535, C1 => n1946, C2 => n2159
                           , A => n536, ZN => n1690);
   U338 : AOI222_X1 port map( A1 => n61, A2 => n2153, B1 => n189, B2 => n2148, 
                           C1 => n2146, C2 => n537, ZN => n536);
   U339 : OAI221_X1 port map( B1 => n2167, B2 => n619, C1 => n1921, C2 => n2161
                           , A => n620, ZN => n1665);
   U340 : AOI222_X1 port map( A1 => n36, A2 => n2155, B1 => n2150, B2 => n621, 
                           C1 => n2144, C2 => n622, ZN => n620);
   U341 : OAI221_X1 port map( B1 => n2167, B2 => n623, C1 => n1920, C2 => n2161
                           , A => n624, ZN => n1664);
   U342 : AOI222_X1 port map( A1 => n35, A2 => n2155, B1 => n2150, B2 => n625, 
                           C1 => n99, C2 => n2144, ZN => n624);
   U343 : OAI221_X1 port map( B1 => n2167, B2 => n626, C1 => n1919, C2 => n2161
                           , A => n627, ZN => n1663);
   U344 : AOI222_X1 port map( A1 => n34, A2 => n2155, B1 => n2150, B2 => n628, 
                           C1 => n98, C2 => n2144, ZN => n627);
   U345 : OAI221_X1 port map( B1 => n2167, B2 => n629, C1 => n1918, C2 => n2161
                           , A => n630, ZN => n1662);
   U346 : AOI222_X1 port map( A1 => n33, A2 => n2155, B1 => n2150, B2 => n631, 
                           C1 => n97, C2 => n2144, ZN => n630);
   U347 : OAI221_X1 port map( B1 => n2167, B2 => n632, C1 => n1917, C2 => n2161
                           , A => n633, ZN => n1661);
   U348 : AOI222_X1 port map( A1 => n32, A2 => n2155, B1 => n2150, B2 => n634, 
                           C1 => n96, C2 => n2144, ZN => n633);
   U349 : OAI221_X1 port map( B1 => n2167, B2 => n635, C1 => n1916, C2 => n2161
                           , A => n636, ZN => n1660);
   U350 : AOI222_X1 port map( A1 => n31, A2 => n2155, B1 => n2150, B2 => n637, 
                           C1 => n95, C2 => n2144, ZN => n636);
   U351 : OAI221_X1 port map( B1 => n2167, B2 => n638, C1 => n1915, C2 => n2161
                           , A => n639, ZN => n1659);
   U352 : AOI222_X1 port map( A1 => n30, A2 => n2155, B1 => n2150, B2 => n640, 
                           C1 => n94, C2 => n2144, ZN => n639);
   U353 : OAI221_X1 port map( B1 => n2167, B2 => n641, C1 => n1914, C2 => n2161
                           , A => n642, ZN => n1658);
   U354 : AOI222_X1 port map( A1 => n29, A2 => n2155, B1 => n2150, B2 => n643, 
                           C1 => n93, C2 => n2144, ZN => n642);
   U355 : OAI221_X1 port map( B1 => n2167, B2 => n644, C1 => n1913, C2 => n2162
                           , A => n645, ZN => n1657);
   U356 : AOI222_X1 port map( A1 => n28, A2 => n2156, B1 => n2150, B2 => n646, 
                           C1 => n92, C2 => n2144, ZN => n645);
   U357 : OAI221_X1 port map( B1 => n2167, B2 => n647, C1 => n1912, C2 => n2162
                           , A => n648, ZN => n1656);
   U358 : AOI222_X1 port map( A1 => n27, A2 => n2156, B1 => n2151, B2 => n649, 
                           C1 => n91, C2 => n2144, ZN => n648);
   U359 : OAI221_X1 port map( B1 => n2167, B2 => n650, C1 => n1911, C2 => n2162
                           , A => n651, ZN => n1655);
   U360 : AOI222_X1 port map( A1 => n26, A2 => n2156, B1 => n2151, B2 => n652, 
                           C1 => n90, C2 => n2144, ZN => n651);
   U361 : OAI221_X1 port map( B1 => n2167, B2 => n653, C1 => n1910, C2 => n2162
                           , A => n654, ZN => n1654);
   U362 : AOI222_X1 port map( A1 => n25, A2 => n2156, B1 => n2151, B2 => n655, 
                           C1 => n89, C2 => n2144, ZN => n654);
   U363 : OAI221_X1 port map( B1 => n2165, B2 => n716, C1 => n1890, C2 => n2164
                           , A => n717, ZN => n1634);
   U364 : AOI222_X1 port map( A1 => n5, A2 => n2157, B1 => n2152, B2 => n718, 
                           C1 => n69, C2 => n2142, ZN => n717);
   U365 : OAI221_X1 port map( B1 => n2165, B2 => n722, C1 => n1888, C2 => n2164
                           , A => n723, ZN => n1632);
   U366 : AOI222_X1 port map( A1 => n3, A2 => n2157, B1 => n2152, B2 => n724, 
                           C1 => n67, C2 => n2142, ZN => n723);
   U367 : OAI221_X1 port map( B1 => n2165, B2 => n725, C1 => n1887, C2 => n2164
                           , A => n726, ZN => n1631);
   U368 : AOI222_X1 port map( A1 => n2, A2 => n2157, B1 => n2152, B2 => n727, 
                           C1 => n66, C2 => n2142, ZN => n726);
   U369 : OAI221_X1 port map( B1 => n522, B2 => n2141, C1 => n1885, C2 => n2130
                           , A => n737, ZN => n1629);
   U370 : AOI222_X1 port map( A1 => n2129, A2 => n64, B1 => n2123, B2 => n192, 
                           C1 => n2117, C2 => n528, ZN => n737);
   U371 : OAI221_X1 port map( B1 => n529, B2 => n2141, C1 => n1884, C2 => n2130
                           , A => n744, ZN => n1627);
   U372 : AOI222_X1 port map( A1 => n2129, A2 => n63, B1 => n2123, B2 => n191, 
                           C1 => n2117, C2 => n531, ZN => n744);
   U373 : OAI221_X1 port map( B1 => n532, B2 => n2141, C1 => n1883, C2 => n2130
                           , A => n746, ZN => n1625);
   U374 : AOI222_X1 port map( A1 => n2129, A2 => n62, B1 => n2123, B2 => n190, 
                           C1 => n2117, C2 => n534, ZN => n746);
   U375 : OAI221_X1 port map( B1 => n535, B2 => n2141, C1 => n1882, C2 => n2130
                           , A => n748, ZN => n1623);
   U376 : AOI222_X1 port map( A1 => n2129, A2 => n61, B1 => n2123, B2 => n189, 
                           C1 => n2117, C2 => n537, ZN => n748);
   U377 : OAI221_X1 port map( B1 => n583, B2 => n2139, C1 => n1866, C2 => n2131
                           , A => n780, ZN => n1591);
   U378 : AOI222_X1 port map( A1 => n2127, A2 => n45, B1 => n2121, B2 => n585, 
                           C1 => n2115, C2 => n586, ZN => n780);
   U379 : OAI221_X1 port map( B1 => n587, B2 => n2139, C1 => n1865, C2 => n2131
                           , A => n782, ZN => n1589);
   U380 : AOI222_X1 port map( A1 => n2127, A2 => n44, B1 => n2121, B2 => n589, 
                           C1 => n2115, C2 => n590, ZN => n782);
   U381 : OAI221_X1 port map( B1 => n591, B2 => n2139, C1 => n1864, C2 => n2131
                           , A => n784, ZN => n1587);
   U382 : AOI222_X1 port map( A1 => n2127, A2 => n43, B1 => n2121, B2 => n593, 
                           C1 => n2115, C2 => n594, ZN => n784);
   U383 : OAI221_X1 port map( B1 => n595, B2 => n2139, C1 => n1863, C2 => n2131
                           , A => n786, ZN => n1585);
   U384 : AOI222_X1 port map( A1 => n2127, A2 => n42, B1 => n2121, B2 => n597, 
                           C1 => n2115, C2 => n598, ZN => n786);
   U385 : OAI221_X1 port map( B1 => n599, B2 => n2139, C1 => n1862, C2 => n2131
                           , A => n788, ZN => n1583);
   U386 : AOI222_X1 port map( A1 => n2127, A2 => n41, B1 => n2121, B2 => n601, 
                           C1 => n2115, C2 => n602, ZN => n788);
   U387 : OAI221_X1 port map( B1 => n603, B2 => n2139, C1 => n1861, C2 => n2131
                           , A => n790, ZN => n1581);
   U388 : AOI222_X1 port map( A1 => n2127, A2 => n40, B1 => n2121, B2 => n605, 
                           C1 => n2115, C2 => n606, ZN => n790);
   U389 : OAI221_X1 port map( B1 => n607, B2 => n2139, C1 => n1860, C2 => n2132
                           , A => n792, ZN => n1579);
   U390 : AOI222_X1 port map( A1 => n2127, A2 => n39, B1 => n2121, B2 => n609, 
                           C1 => n2115, C2 => n610, ZN => n792);
   U391 : OAI221_X1 port map( B1 => n611, B2 => n2139, C1 => n1859, C2 => n2132
                           , A => n794, ZN => n1577);
   U392 : AOI222_X1 port map( A1 => n2127, A2 => n38, B1 => n2121, B2 => n613, 
                           C1 => n2115, C2 => n614, ZN => n794);
   U393 : OAI221_X1 port map( B1 => n615, B2 => n2139, C1 => n1858, C2 => n2132
                           , A => n796, ZN => n1575);
   U394 : AOI222_X1 port map( A1 => n2127, A2 => n37, B1 => n2121, B2 => n617, 
                           C1 => n2115, C2 => n618, ZN => n796);
   U395 : OAI221_X1 port map( B1 => n619, B2 => n2138, C1 => n1857, C2 => n2132
                           , A => n798, ZN => n1573);
   U396 : AOI222_X1 port map( A1 => n2126, A2 => n36, B1 => n2120, B2 => n621, 
                           C1 => n2114, C2 => n622, ZN => n798);
   U397 : OAI221_X1 port map( B1 => n2169, B2 => n538, C1 => n1945, C2 => n2159
                           , A => n539, ZN => n1689);
   U398 : AOI222_X1 port map( A1 => n60, A2 => n2153, B1 => n188, B2 => n2148, 
                           C1 => n2146, C2 => n540, ZN => n539);
   U399 : OAI221_X1 port map( B1 => n2169, B2 => n541, C1 => n1944, C2 => n2159
                           , A => n542, ZN => n1688);
   U400 : AOI222_X1 port map( A1 => n59, A2 => n2153, B1 => n187, B2 => n2148, 
                           C1 => n2146, C2 => n543, ZN => n542);
   U401 : OAI221_X1 port map( B1 => n2169, B2 => n544, C1 => n1943, C2 => n2159
                           , A => n545, ZN => n1687);
   U402 : AOI222_X1 port map( A1 => n58, A2 => n2153, B1 => n186, B2 => n2148, 
                           C1 => n2146, C2 => n546, ZN => n545);
   U403 : OAI221_X1 port map( B1 => n2169, B2 => n547, C1 => n1942, C2 => n2159
                           , A => n548, ZN => n1686);
   U404 : AOI222_X1 port map( A1 => n57, A2 => n2153, B1 => n185, B2 => n2148, 
                           C1 => n2146, C2 => n549, ZN => n548);
   U405 : OAI221_X1 port map( B1 => n2169, B2 => n550, C1 => n1941, C2 => n2159
                           , A => n551, ZN => n1685);
   U406 : AOI222_X1 port map( A1 => n56, A2 => n2153, B1 => n184, B2 => n2148, 
                           C1 => n2146, C2 => n552, ZN => n551);
   U407 : OAI221_X1 port map( B1 => n2169, B2 => n553, C1 => n1940, C2 => n2159
                           , A => n554, ZN => n1684);
   U408 : AOI222_X1 port map( A1 => n55, A2 => n2153, B1 => n183, B2 => n2148, 
                           C1 => n2146, C2 => n555, ZN => n554);
   U409 : OAI221_X1 port map( B1 => n2169, B2 => n556, C1 => n1939, C2 => n2159
                           , A => n557, ZN => n1683);
   U410 : AOI222_X1 port map( A1 => n54, A2 => n2153, B1 => n182, B2 => n2148, 
                           C1 => n2146, C2 => n558, ZN => n557);
   U411 : OAI221_X1 port map( B1 => n2169, B2 => n559, C1 => n1938, C2 => n2159
                           , A => n560, ZN => n1682);
   U412 : AOI222_X1 port map( A1 => n53, A2 => n2153, B1 => n181, B2 => n2148, 
                           C1 => n2146, C2 => n561, ZN => n560);
   U413 : OAI221_X1 port map( B1 => n2168, B2 => n583, C1 => n1930, C2 => n2160
                           , A => n584, ZN => n1674);
   U414 : AOI222_X1 port map( A1 => n45, A2 => n2154, B1 => n2149, B2 => n585, 
                           C1 => n2145, C2 => n586, ZN => n584);
   U415 : OAI221_X1 port map( B1 => n2168, B2 => n587, C1 => n1929, C2 => n2160
                           , A => n588, ZN => n1673);
   U416 : AOI222_X1 port map( A1 => n44, A2 => n2154, B1 => n2149, B2 => n589, 
                           C1 => n2145, C2 => n590, ZN => n588);
   U417 : OAI221_X1 port map( B1 => n2168, B2 => n591, C1 => n1928, C2 => n2160
                           , A => n592, ZN => n1672);
   U418 : AOI222_X1 port map( A1 => n43, A2 => n2154, B1 => n2149, B2 => n593, 
                           C1 => n2145, C2 => n594, ZN => n592);
   U419 : OAI221_X1 port map( B1 => n2168, B2 => n595, C1 => n1927, C2 => n2160
                           , A => n596, ZN => n1671);
   U420 : AOI222_X1 port map( A1 => n42, A2 => n2154, B1 => n2149, B2 => n597, 
                           C1 => n2145, C2 => n598, ZN => n596);
   U421 : OAI221_X1 port map( B1 => n2168, B2 => n599, C1 => n1926, C2 => n2160
                           , A => n600, ZN => n1670);
   U422 : AOI222_X1 port map( A1 => n41, A2 => n2154, B1 => n2149, B2 => n601, 
                           C1 => n2145, C2 => n602, ZN => n600);
   U423 : OAI221_X1 port map( B1 => n2168, B2 => n603, C1 => n1925, C2 => n2160
                           , A => n604, ZN => n1669);
   U424 : AOI222_X1 port map( A1 => n40, A2 => n2154, B1 => n2150, B2 => n605, 
                           C1 => n2145, C2 => n606, ZN => n604);
   U425 : OAI221_X1 port map( B1 => n2168, B2 => n607, C1 => n1924, C2 => n2161
                           , A => n608, ZN => n1668);
   U426 : AOI222_X1 port map( A1 => n39, A2 => n2155, B1 => n2150, B2 => n609, 
                           C1 => n2145, C2 => n610, ZN => n608);
   U427 : OAI221_X1 port map( B1 => n2168, B2 => n611, C1 => n1923, C2 => n2161
                           , A => n612, ZN => n1667);
   U428 : AOI222_X1 port map( A1 => n38, A2 => n2155, B1 => n2150, B2 => n613, 
                           C1 => n2145, C2 => n614, ZN => n612);
   U429 : OAI221_X1 port map( B1 => n2168, B2 => n615, C1 => n1922, C2 => n2161
                           , A => n616, ZN => n1666);
   U430 : AOI222_X1 port map( A1 => n37, A2 => n2155, B1 => n2150, B2 => n617, 
                           C1 => n2145, C2 => n618, ZN => n616);
   U431 : OAI22_X1 port map( A1 => n1950, A2 => n2099, B1 => n743, B2 => n2093,
                           ZN => n1501);
   U432 : OAI22_X1 port map( A1 => n1951, A2 => n2099, B1 => n745, B2 => n2093,
                           ZN => n1500);
   U433 : OAI22_X1 port map( A1 => n1952, A2 => n2099, B1 => n747, B2 => n2093,
                           ZN => n1499);
   U434 : OAI22_X1 port map( A1 => n1953, A2 => n2099, B1 => n749, B2 => n2093,
                           ZN => n1498);
   U435 : OAI22_X1 port map( A1 => n1821, A2 => n2087, B1 => n743, B2 => n2081,
                           ZN => n1437);
   U436 : OAI22_X1 port map( A1 => n1820, A2 => n2087, B1 => n745, B2 => n2081,
                           ZN => n1436);
   U437 : OAI22_X1 port map( A1 => n1819, A2 => n2087, B1 => n747, B2 => n2081,
                           ZN => n1435);
   U438 : OAI22_X1 port map( A1 => n1818, A2 => n2087, B1 => n749, B2 => n2081,
                           ZN => n1434);
   U439 : OAI22_X1 port map( A1 => n2010, A2 => n2075, B1 => n743, B2 => n2069,
                           ZN => n1373);
   U440 : OAI22_X1 port map( A1 => n2011, A2 => n2075, B1 => n745, B2 => n2069,
                           ZN => n1372);
   U441 : OAI22_X1 port map( A1 => n2012, A2 => n2075, B1 => n747, B2 => n2069,
                           ZN => n1371);
   U442 : OAI22_X1 port map( A1 => n2013, A2 => n2075, B1 => n749, B2 => n2069,
                           ZN => n1370);
   U443 : OAI22_X1 port map( A1 => n1954, A2 => n2099, B1 => n751, B2 => n2092,
                           ZN => n1497);
   U444 : OAI22_X1 port map( A1 => n1955, A2 => n2098, B1 => n753, B2 => n2092,
                           ZN => n1496);
   U445 : OAI22_X1 port map( A1 => n1956, A2 => n2098, B1 => n755, B2 => n2092,
                           ZN => n1495);
   U446 : OAI22_X1 port map( A1 => n1957, A2 => n2098, B1 => n757, B2 => n2092,
                           ZN => n1494);
   U447 : OAI22_X1 port map( A1 => n1958, A2 => n2098, B1 => n759, B2 => n2092,
                           ZN => n1493);
   U448 : OAI22_X1 port map( A1 => n1959, A2 => n2098, B1 => n761, B2 => n2092,
                           ZN => n1492);
   U449 : OAI22_X1 port map( A1 => n1960, A2 => n2098, B1 => n763, B2 => n2092,
                           ZN => n1491);
   U450 : OAI22_X1 port map( A1 => n1961, A2 => n2098, B1 => n765, B2 => n2092,
                           ZN => n1490);
   U451 : OAI22_X1 port map( A1 => n1962, A2 => n2098, B1 => n767, B2 => n2092,
                           ZN => n1489);
   U452 : OAI22_X1 port map( A1 => n1963, A2 => n2098, B1 => n769, B2 => n2092,
                           ZN => n1488);
   U453 : OAI22_X1 port map( A1 => n1964, A2 => n2098, B1 => n771, B2 => n2092,
                           ZN => n1487);
   U454 : OAI22_X1 port map( A1 => n1965, A2 => n2098, B1 => n773, B2 => n2092,
                           ZN => n1486);
   U455 : OAI22_X1 port map( A1 => n1966, A2 => n2098, B1 => n775, B2 => n2091,
                           ZN => n1485);
   U456 : OAI22_X1 port map( A1 => n1967, A2 => n2097, B1 => n777, B2 => n2091,
                           ZN => n1484);
   U457 : OAI22_X1 port map( A1 => n1968, A2 => n2097, B1 => n779, B2 => n2091,
                           ZN => n1483);
   U458 : OAI22_X1 port map( A1 => n1969, A2 => n2097, B1 => n781, B2 => n2091,
                           ZN => n1482);
   U459 : OAI22_X1 port map( A1 => n1970, A2 => n2097, B1 => n783, B2 => n2091,
                           ZN => n1481);
   U460 : OAI22_X1 port map( A1 => n1971, A2 => n2097, B1 => n785, B2 => n2091,
                           ZN => n1480);
   U461 : OAI22_X1 port map( A1 => n1972, A2 => n2097, B1 => n787, B2 => n2091,
                           ZN => n1479);
   U462 : OAI22_X1 port map( A1 => n1973, A2 => n2097, B1 => n789, B2 => n2091,
                           ZN => n1478);
   U463 : OAI22_X1 port map( A1 => n1974, A2 => n2097, B1 => n791, B2 => n2091,
                           ZN => n1477);
   U464 : OAI22_X1 port map( A1 => n1975, A2 => n2097, B1 => n793, B2 => n2091,
                           ZN => n1476);
   U465 : OAI22_X1 port map( A1 => n1976, A2 => n2097, B1 => n795, B2 => n2091,
                           ZN => n1475);
   U466 : OAI22_X1 port map( A1 => n1977, A2 => n2097, B1 => n797, B2 => n2091,
                           ZN => n1474);
   U467 : OAI22_X1 port map( A1 => n1978, A2 => n2097, B1 => n799, B2 => n2090,
                           ZN => n1473);
   U468 : OAI22_X1 port map( A1 => n1979, A2 => n2096, B1 => n801, B2 => n2090,
                           ZN => n1472);
   U469 : OAI22_X1 port map( A1 => n1980, A2 => n2096, B1 => n803, B2 => n2090,
                           ZN => n1471);
   U470 : OAI22_X1 port map( A1 => n1981, A2 => n2096, B1 => n805, B2 => n2090,
                           ZN => n1470);
   U471 : OAI22_X1 port map( A1 => n1982, A2 => n2096, B1 => n807, B2 => n2090,
                           ZN => n1469);
   U472 : OAI22_X1 port map( A1 => n1983, A2 => n2096, B1 => n809, B2 => n2090,
                           ZN => n1468);
   U473 : OAI22_X1 port map( A1 => n1984, A2 => n2096, B1 => n811, B2 => n2090,
                           ZN => n1467);
   U474 : OAI22_X1 port map( A1 => n1985, A2 => n2096, B1 => n813, B2 => n2090,
                           ZN => n1466);
   U475 : OAI22_X1 port map( A1 => n1986, A2 => n2096, B1 => n815, B2 => n2090,
                           ZN => n1465);
   U476 : OAI22_X1 port map( A1 => n1987, A2 => n2096, B1 => n817, B2 => n2090,
                           ZN => n1464);
   U477 : OAI22_X1 port map( A1 => n1988, A2 => n2096, B1 => n819, B2 => n2090,
                           ZN => n1463);
   U478 : OAI22_X1 port map( A1 => n1989, A2 => n2096, B1 => n821, B2 => n2090,
                           ZN => n1462);
   U479 : OAI22_X1 port map( A1 => n1990, A2 => n2096, B1 => n823, B2 => n2089,
                           ZN => n1461);
   U480 : OAI22_X1 port map( A1 => n1991, A2 => n2095, B1 => n825, B2 => n2089,
                           ZN => n1460);
   U481 : OAI22_X1 port map( A1 => n1992, A2 => n2095, B1 => n827, B2 => n2089,
                           ZN => n1459);
   U482 : OAI22_X1 port map( A1 => n1993, A2 => n2095, B1 => n829, B2 => n2089,
                           ZN => n1458);
   U483 : OAI22_X1 port map( A1 => n1994, A2 => n2095, B1 => n831, B2 => n2089,
                           ZN => n1457);
   U484 : OAI22_X1 port map( A1 => n1995, A2 => n2095, B1 => n833, B2 => n2089,
                           ZN => n1456);
   U485 : OAI22_X1 port map( A1 => n1996, A2 => n2095, B1 => n835, B2 => n2089,
                           ZN => n1455);
   U486 : OAI22_X1 port map( A1 => n1997, A2 => n2095, B1 => n837, B2 => n2089,
                           ZN => n1454);
   U487 : OAI22_X1 port map( A1 => n1998, A2 => n2095, B1 => n839, B2 => n2089,
                           ZN => n1453);
   U488 : OAI22_X1 port map( A1 => n1999, A2 => n2095, B1 => n841, B2 => n2089,
                           ZN => n1452);
   U489 : OAI22_X1 port map( A1 => n2000, A2 => n2095, B1 => n843, B2 => n2089,
                           ZN => n1451);
   U490 : OAI22_X1 port map( A1 => n2001, A2 => n2095, B1 => n845, B2 => n2089,
                           ZN => n1450);
   U491 : OAI22_X1 port map( A1 => n1204, A2 => n2095, B1 => n847, B2 => n2088,
                           ZN => n1449);
   U492 : OAI22_X1 port map( A1 => n1202, A2 => n2094, B1 => n849, B2 => n2088,
                           ZN => n1448);
   U493 : OAI22_X1 port map( A1 => n1200, A2 => n2094, B1 => n851, B2 => n2088,
                           ZN => n1447);
   U494 : OAI22_X1 port map( A1 => n2002, A2 => n2094, B1 => n853, B2 => n2088,
                           ZN => n1446);
   U495 : OAI22_X1 port map( A1 => n2003, A2 => n2094, B1 => n855, B2 => n2088,
                           ZN => n1445);
   U496 : OAI22_X1 port map( A1 => n2004, A2 => n2094, B1 => n857, B2 => n2088,
                           ZN => n1444);
   U497 : OAI22_X1 port map( A1 => n2005, A2 => n2094, B1 => n859, B2 => n2088,
                           ZN => n1443);
   U498 : OAI22_X1 port map( A1 => n2006, A2 => n2094, B1 => n861, B2 => n2088,
                           ZN => n1442);
   U499 : OAI22_X1 port map( A1 => n2007, A2 => n2094, B1 => n863, B2 => n2088,
                           ZN => n1441);
   U500 : OAI22_X1 port map( A1 => n2008, A2 => n2094, B1 => n865, B2 => n2088,
                           ZN => n1440);
   U501 : OAI22_X1 port map( A1 => n2009, A2 => n2094, B1 => n867, B2 => n2088,
                           ZN => n1439);
   U502 : OAI22_X1 port map( A1 => n415, A2 => n2094, B1 => n871, B2 => n2088, 
                           ZN => n1438);
   U503 : OAI22_X1 port map( A1 => n1817, A2 => n2087, B1 => n751, B2 => n2080,
                           ZN => n1433);
   U504 : OAI22_X1 port map( A1 => n1816, A2 => n2086, B1 => n753, B2 => n2080,
                           ZN => n1432);
   U505 : OAI22_X1 port map( A1 => n1815, A2 => n2086, B1 => n755, B2 => n2080,
                           ZN => n1431);
   U506 : OAI22_X1 port map( A1 => n1814, A2 => n2086, B1 => n757, B2 => n2080,
                           ZN => n1430);
   U507 : OAI22_X1 port map( A1 => n1813, A2 => n2086, B1 => n759, B2 => n2080,
                           ZN => n1429);
   U508 : OAI22_X1 port map( A1 => n1812, A2 => n2086, B1 => n761, B2 => n2080,
                           ZN => n1428);
   U509 : OAI22_X1 port map( A1 => n1811, A2 => n2086, B1 => n763, B2 => n2080,
                           ZN => n1427);
   U510 : OAI22_X1 port map( A1 => n1810, A2 => n2086, B1 => n765, B2 => n2080,
                           ZN => n1426);
   U511 : OAI22_X1 port map( A1 => n1809, A2 => n2086, B1 => n767, B2 => n2080,
                           ZN => n1425);
   U512 : OAI22_X1 port map( A1 => n1808, A2 => n2086, B1 => n769, B2 => n2080,
                           ZN => n1424);
   U513 : OAI22_X1 port map( A1 => n1807, A2 => n2086, B1 => n771, B2 => n2080,
                           ZN => n1423);
   U514 : OAI22_X1 port map( A1 => n1806, A2 => n2086, B1 => n773, B2 => n2080,
                           ZN => n1422);
   U515 : OAI22_X1 port map( A1 => n1805, A2 => n2086, B1 => n775, B2 => n2079,
                           ZN => n1421);
   U516 : OAI22_X1 port map( A1 => n1804, A2 => n2085, B1 => n777, B2 => n2079,
                           ZN => n1420);
   U517 : OAI22_X1 port map( A1 => n1803, A2 => n2085, B1 => n779, B2 => n2079,
                           ZN => n1419);
   U518 : OAI22_X1 port map( A1 => n1802, A2 => n2085, B1 => n781, B2 => n2079,
                           ZN => n1418);
   U519 : OAI22_X1 port map( A1 => n1801, A2 => n2085, B1 => n783, B2 => n2079,
                           ZN => n1417);
   U520 : OAI22_X1 port map( A1 => n1800, A2 => n2085, B1 => n785, B2 => n2079,
                           ZN => n1416);
   U521 : OAI22_X1 port map( A1 => n1799, A2 => n2085, B1 => n787, B2 => n2079,
                           ZN => n1415);
   U522 : OAI22_X1 port map( A1 => n1798, A2 => n2085, B1 => n789, B2 => n2079,
                           ZN => n1414);
   U523 : OAI22_X1 port map( A1 => n1797, A2 => n2085, B1 => n791, B2 => n2079,
                           ZN => n1413);
   U524 : OAI22_X1 port map( A1 => n1796, A2 => n2085, B1 => n793, B2 => n2079,
                           ZN => n1412);
   U525 : OAI22_X1 port map( A1 => n1795, A2 => n2085, B1 => n795, B2 => n2079,
                           ZN => n1411);
   U526 : OAI22_X1 port map( A1 => n1794, A2 => n2085, B1 => n797, B2 => n2079,
                           ZN => n1410);
   U527 : OAI22_X1 port map( A1 => n1793, A2 => n2085, B1 => n799, B2 => n2078,
                           ZN => n1409);
   U528 : OAI22_X1 port map( A1 => n2029, A2 => n2084, B1 => n801, B2 => n2078,
                           ZN => n1408);
   U529 : OAI22_X1 port map( A1 => n2030, A2 => n2084, B1 => n803, B2 => n2078,
                           ZN => n1407);
   U530 : OAI22_X1 port map( A1 => n2031, A2 => n2084, B1 => n805, B2 => n2078,
                           ZN => n1406);
   U531 : OAI22_X1 port map( A1 => n2032, A2 => n2084, B1 => n807, B2 => n2078,
                           ZN => n1405);
   U532 : OAI22_X1 port map( A1 => n2033, A2 => n2084, B1 => n809, B2 => n2078,
                           ZN => n1404);
   U533 : OAI22_X1 port map( A1 => n2034, A2 => n2084, B1 => n811, B2 => n2078,
                           ZN => n1403);
   U534 : OAI22_X1 port map( A1 => n2035, A2 => n2084, B1 => n813, B2 => n2078,
                           ZN => n1402);
   U535 : OAI22_X1 port map( A1 => n2036, A2 => n2084, B1 => n815, B2 => n2078,
                           ZN => n1401);
   U536 : OAI22_X1 port map( A1 => n2037, A2 => n2084, B1 => n817, B2 => n2078,
                           ZN => n1400);
   U537 : OAI22_X1 port map( A1 => n2038, A2 => n2084, B1 => n819, B2 => n2078,
                           ZN => n1399);
   U538 : OAI22_X1 port map( A1 => n2039, A2 => n2084, B1 => n821, B2 => n2078,
                           ZN => n1398);
   U539 : OAI22_X1 port map( A1 => n2040, A2 => n2084, B1 => n823, B2 => n2077,
                           ZN => n1397);
   U540 : OAI22_X1 port map( A1 => n2041, A2 => n2083, B1 => n825, B2 => n2077,
                           ZN => n1396);
   U541 : OAI22_X1 port map( A1 => n2042, A2 => n2083, B1 => n827, B2 => n2077,
                           ZN => n1395);
   U542 : OAI22_X1 port map( A1 => n2043, A2 => n2083, B1 => n829, B2 => n2077,
                           ZN => n1394);
   U543 : OAI22_X1 port map( A1 => n2044, A2 => n2083, B1 => n831, B2 => n2077,
                           ZN => n1393);
   U544 : OAI22_X1 port map( A1 => n2045, A2 => n2083, B1 => n833, B2 => n2077,
                           ZN => n1392);
   U545 : OAI22_X1 port map( A1 => n2046, A2 => n2083, B1 => n835, B2 => n2077,
                           ZN => n1391);
   U546 : OAI22_X1 port map( A1 => n2047, A2 => n2083, B1 => n837, B2 => n2077,
                           ZN => n1390);
   U547 : OAI22_X1 port map( A1 => n2048, A2 => n2083, B1 => n839, B2 => n2077,
                           ZN => n1389);
   U548 : OAI22_X1 port map( A1 => n2049, A2 => n2083, B1 => n841, B2 => n2077,
                           ZN => n1388);
   U549 : OAI22_X1 port map( A1 => n2050, A2 => n2083, B1 => n843, B2 => n2077,
                           ZN => n1387);
   U550 : OAI22_X1 port map( A1 => n2051, A2 => n2083, B1 => n845, B2 => n2077,
                           ZN => n1386);
   U551 : OAI22_X1 port map( A1 => n2052, A2 => n2083, B1 => n847, B2 => n2076,
                           ZN => n1385);
   U552 : OAI22_X1 port map( A1 => n2053, A2 => n2082, B1 => n849, B2 => n2076,
                           ZN => n1384);
   U553 : OAI22_X1 port map( A1 => n2054, A2 => n2082, B1 => n851, B2 => n2076,
                           ZN => n1383);
   U554 : OAI22_X1 port map( A1 => n2055, A2 => n2082, B1 => n853, B2 => n2076,
                           ZN => n1382);
   U555 : OAI22_X1 port map( A1 => n2056, A2 => n2082, B1 => n855, B2 => n2076,
                           ZN => n1381);
   U556 : OAI22_X1 port map( A1 => n2057, A2 => n2082, B1 => n857, B2 => n2076,
                           ZN => n1380);
   U557 : OAI22_X1 port map( A1 => n2058, A2 => n2082, B1 => n859, B2 => n2076,
                           ZN => n1379);
   U558 : OAI22_X1 port map( A1 => n2059, A2 => n2082, B1 => n861, B2 => n2076,
                           ZN => n1378);
   U559 : OAI22_X1 port map( A1 => n2060, A2 => n2082, B1 => n863, B2 => n2076,
                           ZN => n1377);
   U560 : OAI22_X1 port map( A1 => n2061, A2 => n2082, B1 => n865, B2 => n2076,
                           ZN => n1376);
   U561 : OAI22_X1 port map( A1 => n2062, A2 => n2082, B1 => n867, B2 => n2076,
                           ZN => n1375);
   U562 : OAI22_X1 port map( A1 => n2063, A2 => n2082, B1 => n871, B2 => n2076,
                           ZN => n1374);
   U563 : OAI22_X1 port map( A1 => n2014, A2 => n2075, B1 => n751, B2 => n2068,
                           ZN => n1369);
   U564 : OAI22_X1 port map( A1 => n2015, A2 => n2074, B1 => n753, B2 => n2068,
                           ZN => n1368);
   U565 : OAI22_X1 port map( A1 => n2016, A2 => n2074, B1 => n755, B2 => n2068,
                           ZN => n1367);
   U566 : OAI22_X1 port map( A1 => n2017, A2 => n2074, B1 => n757, B2 => n2068,
                           ZN => n1366);
   U567 : OAI22_X1 port map( A1 => n2018, A2 => n2074, B1 => n759, B2 => n2068,
                           ZN => n1365);
   U568 : OAI22_X1 port map( A1 => n2019, A2 => n2074, B1 => n761, B2 => n2068,
                           ZN => n1364);
   U569 : OAI22_X1 port map( A1 => n2020, A2 => n2074, B1 => n763, B2 => n2068,
                           ZN => n1363);
   U570 : OAI22_X1 port map( A1 => n2021, A2 => n2074, B1 => n765, B2 => n2068,
                           ZN => n1362);
   U571 : OAI22_X1 port map( A1 => n2022, A2 => n2074, B1 => n767, B2 => n2068,
                           ZN => n1361);
   U572 : OAI22_X1 port map( A1 => n2023, A2 => n2074, B1 => n769, B2 => n2068,
                           ZN => n1360);
   U573 : OAI22_X1 port map( A1 => n2024, A2 => n2074, B1 => n771, B2 => n2068,
                           ZN => n1359);
   U574 : OAI22_X1 port map( A1 => n2025, A2 => n2074, B1 => n773, B2 => n2068,
                           ZN => n1358);
   U575 : OAI22_X1 port map( A1 => n2026, A2 => n2074, B1 => n775, B2 => n2067,
                           ZN => n1357);
   U576 : OAI22_X1 port map( A1 => n2027, A2 => n2073, B1 => n777, B2 => n2067,
                           ZN => n1356);
   U577 : OAI22_X1 port map( A1 => n2028, A2 => n2073, B1 => n779, B2 => n2067,
                           ZN => n1355);
   U578 : OAI22_X1 port map( A1 => n1738, A2 => n2073, B1 => n781, B2 => n2067,
                           ZN => n1354);
   U579 : OAI22_X1 port map( A1 => n1737, A2 => n2073, B1 => n783, B2 => n2067,
                           ZN => n1353);
   U580 : OAI22_X1 port map( A1 => n1736, A2 => n2073, B1 => n785, B2 => n2067,
                           ZN => n1352);
   U581 : OAI22_X1 port map( A1 => n1735, A2 => n2073, B1 => n787, B2 => n2067,
                           ZN => n1351);
   U582 : OAI22_X1 port map( A1 => n1734, A2 => n2073, B1 => n789, B2 => n2067,
                           ZN => n1350);
   U583 : OAI22_X1 port map( A1 => n1733, A2 => n2073, B1 => n791, B2 => n2067,
                           ZN => n1349);
   U584 : OAI22_X1 port map( A1 => n1732, A2 => n2073, B1 => n793, B2 => n2067,
                           ZN => n1348);
   U585 : OAI22_X1 port map( A1 => n1731, A2 => n2073, B1 => n795, B2 => n2067,
                           ZN => n1347);
   U586 : OAI22_X1 port map( A1 => n1730, A2 => n2073, B1 => n797, B2 => n2067,
                           ZN => n1346);
   U587 : OAI22_X1 port map( A1 => n1729, A2 => n2073, B1 => n799, B2 => n2066,
                           ZN => n1345);
   U588 : OAI22_X1 port map( A1 => n1728, A2 => n2072, B1 => n801, B2 => n2066,
                           ZN => n1344);
   U589 : OAI22_X1 port map( A1 => n1727, A2 => n2072, B1 => n803, B2 => n2066,
                           ZN => n1343);
   U590 : OAI22_X1 port map( A1 => n1726, A2 => n2072, B1 => n805, B2 => n2066,
                           ZN => n1342);
   U591 : OAI22_X1 port map( A1 => n1725, A2 => n2072, B1 => n807, B2 => n2066,
                           ZN => n1341);
   U592 : OAI22_X1 port map( A1 => n1724, A2 => n2072, B1 => n809, B2 => n2066,
                           ZN => n1340);
   U593 : OAI22_X1 port map( A1 => n1723, A2 => n2072, B1 => n811, B2 => n2066,
                           ZN => n1339);
   U594 : OAI22_X1 port map( A1 => n1722, A2 => n2072, B1 => n813, B2 => n2066,
                           ZN => n1338);
   U595 : OAI22_X1 port map( A1 => n1721, A2 => n2072, B1 => n815, B2 => n2066,
                           ZN => n1337);
   U596 : OAI22_X1 port map( A1 => n1720, A2 => n2072, B1 => n817, B2 => n2066,
                           ZN => n1336);
   U597 : OAI22_X1 port map( A1 => n1719, A2 => n2072, B1 => n819, B2 => n2066,
                           ZN => n1335);
   U598 : OAI22_X1 port map( A1 => n1718, A2 => n2072, B1 => n821, B2 => n2066,
                           ZN => n1334);
   U599 : OAI22_X1 port map( A1 => n1717, A2 => n2072, B1 => n823, B2 => n2065,
                           ZN => n1333);
   U600 : OAI22_X1 port map( A1 => n1716, A2 => n2071, B1 => n825, B2 => n2065,
                           ZN => n1332);
   U601 : OAI22_X1 port map( A1 => n1715, A2 => n2071, B1 => n827, B2 => n2065,
                           ZN => n1331);
   U602 : OAI22_X1 port map( A1 => n1714, A2 => n2071, B1 => n829, B2 => n2065,
                           ZN => n1330);
   U603 : OAI22_X1 port map( A1 => n1713, A2 => n2071, B1 => n831, B2 => n2065,
                           ZN => n1329);
   U604 : OAI22_X1 port map( A1 => n1712, A2 => n2071, B1 => n833, B2 => n2065,
                           ZN => n1328);
   U605 : OAI22_X1 port map( A1 => n1711, A2 => n2071, B1 => n835, B2 => n2065,
                           ZN => n1327);
   U606 : OAI22_X1 port map( A1 => n1710, A2 => n2071, B1 => n837, B2 => n2065,
                           ZN => n1326);
   U607 : OAI22_X1 port map( A1 => n1709, A2 => n2071, B1 => n839, B2 => n2065,
                           ZN => n1325);
   U608 : OAI22_X1 port map( A1 => n1708, A2 => n2071, B1 => n841, B2 => n2065,
                           ZN => n1324);
   U609 : OAI22_X1 port map( A1 => n1707, A2 => n2071, B1 => n843, B2 => n2065,
                           ZN => n1323);
   U610 : OAI22_X1 port map( A1 => n1706, A2 => n2071, B1 => n845, B2 => n2065,
                           ZN => n1322);
   U611 : OAI22_X1 port map( A1 => n1705, A2 => n2071, B1 => n847, B2 => n2064,
                           ZN => n1321);
   U612 : OAI22_X1 port map( A1 => n1704, A2 => n2070, B1 => n849, B2 => n2064,
                           ZN => n1320);
   U613 : OAI22_X1 port map( A1 => n1703, A2 => n2070, B1 => n851, B2 => n2064,
                           ZN => n1319);
   U614 : OAI22_X1 port map( A1 => n1702, A2 => n2070, B1 => n853, B2 => n2064,
                           ZN => n1318);
   U615 : OAI22_X1 port map( A1 => n1701, A2 => n2070, B1 => n855, B2 => n2064,
                           ZN => n1317);
   U616 : OAI22_X1 port map( A1 => n1700, A2 => n2070, B1 => n857, B2 => n2064,
                           ZN => n1316);
   U617 : OAI22_X1 port map( A1 => n1699, A2 => n2070, B1 => n859, B2 => n2064,
                           ZN => n1315);
   U618 : OAI22_X1 port map( A1 => n1698, A2 => n2070, B1 => n861, B2 => n2064,
                           ZN => n1314);
   U619 : OAI22_X1 port map( A1 => n1697, A2 => n2070, B1 => n863, B2 => n2064,
                           ZN => n1313);
   U620 : OAI22_X1 port map( A1 => n1696, A2 => n2070, B1 => n865, B2 => n2064,
                           ZN => n1312);
   U621 : OAI22_X1 port map( A1 => n1695, A2 => n2070, B1 => n867, B2 => n2064,
                           ZN => n1311);
   U622 : OAI22_X1 port map( A1 => n1694, A2 => n2070, B1 => n871, B2 => n2064,
                           ZN => n1310);
   U623 : INV_X1 port map( A => DATAIN(0), ZN => n743);
   U624 : INV_X1 port map( A => DATAIN(1), ZN => n745);
   U625 : INV_X1 port map( A => DATAIN(2), ZN => n747);
   U626 : INV_X1 port map( A => DATAIN(3), ZN => n749);
   U627 : INV_X1 port map( A => DATAIN(4), ZN => n751);
   U628 : INV_X1 port map( A => DATAIN(5), ZN => n753);
   U629 : INV_X1 port map( A => DATAIN(6), ZN => n755);
   U630 : INV_X1 port map( A => DATAIN(7), ZN => n757);
   U631 : INV_X1 port map( A => DATAIN(8), ZN => n759);
   U632 : INV_X1 port map( A => DATAIN(9), ZN => n761);
   U633 : INV_X1 port map( A => DATAIN(10), ZN => n763);
   U634 : INV_X1 port map( A => DATAIN(11), ZN => n765);
   U635 : INV_X1 port map( A => DATAIN(12), ZN => n767);
   U636 : INV_X1 port map( A => DATAIN(13), ZN => n769);
   U637 : INV_X1 port map( A => DATAIN(14), ZN => n771);
   U638 : INV_X1 port map( A => DATAIN(15), ZN => n773);
   U639 : INV_X1 port map( A => DATAIN(16), ZN => n775);
   U640 : INV_X1 port map( A => DATAIN(17), ZN => n777);
   U641 : INV_X1 port map( A => DATAIN(18), ZN => n779);
   U642 : INV_X1 port map( A => DATAIN(19), ZN => n781);
   U643 : INV_X1 port map( A => DATAIN(20), ZN => n783);
   U644 : INV_X1 port map( A => DATAIN(21), ZN => n785);
   U645 : INV_X1 port map( A => DATAIN(22), ZN => n787);
   U646 : INV_X1 port map( A => DATAIN(23), ZN => n789);
   U647 : INV_X1 port map( A => DATAIN(24), ZN => n791);
   U648 : INV_X1 port map( A => DATAIN(25), ZN => n793);
   U649 : INV_X1 port map( A => DATAIN(26), ZN => n795);
   U650 : INV_X1 port map( A => DATAIN(27), ZN => n797);
   U651 : INV_X1 port map( A => DATAIN(28), ZN => n799);
   U652 : INV_X1 port map( A => DATAIN(29), ZN => n801);
   U653 : INV_X1 port map( A => DATAIN(30), ZN => n803);
   U654 : INV_X1 port map( A => DATAIN(31), ZN => n805);
   U655 : INV_X1 port map( A => DATAIN(32), ZN => n807);
   U656 : INV_X1 port map( A => DATAIN(33), ZN => n809);
   U657 : INV_X1 port map( A => DATAIN(34), ZN => n811);
   U658 : INV_X1 port map( A => DATAIN(35), ZN => n813);
   U659 : INV_X1 port map( A => DATAIN(36), ZN => n815);
   U660 : INV_X1 port map( A => DATAIN(37), ZN => n817);
   U661 : INV_X1 port map( A => DATAIN(38), ZN => n819);
   U662 : INV_X1 port map( A => DATAIN(39), ZN => n821);
   U663 : INV_X1 port map( A => DATAIN(40), ZN => n823);
   U664 : INV_X1 port map( A => DATAIN(41), ZN => n825);
   U665 : INV_X1 port map( A => DATAIN(42), ZN => n827);
   U666 : INV_X1 port map( A => DATAIN(43), ZN => n829);
   U667 : INV_X1 port map( A => DATAIN(44), ZN => n831);
   U668 : INV_X1 port map( A => DATAIN(45), ZN => n833);
   U669 : INV_X1 port map( A => DATAIN(46), ZN => n835);
   U670 : INV_X1 port map( A => DATAIN(47), ZN => n837);
   U671 : INV_X1 port map( A => DATAIN(48), ZN => n839);
   U672 : INV_X1 port map( A => DATAIN(49), ZN => n841);
   U673 : INV_X1 port map( A => DATAIN(50), ZN => n843);
   U674 : INV_X1 port map( A => DATAIN(51), ZN => n845);
   U675 : INV_X1 port map( A => DATAIN(52), ZN => n847);
   U676 : INV_X1 port map( A => DATAIN(53), ZN => n849);
   U677 : INV_X1 port map( A => DATAIN(54), ZN => n851);
   U678 : INV_X1 port map( A => DATAIN(55), ZN => n853);
   U679 : INV_X1 port map( A => DATAIN(56), ZN => n855);
   U680 : INV_X1 port map( A => DATAIN(57), ZN => n857);
   U681 : INV_X1 port map( A => DATAIN(58), ZN => n859);
   U682 : INV_X1 port map( A => DATAIN(59), ZN => n861);
   U683 : INV_X1 port map( A => DATAIN(60), ZN => n863);
   U684 : INV_X1 port map( A => DATAIN(61), ZN => n865);
   U685 : INV_X1 port map( A => DATAIN(62), ZN => n867);
   U686 : INV_X1 port map( A => DATAIN(63), ZN => n871);
   U687 : CLKBUF_X1 port map( A => n979, Z => n2069);
   U688 : CLKBUF_X1 port map( A => n978, Z => n2075);
   U689 : CLKBUF_X1 port map( A => n939, Z => n2081);
   U690 : CLKBUF_X1 port map( A => n938, Z => n2087);
   U691 : CLKBUF_X1 port map( A => n876, Z => n2093);
   U692 : CLKBUF_X1 port map( A => n875, Z => n2099);
   U693 : CLKBUF_X1 port map( A => n742, Z => n2105);
   U694 : CLKBUF_X1 port map( A => n741, Z => n2111);
   U695 : CLKBUF_X1 port map( A => n740, Z => n2117);
   U696 : CLKBUF_X1 port map( A => n739, Z => n2123);
   U697 : CLKBUF_X1 port map( A => n738, Z => n2129);
   U698 : CLKBUF_X1 port map( A => n736, Z => n2135);
   U699 : CLKBUF_X1 port map( A => n735, Z => n2141);
   U700 : CLKBUF_X1 port map( A => n527, Z => n2147);
   U701 : CLKBUF_X1 port map( A => n525, Z => n2158);
   U702 : CLKBUF_X1 port map( A => n523, Z => n2164);
   U703 : CLKBUF_X1 port map( A => n521, Z => n2170);
   U704 : INV_X1 port map( A => ADD_RD2(0), ZN => n2171);
   U705 : INV_X1 port map( A => ADD_RD2(1), ZN => n2172);
   U706 : INV_X1 port map( A => ADD_RD1(0), ZN => n2173);
   U707 : INV_X1 port map( A => ADD_RD1(1), ZN => n2174);
   U708 : INV_X1 port map( A => ADD_WR(0), ZN => n2175);
   U709 : INV_X1 port map( A => ADD_WR(1), ZN => n2176);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4.all;

entity register_file_reg_size64_file_size4_2 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_reg_size64_file_size4_2;

architecture SYN_BEHAVIORAL of register_file_reg_size64_file_size4_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n415, n1200, n1202, n1204, n1310, n1311, n1312, n1313, n1314, n1315
      , n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n871, n872, 
      n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, 
      n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, 
      n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, 
      n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, 
      n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, 
      n933, n934, n935, n936, n938, n939, n940, n941, n942, n943, n944, n945, 
      n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, 
      n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, 
      n970, n971, n972, n973, n974, n975, n977, n978, n979, n980, n981, n982, 
      n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, 
      n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, 
      n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, 
      n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, 
      n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, 
      n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, 
      n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, 
      n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062 : 
      std_logic;

begin
   
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => n174,
                           QN => n997);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => n175,
                           QN => n996);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => n176,
                           QN => n995);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => n177,
                           QN => n994);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => n178,
                           QN => n993);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => n179,
                           QN => n992);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => n180,
                           QN => n991);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => n181,
                           QN => n990);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => n182,
                           QN => n989);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => n183, 
                           QN => n988);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => n184, 
                           QN => n987);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => n185, 
                           QN => n986);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => n186, 
                           QN => n985);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => n187, 
                           QN => n984);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => n188, 
                           QN => n983);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => n189, 
                           QN => n982);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => n190, 
                           QN => n981);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => n191, 
                           QN => n980);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => n192, 
                           QN => n977);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => n65, 
                           QN => n974);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => n66, 
                           QN => n973);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n67, 
                           QN => n972);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => n68, 
                           QN => n971);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => n69, 
                           QN => n970);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => n70, 
                           QN => n969);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => n71, 
                           QN => n968);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => n72, 
                           QN => n967);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => n73, 
                           QN => n966);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => n74, 
                           QN => n965);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => n75, 
                           QN => n964);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => n76, 
                           QN => n963);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => n77, 
                           QN => n962);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => n78, 
                           QN => n961);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => n79, 
                           QN => n960);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => n80, 
                           QN => n959);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => n81, 
                           QN => n958);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => n82, 
                           QN => n957);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => n83, 
                           QN => n956);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => n84, 
                           QN => n955);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => n85, 
                           QN => n954);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => n86, 
                           QN => n953);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => n87, 
                           QN => n952);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => n88, 
                           QN => n951);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => n89, 
                           QN => n950);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => n90, 
                           QN => n949);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => n91, 
                           QN => n948);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => n92, 
                           QN => n947);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => n93, 
                           QN => n946);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => n94, 
                           QN => n945);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => n95, 
                           QN => n944);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => n96, 
                           QN => n943);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => n97, 
                           QN => n942);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => n98, 
                           QN => n941);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => n99, 
                           QN => n940);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => n2, 
                           QN => n935);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => n3, 
                           QN => n934);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => n4, 
                           QN => n933);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => n5, 
                           QN => n932);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => n6, 
                           QN => n931);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => n7, 
                           QN => n930);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => n8, 
                           QN => n929);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => n9, 
                           QN => n928);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => n13, 
                           QN => n927);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => n14, 
                           QN => n926);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => n15, 
                           QN => n925);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => n16, 
                           QN => n924);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => n17, 
                           QN => n923);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => n18, 
                           QN => n922);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => n19, 
                           QN => n921);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => n20, 
                           QN => n920);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => n21, 
                           QN => n919);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => n22, 
                           QN => n918);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => n23, 
                           QN => n917);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => n24, 
                           QN => n916);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => n25, 
                           QN => n915);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => n26, 
                           QN => n914);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n27, 
                           QN => n913);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => n28, 
                           QN => n912);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n29, 
                           QN => n911);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => n30, 
                           QN => n910);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n31, 
                           QN => n909);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => n32, 
                           QN => n908);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n33, 
                           QN => n907);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => n34, 
                           QN => n906);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n35, 
                           QN => n905);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => n36, 
                           QN => n904);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => n37, 
                           QN => n903);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => n38, 
                           QN => n902);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => n39, 
                           QN => n901);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => n40, 
                           QN => n900);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => n41, 
                           QN => n899);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => n42, 
                           QN => n898);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => n43, 
                           QN => n897);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => n44, 
                           QN => n896);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => n45, 
                           QN => n895);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => n46, 
                           QN => n894);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => n47, 
                           QN => n893);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => n48, 
                           QN => n892);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => n49, 
                           QN => n891);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => n50, 
                           QN => n890);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => n51, 
                           QN => n889);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => n52, 
                           QN => n888);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => n53, 
                           QN => n887);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => n54, 
                           QN => n886);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n55, 
                           QN => n885);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => n56, 
                           QN => n884);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n57, 
                           QN => n883);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => n58, 
                           QN => n882);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n59, 
                           QN => n881);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => n60, 
                           QN => n880);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n61, 
                           QN => n879);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => n62, 
                           QN => n878);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n63, 
                           QN => n877);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => n64, 
                           QN => n874);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n999,
                           QN => n728);
   OUT2_reg_63_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => OUT2(63), QN
                           => n1822);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n1000
                           , QN => n725);
   OUT2_reg_62_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => OUT2(62), QN
                           => n1823);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n1001
                           , QN => n722);
   OUT2_reg_61_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => OUT2(61), QN
                           => n1824);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n1002
                           , QN => n719);
   OUT2_reg_60_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => OUT2(60), QN
                           => n1825);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n1003
                           , QN => n716);
   OUT2_reg_59_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => OUT2(59), QN
                           => n1826);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n1004
                           , QN => n713);
   OUT2_reg_58_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => OUT2(58), QN
                           => n1827);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n1005
                           , QN => n710);
   OUT2_reg_57_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => OUT2(57), QN
                           => n1828);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n1006
                           , QN => n707);
   OUT2_reg_56_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => OUT2(56), QN
                           => n1829);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n1007
                           , QN => n704);
   OUT2_reg_55_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => OUT2(55), QN
                           => n1830);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n1008
                           , QN => n700);
   OUT2_reg_54_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => OUT2(54), QN
                           => n1831);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n1009
                           , QN => n696);
   OUT2_reg_53_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => OUT2(53), QN
                           => n1832);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n1010
                           , QN => n692);
   OUT2_reg_52_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => OUT2(52), QN
                           => n1833);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n1011
                           , QN => n689);
   OUT2_reg_51_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => OUT2(51), QN
                           => n1834);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n1012
                           , QN => n686);
   OUT2_reg_50_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => OUT2(50), QN
                           => n1835);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n1013
                           , QN => n683);
   OUT2_reg_49_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => OUT2(49), QN
                           => n1836);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n1014
                           , QN => n680);
   OUT2_reg_48_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => OUT2(48), QN
                           => n1837);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n1015
                           , QN => n677);
   OUT2_reg_47_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => OUT2(47), QN
                           => n1838);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n1016
                           , QN => n674);
   OUT2_reg_46_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => OUT2(46), QN
                           => n1839);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n1017
                           , QN => n671);
   OUT2_reg_45_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => OUT2(45), QN
                           => n1840);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n1018
                           , QN => n668);
   OUT2_reg_44_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => OUT2(44), QN
                           => n1841);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n1019
                           , QN => n665);
   OUT2_reg_43_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => OUT2(43), QN
                           => n1842);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n1020
                           , QN => n662);
   OUT2_reg_42_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => OUT2(42), QN
                           => n1843);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n1021
                           , QN => n659);
   OUT2_reg_41_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => OUT2(41), QN
                           => n1844);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n1022
                           , QN => n656);
   OUT2_reg_40_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => OUT2(40), QN
                           => n1845);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n1023
                           , QN => n653);
   OUT2_reg_39_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => OUT2(39), QN
                           => n1846);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n1024
                           , QN => n650);
   OUT2_reg_38_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => OUT2(38), QN
                           => n1847);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n1025
                           , QN => n647);
   OUT2_reg_37_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => OUT2(37), QN
                           => n1848);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n1026
                           , QN => n644);
   OUT2_reg_36_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => OUT2(36), QN
                           => n1849);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n1027
                           , QN => n641);
   OUT2_reg_35_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => OUT2(35), QN
                           => n1850);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n1028
                           , QN => n638);
   OUT2_reg_34_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => OUT2(34), QN
                           => n1851);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n1029
                           , QN => n635);
   OUT2_reg_33_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => OUT2(33), QN
                           => n1852);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n1030
                           , QN => n632);
   OUT2_reg_32_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => OUT2(32), QN
                           => n1853);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n1031
                           , QN => n629);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => OUT2(31), QN
                           => n1854);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n1032
                           , QN => n626);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => OUT2(30), QN
                           => n1855);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n1033
                           , QN => n623);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => OUT2(29), QN
                           => n1856);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n1034
                           , QN => n619);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => OUT2(28), QN
                           => n1857);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n1035
                           , QN => n615);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => OUT2(27), QN
                           => n1858);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n1036
                           , QN => n611);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => OUT2(26), QN
                           => n1859);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n1037
                           , QN => n607);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => OUT2(25), QN
                           => n1860);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n1038
                           , QN => n603);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => OUT2(24), QN
                           => n1861);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n1039
                           , QN => n599);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => OUT2(23), QN
                           => n1862);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n1040
                           , QN => n595);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => OUT2(22), QN
                           => n1863);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n1041
                           , QN => n591);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => OUT2(21), QN
                           => n1864);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n1042
                           , QN => n587);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => OUT2(20), QN
                           => n1865);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n1043
                           , QN => n583);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => OUT2(19), QN
                           => n1866);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n1044
                           , QN => n580);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => OUT2(18), QN
                           => n1867);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n1045
                           , QN => n577);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => OUT2(17), QN
                           => n1868);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n1046
                           , QN => n574);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => OUT2(16), QN
                           => n1869);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n1047
                           , QN => n571);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => OUT2(15), QN
                           => n1870);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n1048
                           , QN => n568);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => OUT2(14), QN
                           => n1871);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n1049
                           , QN => n565);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => OUT2(13), QN
                           => n1872);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n1050
                           , QN => n562);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => OUT2(12), QN
                           => n1873);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n1051
                           , QN => n559);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => OUT2(11), QN
                           => n1874);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n1052
                           , QN => n556);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => OUT2(10), QN
                           => n1875);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n1053,
                           QN => n553);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => OUT2(9), QN 
                           => n1876);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => n1054,
                           QN => n550);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => OUT2(8), QN 
                           => n1877);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => n1055,
                           QN => n547);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => OUT2(7), QN 
                           => n1878);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => n1056,
                           QN => n544);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => OUT2(6), QN 
                           => n1879);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => n1057,
                           QN => n541);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => OUT2(5), QN 
                           => n1880);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => n1058,
                           QN => n538);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => OUT2(4), QN 
                           => n1881);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => n1059,
                           QN => n535);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => OUT2(3), QN 
                           => n1882);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n1060,
                           QN => n532);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => OUT2(2), QN 
                           => n1883);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n1061,
                           QN => n529);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => OUT2(1), QN 
                           => n1884);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n1062,
                           QN => n522);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => OUT2(0), QN 
                           => n1885);
   OUT1_reg_63_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => OUT1(63), QN
                           => n1886);
   OUT1_reg_62_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => OUT1(62), QN
                           => n1887);
   OUT1_reg_61_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => OUT1(61), QN
                           => n1888);
   OUT1_reg_60_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => OUT1(60), QN
                           => n1889);
   OUT1_reg_59_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => OUT1(59), QN
                           => n1890);
   OUT1_reg_58_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => OUT1(58), QN
                           => n1891);
   OUT1_reg_57_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => OUT1(57), QN
                           => n1892);
   OUT1_reg_56_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => OUT1(56), QN
                           => n1893);
   OUT1_reg_55_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => OUT1(55), QN
                           => n1894);
   OUT1_reg_54_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => OUT1(54), QN
                           => n1895);
   OUT1_reg_53_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => OUT1(53), QN
                           => n1896);
   OUT1_reg_52_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => OUT1(52), QN
                           => n1897);
   OUT1_reg_51_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => OUT1(51), QN
                           => n1898);
   OUT1_reg_50_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => OUT1(50), QN
                           => n1899);
   OUT1_reg_49_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => OUT1(49), QN
                           => n1900);
   OUT1_reg_48_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => OUT1(48), QN
                           => n1901);
   OUT1_reg_47_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => OUT1(47), QN
                           => n1902);
   OUT1_reg_46_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => OUT1(46), QN
                           => n1903);
   OUT1_reg_45_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => OUT1(45), QN
                           => n1904);
   OUT1_reg_44_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => OUT1(44), QN
                           => n1905);
   OUT1_reg_43_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => OUT1(43), QN
                           => n1906);
   OUT1_reg_42_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => OUT1(42), QN
                           => n1907);
   OUT1_reg_41_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => OUT1(41), QN
                           => n1908);
   OUT1_reg_40_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => OUT1(40), QN
                           => n1909);
   OUT1_reg_39_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => OUT1(39), QN
                           => n1910);
   OUT1_reg_38_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => OUT1(38), QN
                           => n1911);
   OUT1_reg_37_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => OUT1(37), QN
                           => n1912);
   OUT1_reg_36_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => OUT1(36), QN
                           => n1913);
   OUT1_reg_35_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => OUT1(35), QN
                           => n1914);
   OUT1_reg_34_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => OUT1(34), QN
                           => n1915);
   OUT1_reg_33_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => OUT1(33), QN
                           => n1916);
   OUT1_reg_32_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => OUT1(32), QN
                           => n1917);
   OUT1_reg_31_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => OUT1(31), QN
                           => n1918);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => OUT1(30), QN
                           => n1919);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => OUT1(29), QN
                           => n1920);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => OUT1(28), QN
                           => n1921);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => OUT1(27), QN
                           => n1922);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => OUT1(26), QN
                           => n1923);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => OUT1(25), QN
                           => n1924);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => OUT1(24), QN
                           => n1925);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => OUT1(23), QN
                           => n1926);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => OUT1(22), QN
                           => n1927);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => OUT1(21), QN
                           => n1928);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => OUT1(20), QN
                           => n1929);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => OUT1(19), QN
                           => n1930);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => OUT1(18), QN
                           => n1931);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => OUT1(17), QN
                           => n1932);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => OUT1(16), QN
                           => n1933);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => OUT1(15), QN
                           => n1934);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => OUT1(14), QN
                           => n1935);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => OUT1(13), QN
                           => n1936);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => OUT1(12), QN
                           => n1937);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => OUT1(11), QN
                           => n1938);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => OUT1(10), QN
                           => n1939);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => OUT1(9), QN 
                           => n1940);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => OUT1(8), QN 
                           => n1941);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => OUT1(7), QN 
                           => n1942);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => OUT1(6), QN 
                           => n1943);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => OUT1(5), QN 
                           => n1944);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => OUT1(4), QN 
                           => n1945);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => OUT1(3), QN 
                           => n1946);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => OUT1(2), QN 
                           => n1947);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => OUT1(1), QN 
                           => n1948);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => OUT1(0), QN 
                           => n1949);
   U859 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n2050, A3 => ADD_RD1(1), 
                           ZN => n521);
   U860 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n2021, A3 => ADD_RD2(1), 
                           ZN => n735);
   U861 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n873, A3 => ADD_WR(1), ZN 
                           => n872);
   U862 : NAND3_X1 port map( A1 => n873, A2 => n2061, A3 => ADD_WR(1), ZN => 
                           n936);
   U863 : NAND3_X1 port map( A1 => n873, A2 => n2062, A3 => ADD_WR(0), ZN => 
                           n975);
   U864 : NAND3_X1 port map( A1 => n2061, A2 => n2062, A3 => n873, ZN => n998);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => n537, 
                           QN => n1818);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => n534, 
                           QN => n1819);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => n531, 
                           QN => n1820);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => n528, 
                           QN => n1821);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => n730,
                           QN => n415);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => n702,
                           QN => n1200);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => n698,
                           QN => n1202);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => n694,
                           QN => n1204);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => n622,
                           QN => n1793);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => n618,
                           QN => n1794);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => n614,
                           QN => n1795);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => n610,
                           QN => n1796);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => n606,
                           QN => n1797);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => n602,
                           QN => n1798);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => n598,
                           QN => n1799);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => n594,
                           QN => n1800);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => n590,
                           QN => n1801);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => n586,
                           QN => n1802);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => n582,
                           QN => n1803);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => n579,
                           QN => n1804);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => n576,
                           QN => n1805);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => n573,
                           QN => n1806);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => n570,
                           QN => n1807);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => n567,
                           QN => n1808);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => n564,
                           QN => n1809);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => n561,
                           QN => n1810);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => n558,
                           QN => n1811);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => n555, 
                           QN => n1812);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => n552, 
                           QN => n1813);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => n549, 
                           QN => n1814);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => n546, 
                           QN => n1815);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => n543, 
                           QN => n1816);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => n540, 
                           QN => n1817);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => n731,
                           QN => n1694);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => n727,
                           QN => n1695);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => n724,
                           QN => n1696);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => n721,
                           QN => n1697);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => n718,
                           QN => n1698);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => n715,
                           QN => n1699);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => n712,
                           QN => n1700);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => n709,
                           QN => n1701);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => n706,
                           QN => n1702);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => n703,
                           QN => n1703);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => n699,
                           QN => n1704);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => n695,
                           QN => n1705);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => n691,
                           QN => n1706);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => n688,
                           QN => n1707);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => n685,
                           QN => n1708);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => n682,
                           QN => n1709);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => n679,
                           QN => n1710);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => n676,
                           QN => n1711);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => n673,
                           QN => n1712);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => n670,
                           QN => n1713);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => n667,
                           QN => n1714);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => n664,
                           QN => n1715);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => n661,
                           QN => n1716);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => n658,
                           QN => n1717);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => n655,
                           QN => n1718);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => n652,
                           QN => n1719);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => n649,
                           QN => n1720);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => n646,
                           QN => n1721);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => n643,
                           QN => n1722);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => n640,
                           QN => n1723);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => n637,
                           QN => n1724);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => n634,
                           QN => n1725);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => n631,
                           QN => n1726);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => n628,
                           QN => n1727);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n625,
                           QN => n1728);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => n621,
                           QN => n1729);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => n617,
                           QN => n1730);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => n613,
                           QN => n1731);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => n609,
                           QN => n1732);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => n605,
                           QN => n1733);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => n601,
                           QN => n1734);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => n597,
                           QN => n1735);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => n593,
                           QN => n1736);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => n589,
                           QN => n1737);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => n585,
                           QN => n1738);
   U3 : BUF_X1 port map( A => n521, Z => n2053);
   U4 : BUF_X1 port map( A => n521, Z => n2052);
   U5 : BUF_X1 port map( A => n521, Z => n2051);
   U6 : BUF_X1 port map( A => n735, Z => n2025);
   U7 : BUF_X1 port map( A => n735, Z => n2024);
   U8 : BUF_X1 port map( A => n735, Z => n2023);
   U9 : BUF_X1 port map( A => n735, Z => n2022);
   U10 : BUF_X1 port map( A => n521, Z => n2055);
   U11 : BUF_X1 port map( A => n521, Z => n2054);
   U12 : BUF_X1 port map( A => n735, Z => n2026);
   U13 : BUF_X1 port map( A => n742, Z => n1990);
   U14 : BUF_X1 port map( A => n742, Z => n1989);
   U15 : BUF_X1 port map( A => n742, Z => n1988);
   U16 : BUF_X1 port map( A => n742, Z => n1987);
   U17 : BUF_X1 port map( A => n741, Z => n1992);
   U18 : BUF_X1 port map( A => n875, Z => n1980);
   U19 : BUF_X1 port map( A => n938, Z => n1968);
   U20 : BUF_X1 port map( A => n978, Z => n1956);
   U21 : BUF_X1 port map( A => n876, Z => n1978);
   U22 : BUF_X1 port map( A => n876, Z => n1977);
   U23 : BUF_X1 port map( A => n876, Z => n1976);
   U24 : BUF_X1 port map( A => n876, Z => n1975);
   U25 : BUF_X1 port map( A => n876, Z => n1974);
   U26 : BUF_X1 port map( A => n939, Z => n1966);
   U27 : BUF_X1 port map( A => n939, Z => n1965);
   U28 : BUF_X1 port map( A => n939, Z => n1964);
   U29 : BUF_X1 port map( A => n939, Z => n1963);
   U30 : BUF_X1 port map( A => n939, Z => n1962);
   U31 : BUF_X1 port map( A => n979, Z => n1954);
   U32 : BUF_X1 port map( A => n979, Z => n1953);
   U33 : BUF_X1 port map( A => n979, Z => n1952);
   U34 : BUF_X1 port map( A => n979, Z => n1951);
   U35 : BUF_X1 port map( A => n979, Z => n1950);
   U36 : BUF_X1 port map( A => n742, Z => n1986);
   U37 : BUF_X1 port map( A => n526, Z => n2037);
   U38 : BUF_X1 port map( A => n526, Z => n2038);
   U39 : BUF_X1 port map( A => n527, Z => n2030);
   U40 : BUF_X1 port map( A => n527, Z => n2032);
   U41 : BUF_X1 port map( A => n527, Z => n2031);
   U42 : BUF_X1 port map( A => n523, Z => n2045);
   U43 : BUF_X1 port map( A => n523, Z => n2046);
   U44 : BUF_X1 port map( A => n523, Z => n2047);
   U45 : BUF_X1 port map( A => n523, Z => n2048);
   U46 : BUF_X1 port map( A => n523, Z => n2049);
   U47 : BUF_X1 port map( A => n736, Z => n2016);
   U48 : BUF_X1 port map( A => n736, Z => n2017);
   U49 : BUF_X1 port map( A => n736, Z => n2018);
   U50 : BUF_X1 port map( A => n736, Z => n2019);
   U51 : BUF_X1 port map( A => n736, Z => n2020);
   U52 : BUF_X1 port map( A => n525, Z => n2040);
   U53 : BUF_X1 port map( A => n525, Z => n2041);
   U54 : BUF_X1 port map( A => n525, Z => n2042);
   U55 : BUF_X1 port map( A => n525, Z => n2043);
   U56 : BUF_X1 port map( A => n738, Z => n2014);
   U57 : BUF_X1 port map( A => n738, Z => n2013);
   U58 : BUF_X1 port map( A => n738, Z => n2012);
   U59 : BUF_X1 port map( A => n738, Z => n2011);
   U60 : BUF_X1 port map( A => n738, Z => n2010);
   U61 : BUF_X1 port map( A => n739, Z => n2008);
   U62 : BUF_X1 port map( A => n739, Z => n2007);
   U63 : BUF_X1 port map( A => n739, Z => n2006);
   U64 : BUF_X1 port map( A => n739, Z => n2005);
   U65 : BUF_X1 port map( A => n739, Z => n2004);
   U66 : BUF_X1 port map( A => n740, Z => n2002);
   U67 : BUF_X1 port map( A => n740, Z => n2001);
   U68 : BUF_X1 port map( A => n740, Z => n2000);
   U69 : BUF_X1 port map( A => n740, Z => n1999);
   U70 : BUF_X1 port map( A => n740, Z => n1998);
   U71 : BUF_X1 port map( A => n741, Z => n1996);
   U72 : BUF_X1 port map( A => n741, Z => n1995);
   U73 : BUF_X1 port map( A => n741, Z => n1994);
   U74 : BUF_X1 port map( A => n741, Z => n1993);
   U75 : BUF_X1 port map( A => n875, Z => n1984);
   U76 : BUF_X1 port map( A => n875, Z => n1983);
   U77 : BUF_X1 port map( A => n875, Z => n1982);
   U78 : BUF_X1 port map( A => n875, Z => n1981);
   U79 : BUF_X1 port map( A => n938, Z => n1972);
   U80 : BUF_X1 port map( A => n938, Z => n1971);
   U81 : BUF_X1 port map( A => n938, Z => n1970);
   U82 : BUF_X1 port map( A => n938, Z => n1969);
   U83 : BUF_X1 port map( A => n978, Z => n1960);
   U84 : BUF_X1 port map( A => n978, Z => n1959);
   U85 : BUF_X1 port map( A => n978, Z => n1958);
   U86 : BUF_X1 port map( A => n978, Z => n1957);
   U87 : BUF_X1 port map( A => n526, Z => n2034);
   U88 : BUF_X1 port map( A => n526, Z => n2036);
   U89 : BUF_X1 port map( A => n527, Z => n2029);
   U90 : BUF_X1 port map( A => n527, Z => n2028);
   U91 : BUF_X1 port map( A => n526, Z => n2035);
   U92 : BUF_X1 port map( A => n525, Z => n2039);
   U93 : NAND2_X1 port map( A1 => n734, A2 => n872, ZN => n741);
   U94 : NAND2_X1 port map( A1 => n734, A2 => n936, ZN => n875);
   U95 : NAND2_X1 port map( A1 => n734, A2 => n1980, ZN => n876);
   U96 : NAND2_X1 port map( A1 => n734, A2 => n975, ZN => n938);
   U97 : NAND2_X1 port map( A1 => n734, A2 => n1968, ZN => n939);
   U98 : NAND2_X1 port map( A1 => n734, A2 => n998, ZN => n978);
   U99 : NAND2_X1 port map( A1 => n734, A2 => n1956, ZN => n979);
   U100 : OAI22_X1 port map( A1 => n538, A2 => n1997, B1 => n1990, B2 => n751, 
                           ZN => n1620);
   U101 : OAI22_X1 port map( A1 => n541, A2 => n1996, B1 => n1990, B2 => n753, 
                           ZN => n1618);
   U102 : OAI22_X1 port map( A1 => n544, A2 => n1996, B1 => n1990, B2 => n755, 
                           ZN => n1616);
   U103 : OAI22_X1 port map( A1 => n547, A2 => n1996, B1 => n1990, B2 => n757, 
                           ZN => n1614);
   U104 : OAI22_X1 port map( A1 => n550, A2 => n1996, B1 => n1990, B2 => n759, 
                           ZN => n1612);
   U105 : OAI22_X1 port map( A1 => n553, A2 => n1996, B1 => n1990, B2 => n761, 
                           ZN => n1610);
   U106 : OAI22_X1 port map( A1 => n556, A2 => n1996, B1 => n1990, B2 => n763, 
                           ZN => n1608);
   U107 : OAI22_X1 port map( A1 => n559, A2 => n1996, B1 => n1990, B2 => n765, 
                           ZN => n1606);
   U108 : OAI22_X1 port map( A1 => n562, A2 => n1996, B1 => n1990, B2 => n767, 
                           ZN => n1604);
   U109 : OAI22_X1 port map( A1 => n565, A2 => n1996, B1 => n1990, B2 => n769, 
                           ZN => n1602);
   U110 : OAI22_X1 port map( A1 => n568, A2 => n1996, B1 => n1990, B2 => n771, 
                           ZN => n1600);
   U111 : OAI22_X1 port map( A1 => n571, A2 => n1996, B1 => n1990, B2 => n773, 
                           ZN => n1598);
   U112 : OAI22_X1 port map( A1 => n574, A2 => n1996, B1 => n1989, B2 => n775, 
                           ZN => n1596);
   U113 : OAI22_X1 port map( A1 => n577, A2 => n1995, B1 => n1989, B2 => n777, 
                           ZN => n1594);
   U114 : OAI22_X1 port map( A1 => n580, A2 => n1995, B1 => n1989, B2 => n779, 
                           ZN => n1592);
   U115 : OAI22_X1 port map( A1 => n583, A2 => n1995, B1 => n1989, B2 => n781, 
                           ZN => n1590);
   U116 : OAI22_X1 port map( A1 => n587, A2 => n1995, B1 => n1989, B2 => n783, 
                           ZN => n1588);
   U117 : OAI22_X1 port map( A1 => n591, A2 => n1995, B1 => n1989, B2 => n785, 
                           ZN => n1586);
   U118 : OAI22_X1 port map( A1 => n595, A2 => n1995, B1 => n1989, B2 => n787, 
                           ZN => n1584);
   U119 : OAI22_X1 port map( A1 => n599, A2 => n1995, B1 => n1989, B2 => n789, 
                           ZN => n1582);
   U120 : OAI22_X1 port map( A1 => n603, A2 => n1995, B1 => n1989, B2 => n791, 
                           ZN => n1580);
   U121 : OAI22_X1 port map( A1 => n607, A2 => n1995, B1 => n1989, B2 => n793, 
                           ZN => n1578);
   U122 : OAI22_X1 port map( A1 => n611, A2 => n1995, B1 => n1989, B2 => n795, 
                           ZN => n1576);
   U123 : OAI22_X1 port map( A1 => n615, A2 => n1995, B1 => n1989, B2 => n797, 
                           ZN => n1574);
   U124 : OAI22_X1 port map( A1 => n619, A2 => n1995, B1 => n1988, B2 => n799, 
                           ZN => n1572);
   U125 : OAI22_X1 port map( A1 => n623, A2 => n1994, B1 => n1988, B2 => n801, 
                           ZN => n1570);
   U126 : OAI22_X1 port map( A1 => n626, A2 => n1994, B1 => n1988, B2 => n803, 
                           ZN => n1568);
   U127 : OAI22_X1 port map( A1 => n629, A2 => n1994, B1 => n1988, B2 => n805, 
                           ZN => n1566);
   U128 : OAI22_X1 port map( A1 => n632, A2 => n1994, B1 => n1988, B2 => n807, 
                           ZN => n1564);
   U129 : OAI22_X1 port map( A1 => n635, A2 => n1994, B1 => n1988, B2 => n809, 
                           ZN => n1562);
   U130 : OAI22_X1 port map( A1 => n638, A2 => n1994, B1 => n1988, B2 => n811, 
                           ZN => n1560);
   U131 : OAI22_X1 port map( A1 => n641, A2 => n1994, B1 => n1988, B2 => n813, 
                           ZN => n1558);
   U132 : OAI22_X1 port map( A1 => n644, A2 => n1994, B1 => n1988, B2 => n815, 
                           ZN => n1556);
   U133 : OAI22_X1 port map( A1 => n647, A2 => n1994, B1 => n1988, B2 => n817, 
                           ZN => n1554);
   U134 : OAI22_X1 port map( A1 => n650, A2 => n1994, B1 => n1988, B2 => n819, 
                           ZN => n1552);
   U135 : OAI22_X1 port map( A1 => n653, A2 => n1994, B1 => n1988, B2 => n821, 
                           ZN => n1550);
   U136 : OAI22_X1 port map( A1 => n656, A2 => n1994, B1 => n1987, B2 => n823, 
                           ZN => n1548);
   U137 : OAI22_X1 port map( A1 => n659, A2 => n1993, B1 => n1987, B2 => n825, 
                           ZN => n1546);
   U138 : OAI22_X1 port map( A1 => n662, A2 => n1993, B1 => n1987, B2 => n827, 
                           ZN => n1544);
   U139 : OAI22_X1 port map( A1 => n665, A2 => n1993, B1 => n1987, B2 => n829, 
                           ZN => n1542);
   U140 : OAI22_X1 port map( A1 => n668, A2 => n1993, B1 => n1987, B2 => n831, 
                           ZN => n1540);
   U141 : OAI22_X1 port map( A1 => n671, A2 => n1993, B1 => n1987, B2 => n833, 
                           ZN => n1538);
   U142 : OAI22_X1 port map( A1 => n674, A2 => n1993, B1 => n1987, B2 => n835, 
                           ZN => n1536);
   U143 : OAI22_X1 port map( A1 => n677, A2 => n1993, B1 => n1987, B2 => n837, 
                           ZN => n1534);
   U144 : OAI22_X1 port map( A1 => n680, A2 => n1993, B1 => n1987, B2 => n839, 
                           ZN => n1532);
   U145 : OAI22_X1 port map( A1 => n683, A2 => n1993, B1 => n1987, B2 => n841, 
                           ZN => n1530);
   U146 : OAI22_X1 port map( A1 => n686, A2 => n1993, B1 => n1987, B2 => n843, 
                           ZN => n1528);
   U147 : OAI22_X1 port map( A1 => n689, A2 => n1993, B1 => n1987, B2 => n845, 
                           ZN => n1526);
   U148 : OAI22_X1 port map( A1 => n522, A2 => n1997, B1 => n1991, B2 => n743, 
                           ZN => n1628);
   U149 : OAI22_X1 port map( A1 => n529, A2 => n1997, B1 => n1991, B2 => n745, 
                           ZN => n1626);
   U150 : OAI22_X1 port map( A1 => n532, A2 => n1997, B1 => n1991, B2 => n747, 
                           ZN => n1624);
   U151 : OAI22_X1 port map( A1 => n535, A2 => n1997, B1 => n1991, B2 => n749, 
                           ZN => n1622);
   U152 : OAI22_X1 port map( A1 => n692, A2 => n1993, B1 => n1986, B2 => n847, 
                           ZN => n1524);
   U153 : OAI22_X1 port map( A1 => n696, A2 => n1992, B1 => n1986, B2 => n849, 
                           ZN => n1522);
   U154 : OAI22_X1 port map( A1 => n700, A2 => n1992, B1 => n1986, B2 => n851, 
                           ZN => n1520);
   U155 : OAI22_X1 port map( A1 => n704, A2 => n1992, B1 => n1986, B2 => n853, 
                           ZN => n1518);
   U156 : OAI22_X1 port map( A1 => n707, A2 => n1992, B1 => n1986, B2 => n855, 
                           ZN => n1516);
   U157 : OAI22_X1 port map( A1 => n710, A2 => n1992, B1 => n1986, B2 => n857, 
                           ZN => n1514);
   U158 : OAI22_X1 port map( A1 => n713, A2 => n1992, B1 => n1986, B2 => n859, 
                           ZN => n1512);
   U159 : OAI22_X1 port map( A1 => n716, A2 => n1992, B1 => n1986, B2 => n861, 
                           ZN => n1510);
   U160 : OAI22_X1 port map( A1 => n719, A2 => n1992, B1 => n1986, B2 => n863, 
                           ZN => n1508);
   U161 : OAI22_X1 port map( A1 => n722, A2 => n1992, B1 => n1986, B2 => n865, 
                           ZN => n1506);
   U162 : OAI22_X1 port map( A1 => n725, A2 => n1992, B1 => n1986, B2 => n867, 
                           ZN => n1504);
   U163 : OAI22_X1 port map( A1 => n728, A2 => n1992, B1 => n1986, B2 => n871, 
                           ZN => n1502);
   U164 : NAND2_X1 port map( A1 => n734, A2 => n1992, ZN => n742);
   U165 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n873);
   U166 : AND3_X1 port map( A1 => n2059, A2 => n2060, A3 => n2050, ZN => n526);
   U167 : AND3_X1 port map( A1 => n2050, A2 => n2060, A3 => ADD_RD1(0), ZN => 
                           n527);
   U168 : AND3_X1 port map( A1 => n2050, A2 => n2059, A3 => ADD_RD1(1), ZN => 
                           n525);
   U169 : AND3_X1 port map( A1 => n2021, A2 => n2058, A3 => ADD_RD2(0), ZN => 
                           n740);
   U170 : AND3_X1 port map( A1 => n2021, A2 => n2057, A3 => ADD_RD2(1), ZN => 
                           n738);
   U171 : AND3_X1 port map( A1 => n2057, A2 => n2058, A3 => n2021, ZN => n739);
   U172 : AND2_X1 port map( A1 => RD2, A2 => n734, ZN => n736);
   U173 : AND2_X1 port map( A1 => RD1, A2 => n734, ZN => n523);
   U174 : OAI22_X1 port map( A1 => n874, A2 => n1985, B1 => n743, B2 => n1979, 
                           ZN => n1501);
   U175 : OAI22_X1 port map( A1 => n877, A2 => n1985, B1 => n745, B2 => n1979, 
                           ZN => n1500);
   U176 : OAI22_X1 port map( A1 => n878, A2 => n1985, B1 => n747, B2 => n1979, 
                           ZN => n1499);
   U177 : OAI22_X1 port map( A1 => n879, A2 => n1985, B1 => n749, B2 => n1979, 
                           ZN => n1498);
   U178 : OAI22_X1 port map( A1 => n1821, A2 => n1973, B1 => n743, B2 => n1967,
                           ZN => n1437);
   U179 : OAI22_X1 port map( A1 => n1820, A2 => n1973, B1 => n745, B2 => n1967,
                           ZN => n1436);
   U180 : OAI22_X1 port map( A1 => n1819, A2 => n1973, B1 => n747, B2 => n1967,
                           ZN => n1435);
   U181 : OAI22_X1 port map( A1 => n1818, A2 => n1973, B1 => n749, B2 => n1967,
                           ZN => n1434);
   U182 : OAI22_X1 port map( A1 => n977, A2 => n1961, B1 => n743, B2 => n1955, 
                           ZN => n1373);
   U183 : OAI22_X1 port map( A1 => n980, A2 => n1961, B1 => n745, B2 => n1955, 
                           ZN => n1372);
   U184 : OAI22_X1 port map( A1 => n981, A2 => n1961, B1 => n747, B2 => n1955, 
                           ZN => n1371);
   U185 : OAI22_X1 port map( A1 => n982, A2 => n1961, B1 => n749, B2 => n1955, 
                           ZN => n1370);
   U186 : OAI22_X1 port map( A1 => n880, A2 => n1985, B1 => n751, B2 => n1978, 
                           ZN => n1497);
   U187 : OAI22_X1 port map( A1 => n881, A2 => n1984, B1 => n753, B2 => n1978, 
                           ZN => n1496);
   U188 : OAI22_X1 port map( A1 => n882, A2 => n1984, B1 => n755, B2 => n1978, 
                           ZN => n1495);
   U189 : OAI22_X1 port map( A1 => n883, A2 => n1984, B1 => n757, B2 => n1978, 
                           ZN => n1494);
   U190 : OAI22_X1 port map( A1 => n884, A2 => n1984, B1 => n759, B2 => n1978, 
                           ZN => n1493);
   U191 : OAI22_X1 port map( A1 => n885, A2 => n1984, B1 => n761, B2 => n1978, 
                           ZN => n1492);
   U192 : OAI22_X1 port map( A1 => n886, A2 => n1984, B1 => n763, B2 => n1978, 
                           ZN => n1491);
   U193 : OAI22_X1 port map( A1 => n887, A2 => n1984, B1 => n765, B2 => n1978, 
                           ZN => n1490);
   U194 : OAI22_X1 port map( A1 => n888, A2 => n1984, B1 => n767, B2 => n1978, 
                           ZN => n1489);
   U195 : OAI22_X1 port map( A1 => n889, A2 => n1984, B1 => n769, B2 => n1978, 
                           ZN => n1488);
   U196 : OAI22_X1 port map( A1 => n890, A2 => n1984, B1 => n771, B2 => n1978, 
                           ZN => n1487);
   U197 : OAI22_X1 port map( A1 => n891, A2 => n1984, B1 => n773, B2 => n1978, 
                           ZN => n1486);
   U198 : OAI22_X1 port map( A1 => n892, A2 => n1984, B1 => n775, B2 => n1977, 
                           ZN => n1485);
   U199 : OAI22_X1 port map( A1 => n893, A2 => n1983, B1 => n777, B2 => n1977, 
                           ZN => n1484);
   U200 : OAI22_X1 port map( A1 => n894, A2 => n1983, B1 => n779, B2 => n1977, 
                           ZN => n1483);
   U201 : OAI22_X1 port map( A1 => n895, A2 => n1983, B1 => n781, B2 => n1977, 
                           ZN => n1482);
   U202 : OAI22_X1 port map( A1 => n896, A2 => n1983, B1 => n783, B2 => n1977, 
                           ZN => n1481);
   U203 : OAI22_X1 port map( A1 => n897, A2 => n1983, B1 => n785, B2 => n1977, 
                           ZN => n1480);
   U204 : OAI22_X1 port map( A1 => n898, A2 => n1983, B1 => n787, B2 => n1977, 
                           ZN => n1479);
   U205 : OAI22_X1 port map( A1 => n899, A2 => n1983, B1 => n789, B2 => n1977, 
                           ZN => n1478);
   U206 : OAI22_X1 port map( A1 => n900, A2 => n1983, B1 => n791, B2 => n1977, 
                           ZN => n1477);
   U207 : OAI22_X1 port map( A1 => n901, A2 => n1983, B1 => n793, B2 => n1977, 
                           ZN => n1476);
   U208 : OAI22_X1 port map( A1 => n902, A2 => n1983, B1 => n795, B2 => n1977, 
                           ZN => n1475);
   U209 : OAI22_X1 port map( A1 => n903, A2 => n1983, B1 => n797, B2 => n1977, 
                           ZN => n1474);
   U210 : OAI22_X1 port map( A1 => n904, A2 => n1983, B1 => n799, B2 => n1976, 
                           ZN => n1473);
   U211 : OAI22_X1 port map( A1 => n905, A2 => n1982, B1 => n801, B2 => n1976, 
                           ZN => n1472);
   U212 : OAI22_X1 port map( A1 => n906, A2 => n1982, B1 => n803, B2 => n1976, 
                           ZN => n1471);
   U213 : OAI22_X1 port map( A1 => n907, A2 => n1982, B1 => n805, B2 => n1976, 
                           ZN => n1470);
   U214 : OAI22_X1 port map( A1 => n908, A2 => n1982, B1 => n807, B2 => n1976, 
                           ZN => n1469);
   U215 : OAI22_X1 port map( A1 => n909, A2 => n1982, B1 => n809, B2 => n1976, 
                           ZN => n1468);
   U216 : OAI22_X1 port map( A1 => n910, A2 => n1982, B1 => n811, B2 => n1976, 
                           ZN => n1467);
   U217 : OAI22_X1 port map( A1 => n911, A2 => n1982, B1 => n813, B2 => n1976, 
                           ZN => n1466);
   U218 : OAI22_X1 port map( A1 => n912, A2 => n1982, B1 => n815, B2 => n1976, 
                           ZN => n1465);
   U219 : OAI22_X1 port map( A1 => n913, A2 => n1982, B1 => n817, B2 => n1976, 
                           ZN => n1464);
   U220 : OAI22_X1 port map( A1 => n914, A2 => n1982, B1 => n819, B2 => n1976, 
                           ZN => n1463);
   U221 : OAI22_X1 port map( A1 => n915, A2 => n1982, B1 => n821, B2 => n1976, 
                           ZN => n1462);
   U222 : OAI22_X1 port map( A1 => n916, A2 => n1982, B1 => n823, B2 => n1975, 
                           ZN => n1461);
   U223 : OAI22_X1 port map( A1 => n917, A2 => n1981, B1 => n825, B2 => n1975, 
                           ZN => n1460);
   U224 : OAI22_X1 port map( A1 => n918, A2 => n1981, B1 => n827, B2 => n1975, 
                           ZN => n1459);
   U225 : OAI22_X1 port map( A1 => n919, A2 => n1981, B1 => n829, B2 => n1975, 
                           ZN => n1458);
   U226 : OAI22_X1 port map( A1 => n920, A2 => n1981, B1 => n831, B2 => n1975, 
                           ZN => n1457);
   U227 : OAI22_X1 port map( A1 => n921, A2 => n1981, B1 => n833, B2 => n1975, 
                           ZN => n1456);
   U228 : OAI22_X1 port map( A1 => n922, A2 => n1981, B1 => n835, B2 => n1975, 
                           ZN => n1455);
   U229 : OAI22_X1 port map( A1 => n923, A2 => n1981, B1 => n837, B2 => n1975, 
                           ZN => n1454);
   U230 : OAI22_X1 port map( A1 => n924, A2 => n1981, B1 => n839, B2 => n1975, 
                           ZN => n1453);
   U231 : OAI22_X1 port map( A1 => n925, A2 => n1981, B1 => n841, B2 => n1975, 
                           ZN => n1452);
   U232 : OAI22_X1 port map( A1 => n926, A2 => n1981, B1 => n843, B2 => n1975, 
                           ZN => n1451);
   U233 : OAI22_X1 port map( A1 => n927, A2 => n1981, B1 => n845, B2 => n1975, 
                           ZN => n1450);
   U234 : OAI22_X1 port map( A1 => n1204, A2 => n1981, B1 => n847, B2 => n1974,
                           ZN => n1449);
   U235 : OAI22_X1 port map( A1 => n1202, A2 => n1980, B1 => n849, B2 => n1974,
                           ZN => n1448);
   U236 : OAI22_X1 port map( A1 => n1200, A2 => n1980, B1 => n851, B2 => n1974,
                           ZN => n1447);
   U237 : OAI22_X1 port map( A1 => n928, A2 => n1980, B1 => n853, B2 => n1974, 
                           ZN => n1446);
   U238 : OAI22_X1 port map( A1 => n929, A2 => n1980, B1 => n855, B2 => n1974, 
                           ZN => n1445);
   U239 : OAI22_X1 port map( A1 => n930, A2 => n1980, B1 => n857, B2 => n1974, 
                           ZN => n1444);
   U240 : OAI22_X1 port map( A1 => n931, A2 => n1980, B1 => n859, B2 => n1974, 
                           ZN => n1443);
   U241 : OAI22_X1 port map( A1 => n932, A2 => n1980, B1 => n861, B2 => n1974, 
                           ZN => n1442);
   U242 : OAI22_X1 port map( A1 => n933, A2 => n1980, B1 => n863, B2 => n1974, 
                           ZN => n1441);
   U243 : OAI22_X1 port map( A1 => n934, A2 => n1980, B1 => n865, B2 => n1974, 
                           ZN => n1440);
   U244 : OAI22_X1 port map( A1 => n935, A2 => n1980, B1 => n867, B2 => n1974, 
                           ZN => n1439);
   U245 : OAI22_X1 port map( A1 => n415, A2 => n1980, B1 => n871, B2 => n1974, 
                           ZN => n1438);
   U246 : OAI22_X1 port map( A1 => n1817, A2 => n1973, B1 => n751, B2 => n1966,
                           ZN => n1433);
   U247 : OAI22_X1 port map( A1 => n1816, A2 => n1972, B1 => n753, B2 => n1966,
                           ZN => n1432);
   U248 : OAI22_X1 port map( A1 => n1815, A2 => n1972, B1 => n755, B2 => n1966,
                           ZN => n1431);
   U249 : OAI22_X1 port map( A1 => n1814, A2 => n1972, B1 => n757, B2 => n1966,
                           ZN => n1430);
   U250 : OAI22_X1 port map( A1 => n1813, A2 => n1972, B1 => n759, B2 => n1966,
                           ZN => n1429);
   U251 : OAI22_X1 port map( A1 => n1812, A2 => n1972, B1 => n761, B2 => n1966,
                           ZN => n1428);
   U252 : OAI22_X1 port map( A1 => n1811, A2 => n1972, B1 => n763, B2 => n1966,
                           ZN => n1427);
   U253 : OAI22_X1 port map( A1 => n1810, A2 => n1972, B1 => n765, B2 => n1966,
                           ZN => n1426);
   U254 : OAI22_X1 port map( A1 => n1809, A2 => n1972, B1 => n767, B2 => n1966,
                           ZN => n1425);
   U255 : OAI22_X1 port map( A1 => n1808, A2 => n1972, B1 => n769, B2 => n1966,
                           ZN => n1424);
   U256 : OAI22_X1 port map( A1 => n1807, A2 => n1972, B1 => n771, B2 => n1966,
                           ZN => n1423);
   U257 : OAI22_X1 port map( A1 => n1806, A2 => n1972, B1 => n773, B2 => n1966,
                           ZN => n1422);
   U258 : OAI22_X1 port map( A1 => n1805, A2 => n1972, B1 => n775, B2 => n1965,
                           ZN => n1421);
   U259 : OAI22_X1 port map( A1 => n1804, A2 => n1971, B1 => n777, B2 => n1965,
                           ZN => n1420);
   U260 : OAI22_X1 port map( A1 => n1803, A2 => n1971, B1 => n779, B2 => n1965,
                           ZN => n1419);
   U261 : OAI22_X1 port map( A1 => n1802, A2 => n1971, B1 => n781, B2 => n1965,
                           ZN => n1418);
   U262 : OAI22_X1 port map( A1 => n1801, A2 => n1971, B1 => n783, B2 => n1965,
                           ZN => n1417);
   U263 : OAI22_X1 port map( A1 => n1800, A2 => n1971, B1 => n785, B2 => n1965,
                           ZN => n1416);
   U264 : OAI22_X1 port map( A1 => n1799, A2 => n1971, B1 => n787, B2 => n1965,
                           ZN => n1415);
   U265 : OAI22_X1 port map( A1 => n1798, A2 => n1971, B1 => n789, B2 => n1965,
                           ZN => n1414);
   U266 : OAI22_X1 port map( A1 => n1797, A2 => n1971, B1 => n791, B2 => n1965,
                           ZN => n1413);
   U267 : OAI22_X1 port map( A1 => n1796, A2 => n1971, B1 => n793, B2 => n1965,
                           ZN => n1412);
   U268 : OAI22_X1 port map( A1 => n1795, A2 => n1971, B1 => n795, B2 => n1965,
                           ZN => n1411);
   U269 : OAI22_X1 port map( A1 => n1794, A2 => n1971, B1 => n797, B2 => n1965,
                           ZN => n1410);
   U270 : OAI22_X1 port map( A1 => n1793, A2 => n1971, B1 => n799, B2 => n1964,
                           ZN => n1409);
   U271 : OAI22_X1 port map( A1 => n940, A2 => n1970, B1 => n801, B2 => n1964, 
                           ZN => n1408);
   U272 : OAI22_X1 port map( A1 => n941, A2 => n1970, B1 => n803, B2 => n1964, 
                           ZN => n1407);
   U273 : OAI22_X1 port map( A1 => n942, A2 => n1970, B1 => n805, B2 => n1964, 
                           ZN => n1406);
   U274 : OAI22_X1 port map( A1 => n943, A2 => n1970, B1 => n807, B2 => n1964, 
                           ZN => n1405);
   U275 : OAI22_X1 port map( A1 => n944, A2 => n1970, B1 => n809, B2 => n1964, 
                           ZN => n1404);
   U276 : OAI22_X1 port map( A1 => n945, A2 => n1970, B1 => n811, B2 => n1964, 
                           ZN => n1403);
   U277 : OAI22_X1 port map( A1 => n946, A2 => n1970, B1 => n813, B2 => n1964, 
                           ZN => n1402);
   U278 : OAI22_X1 port map( A1 => n947, A2 => n1970, B1 => n815, B2 => n1964, 
                           ZN => n1401);
   U279 : OAI22_X1 port map( A1 => n948, A2 => n1970, B1 => n817, B2 => n1964, 
                           ZN => n1400);
   U280 : OAI22_X1 port map( A1 => n949, A2 => n1970, B1 => n819, B2 => n1964, 
                           ZN => n1399);
   U281 : OAI22_X1 port map( A1 => n950, A2 => n1970, B1 => n821, B2 => n1964, 
                           ZN => n1398);
   U282 : OAI22_X1 port map( A1 => n951, A2 => n1970, B1 => n823, B2 => n1963, 
                           ZN => n1397);
   U283 : OAI22_X1 port map( A1 => n952, A2 => n1969, B1 => n825, B2 => n1963, 
                           ZN => n1396);
   U284 : OAI22_X1 port map( A1 => n953, A2 => n1969, B1 => n827, B2 => n1963, 
                           ZN => n1395);
   U285 : OAI22_X1 port map( A1 => n954, A2 => n1969, B1 => n829, B2 => n1963, 
                           ZN => n1394);
   U286 : OAI22_X1 port map( A1 => n955, A2 => n1969, B1 => n831, B2 => n1963, 
                           ZN => n1393);
   U287 : OAI22_X1 port map( A1 => n956, A2 => n1969, B1 => n833, B2 => n1963, 
                           ZN => n1392);
   U288 : OAI22_X1 port map( A1 => n957, A2 => n1969, B1 => n835, B2 => n1963, 
                           ZN => n1391);
   U289 : OAI22_X1 port map( A1 => n958, A2 => n1969, B1 => n837, B2 => n1963, 
                           ZN => n1390);
   U290 : OAI22_X1 port map( A1 => n959, A2 => n1969, B1 => n839, B2 => n1963, 
                           ZN => n1389);
   U291 : OAI22_X1 port map( A1 => n960, A2 => n1969, B1 => n841, B2 => n1963, 
                           ZN => n1388);
   U292 : OAI22_X1 port map( A1 => n961, A2 => n1969, B1 => n843, B2 => n1963, 
                           ZN => n1387);
   U293 : OAI22_X1 port map( A1 => n962, A2 => n1969, B1 => n845, B2 => n1963, 
                           ZN => n1386);
   U294 : OAI22_X1 port map( A1 => n963, A2 => n1969, B1 => n847, B2 => n1962, 
                           ZN => n1385);
   U295 : OAI22_X1 port map( A1 => n964, A2 => n1968, B1 => n849, B2 => n1962, 
                           ZN => n1384);
   U296 : OAI22_X1 port map( A1 => n965, A2 => n1968, B1 => n851, B2 => n1962, 
                           ZN => n1383);
   U297 : OAI22_X1 port map( A1 => n966, A2 => n1968, B1 => n853, B2 => n1962, 
                           ZN => n1382);
   U298 : OAI22_X1 port map( A1 => n967, A2 => n1968, B1 => n855, B2 => n1962, 
                           ZN => n1381);
   U299 : OAI22_X1 port map( A1 => n968, A2 => n1968, B1 => n857, B2 => n1962, 
                           ZN => n1380);
   U300 : OAI22_X1 port map( A1 => n969, A2 => n1968, B1 => n859, B2 => n1962, 
                           ZN => n1379);
   U301 : OAI22_X1 port map( A1 => n970, A2 => n1968, B1 => n861, B2 => n1962, 
                           ZN => n1378);
   U302 : OAI22_X1 port map( A1 => n971, A2 => n1968, B1 => n863, B2 => n1962, 
                           ZN => n1377);
   U303 : OAI22_X1 port map( A1 => n972, A2 => n1968, B1 => n865, B2 => n1962, 
                           ZN => n1376);
   U304 : OAI22_X1 port map( A1 => n973, A2 => n1968, B1 => n867, B2 => n1962, 
                           ZN => n1375);
   U305 : OAI22_X1 port map( A1 => n974, A2 => n1968, B1 => n871, B2 => n1962, 
                           ZN => n1374);
   U306 : OAI22_X1 port map( A1 => n983, A2 => n1961, B1 => n751, B2 => n1954, 
                           ZN => n1369);
   U307 : OAI22_X1 port map( A1 => n984, A2 => n1960, B1 => n753, B2 => n1954, 
                           ZN => n1368);
   U308 : OAI22_X1 port map( A1 => n985, A2 => n1960, B1 => n755, B2 => n1954, 
                           ZN => n1367);
   U309 : OAI22_X1 port map( A1 => n986, A2 => n1960, B1 => n757, B2 => n1954, 
                           ZN => n1366);
   U310 : OAI22_X1 port map( A1 => n987, A2 => n1960, B1 => n759, B2 => n1954, 
                           ZN => n1365);
   U311 : OAI22_X1 port map( A1 => n988, A2 => n1960, B1 => n761, B2 => n1954, 
                           ZN => n1364);
   U312 : OAI22_X1 port map( A1 => n989, A2 => n1960, B1 => n763, B2 => n1954, 
                           ZN => n1363);
   U313 : OAI22_X1 port map( A1 => n990, A2 => n1960, B1 => n765, B2 => n1954, 
                           ZN => n1362);
   U314 : OAI22_X1 port map( A1 => n991, A2 => n1960, B1 => n767, B2 => n1954, 
                           ZN => n1361);
   U315 : OAI22_X1 port map( A1 => n992, A2 => n1960, B1 => n769, B2 => n1954, 
                           ZN => n1360);
   U316 : OAI22_X1 port map( A1 => n993, A2 => n1960, B1 => n771, B2 => n1954, 
                           ZN => n1359);
   U317 : OAI22_X1 port map( A1 => n994, A2 => n1960, B1 => n773, B2 => n1954, 
                           ZN => n1358);
   U318 : OAI22_X1 port map( A1 => n995, A2 => n1960, B1 => n775, B2 => n1953, 
                           ZN => n1357);
   U319 : OAI22_X1 port map( A1 => n996, A2 => n1959, B1 => n777, B2 => n1953, 
                           ZN => n1356);
   U320 : OAI22_X1 port map( A1 => n997, A2 => n1959, B1 => n779, B2 => n1953, 
                           ZN => n1355);
   U321 : OAI22_X1 port map( A1 => n1738, A2 => n1959, B1 => n781, B2 => n1953,
                           ZN => n1354);
   U322 : OAI22_X1 port map( A1 => n1737, A2 => n1959, B1 => n783, B2 => n1953,
                           ZN => n1353);
   U323 : OAI22_X1 port map( A1 => n1736, A2 => n1959, B1 => n785, B2 => n1953,
                           ZN => n1352);
   U324 : OAI22_X1 port map( A1 => n1735, A2 => n1959, B1 => n787, B2 => n1953,
                           ZN => n1351);
   U325 : OAI22_X1 port map( A1 => n1734, A2 => n1959, B1 => n789, B2 => n1953,
                           ZN => n1350);
   U326 : OAI22_X1 port map( A1 => n1733, A2 => n1959, B1 => n791, B2 => n1953,
                           ZN => n1349);
   U327 : OAI22_X1 port map( A1 => n1732, A2 => n1959, B1 => n793, B2 => n1953,
                           ZN => n1348);
   U328 : OAI22_X1 port map( A1 => n1731, A2 => n1959, B1 => n795, B2 => n1953,
                           ZN => n1347);
   U329 : OAI22_X1 port map( A1 => n1730, A2 => n1959, B1 => n797, B2 => n1953,
                           ZN => n1346);
   U330 : OAI22_X1 port map( A1 => n1729, A2 => n1959, B1 => n799, B2 => n1952,
                           ZN => n1345);
   U331 : OAI22_X1 port map( A1 => n1728, A2 => n1958, B1 => n801, B2 => n1952,
                           ZN => n1344);
   U332 : OAI22_X1 port map( A1 => n1727, A2 => n1958, B1 => n803, B2 => n1952,
                           ZN => n1343);
   U333 : OAI22_X1 port map( A1 => n1726, A2 => n1958, B1 => n805, B2 => n1952,
                           ZN => n1342);
   U334 : OAI22_X1 port map( A1 => n1725, A2 => n1958, B1 => n807, B2 => n1952,
                           ZN => n1341);
   U335 : OAI22_X1 port map( A1 => n1724, A2 => n1958, B1 => n809, B2 => n1952,
                           ZN => n1340);
   U336 : OAI22_X1 port map( A1 => n1723, A2 => n1958, B1 => n811, B2 => n1952,
                           ZN => n1339);
   U337 : OAI22_X1 port map( A1 => n1722, A2 => n1958, B1 => n813, B2 => n1952,
                           ZN => n1338);
   U338 : OAI22_X1 port map( A1 => n1721, A2 => n1958, B1 => n815, B2 => n1952,
                           ZN => n1337);
   U339 : OAI22_X1 port map( A1 => n1720, A2 => n1958, B1 => n817, B2 => n1952,
                           ZN => n1336);
   U340 : OAI22_X1 port map( A1 => n1719, A2 => n1958, B1 => n819, B2 => n1952,
                           ZN => n1335);
   U341 : OAI22_X1 port map( A1 => n1718, A2 => n1958, B1 => n821, B2 => n1952,
                           ZN => n1334);
   U342 : OAI22_X1 port map( A1 => n1717, A2 => n1958, B1 => n823, B2 => n1951,
                           ZN => n1333);
   U343 : OAI22_X1 port map( A1 => n1716, A2 => n1957, B1 => n825, B2 => n1951,
                           ZN => n1332);
   U344 : OAI22_X1 port map( A1 => n1715, A2 => n1957, B1 => n827, B2 => n1951,
                           ZN => n1331);
   U345 : OAI22_X1 port map( A1 => n1714, A2 => n1957, B1 => n829, B2 => n1951,
                           ZN => n1330);
   U346 : OAI22_X1 port map( A1 => n1713, A2 => n1957, B1 => n831, B2 => n1951,
                           ZN => n1329);
   U347 : OAI22_X1 port map( A1 => n1712, A2 => n1957, B1 => n833, B2 => n1951,
                           ZN => n1328);
   U348 : OAI22_X1 port map( A1 => n1711, A2 => n1957, B1 => n835, B2 => n1951,
                           ZN => n1327);
   U349 : OAI22_X1 port map( A1 => n1710, A2 => n1957, B1 => n837, B2 => n1951,
                           ZN => n1326);
   U350 : OAI22_X1 port map( A1 => n1709, A2 => n1957, B1 => n839, B2 => n1951,
                           ZN => n1325);
   U351 : OAI22_X1 port map( A1 => n1708, A2 => n1957, B1 => n841, B2 => n1951,
                           ZN => n1324);
   U352 : OAI22_X1 port map( A1 => n1707, A2 => n1957, B1 => n843, B2 => n1951,
                           ZN => n1323);
   U353 : OAI22_X1 port map( A1 => n1706, A2 => n1957, B1 => n845, B2 => n1951,
                           ZN => n1322);
   U354 : OAI22_X1 port map( A1 => n1705, A2 => n1957, B1 => n847, B2 => n1950,
                           ZN => n1321);
   U355 : OAI22_X1 port map( A1 => n1704, A2 => n1956, B1 => n849, B2 => n1950,
                           ZN => n1320);
   U356 : OAI22_X1 port map( A1 => n1703, A2 => n1956, B1 => n851, B2 => n1950,
                           ZN => n1319);
   U357 : OAI22_X1 port map( A1 => n1702, A2 => n1956, B1 => n853, B2 => n1950,
                           ZN => n1318);
   U358 : OAI22_X1 port map( A1 => n1701, A2 => n1956, B1 => n855, B2 => n1950,
                           ZN => n1317);
   U359 : OAI22_X1 port map( A1 => n1700, A2 => n1956, B1 => n857, B2 => n1950,
                           ZN => n1316);
   U360 : OAI22_X1 port map( A1 => n1699, A2 => n1956, B1 => n859, B2 => n1950,
                           ZN => n1315);
   U361 : OAI22_X1 port map( A1 => n1698, A2 => n1956, B1 => n861, B2 => n1950,
                           ZN => n1314);
   U362 : OAI22_X1 port map( A1 => n1697, A2 => n1956, B1 => n863, B2 => n1950,
                           ZN => n1313);
   U363 : OAI22_X1 port map( A1 => n1696, A2 => n1956, B1 => n865, B2 => n1950,
                           ZN => n1312);
   U364 : OAI22_X1 port map( A1 => n1695, A2 => n1956, B1 => n867, B2 => n1950,
                           ZN => n1311);
   U365 : OAI22_X1 port map( A1 => n1694, A2 => n1956, B1 => n871, B2 => n1950,
                           ZN => n1310);
   U366 : OAI221_X1 port map( B1 => n2055, B2 => n562, C1 => n1937, C2 => n2046
                           , A => n563, ZN => n1681);
   U367 : AOI222_X1 port map( A1 => n52, A2 => n2039, B1 => n180, B2 => n2035, 
                           C1 => n2032, C2 => n564, ZN => n563);
   U368 : OAI221_X1 port map( B1 => n2055, B2 => n565, C1 => n1936, C2 => n2046
                           , A => n566, ZN => n1680);
   U369 : AOI222_X1 port map( A1 => n51, A2 => n2040, B1 => n179, B2 => n2035, 
                           C1 => n2032, C2 => n567, ZN => n566);
   U370 : OAI221_X1 port map( B1 => n2055, B2 => n568, C1 => n1935, C2 => n2046
                           , A => n569, ZN => n1679);
   U371 : AOI222_X1 port map( A1 => n50, A2 => n2040, B1 => n178, B2 => n2035, 
                           C1 => n2032, C2 => n570, ZN => n569);
   U372 : OAI221_X1 port map( B1 => n2055, B2 => n571, C1 => n1934, C2 => n2047
                           , A => n572, ZN => n1678);
   U373 : AOI222_X1 port map( A1 => n49, A2 => n2040, B1 => n177, B2 => n2035, 
                           C1 => n2031, C2 => n573, ZN => n572);
   U374 : OAI221_X1 port map( B1 => n2054, B2 => n574, C1 => n1933, C2 => n2046
                           , A => n575, ZN => n1677);
   U375 : AOI222_X1 port map( A1 => n48, A2 => n2040, B1 => n176, B2 => n2035, 
                           C1 => n2031, C2 => n576, ZN => n575);
   U376 : OAI221_X1 port map( B1 => n2054, B2 => n577, C1 => n1932, C2 => n2046
                           , A => n578, ZN => n1676);
   U377 : AOI222_X1 port map( A1 => n47, A2 => n2040, B1 => n175, B2 => n2035, 
                           C1 => n2031, C2 => n579, ZN => n578);
   U378 : OAI221_X1 port map( B1 => n2054, B2 => n580, C1 => n1931, C2 => n2046
                           , A => n581, ZN => n1675);
   U379 : AOI222_X1 port map( A1 => n46, A2 => n2040, B1 => n174, B2 => n2035, 
                           C1 => n2031, C2 => n582, ZN => n581);
   U380 : OAI221_X1 port map( B1 => n538, B2 => n2026, C1 => n1881, C2 => n2016
                           , A => n750, ZN => n1621);
   U381 : AOI222_X1 port map( A1 => n2014, A2 => n60, B1 => n2008, B2 => n188, 
                           C1 => n2002, C2 => n540, ZN => n750);
   U382 : OAI221_X1 port map( B1 => n541, B2 => n2026, C1 => n1880, C2 => n2016
                           , A => n752, ZN => n1619);
   U383 : AOI222_X1 port map( A1 => n2014, A2 => n59, B1 => n2008, B2 => n187, 
                           C1 => n2002, C2 => n543, ZN => n752);
   U384 : OAI221_X1 port map( B1 => n544, B2 => n2026, C1 => n1879, C2 => n2016
                           , A => n754, ZN => n1617);
   U385 : AOI222_X1 port map( A1 => n2014, A2 => n58, B1 => n2008, B2 => n186, 
                           C1 => n2002, C2 => n546, ZN => n754);
   U386 : OAI221_X1 port map( B1 => n547, B2 => n2026, C1 => n1878, C2 => n2016
                           , A => n756, ZN => n1615);
   U387 : AOI222_X1 port map( A1 => n2014, A2 => n57, B1 => n2008, B2 => n185, 
                           C1 => n2002, C2 => n549, ZN => n756);
   U388 : OAI221_X1 port map( B1 => n550, B2 => n2026, C1 => n1877, C2 => n2016
                           , A => n758, ZN => n1613);
   U389 : AOI222_X1 port map( A1 => n2014, A2 => n56, B1 => n2008, B2 => n184, 
                           C1 => n2002, C2 => n552, ZN => n758);
   U390 : OAI221_X1 port map( B1 => n553, B2 => n2026, C1 => n1876, C2 => n2016
                           , A => n760, ZN => n1611);
   U391 : AOI222_X1 port map( A1 => n2014, A2 => n55, B1 => n2008, B2 => n183, 
                           C1 => n2002, C2 => n555, ZN => n760);
   U392 : OAI221_X1 port map( B1 => n556, B2 => n2026, C1 => n1875, C2 => n2016
                           , A => n762, ZN => n1609);
   U393 : AOI222_X1 port map( A1 => n2014, A2 => n54, B1 => n2008, B2 => n182, 
                           C1 => n2002, C2 => n558, ZN => n762);
   U394 : OAI221_X1 port map( B1 => n559, B2 => n2026, C1 => n1874, C2 => n2016
                           , A => n764, ZN => n1607);
   U395 : AOI222_X1 port map( A1 => n2014, A2 => n53, B1 => n2008, B2 => n181, 
                           C1 => n2002, C2 => n561, ZN => n764);
   U396 : OAI221_X1 port map( B1 => n562, B2 => n2026, C1 => n1873, C2 => n2017
                           , A => n766, ZN => n1605);
   U397 : AOI222_X1 port map( A1 => n2014, A2 => n52, B1 => n2008, B2 => n180, 
                           C1 => n2002, C2 => n564, ZN => n766);
   U398 : OAI221_X1 port map( B1 => n565, B2 => n2026, C1 => n1872, C2 => n2017
                           , A => n768, ZN => n1603);
   U399 : AOI222_X1 port map( A1 => n2014, A2 => n51, B1 => n2008, B2 => n179, 
                           C1 => n2002, C2 => n567, ZN => n768);
   U400 : OAI221_X1 port map( B1 => n568, B2 => n2026, C1 => n1871, C2 => n2017
                           , A => n770, ZN => n1601);
   U401 : AOI222_X1 port map( A1 => n2014, A2 => n50, B1 => n2008, B2 => n178, 
                           C1 => n2002, C2 => n570, ZN => n770);
   U402 : OAI221_X1 port map( B1 => n571, B2 => n2026, C1 => n1870, C2 => n2018
                           , A => n772, ZN => n1599);
   U403 : AOI222_X1 port map( A1 => n2014, A2 => n49, B1 => n2008, B2 => n177, 
                           C1 => n2002, C2 => n573, ZN => n772);
   U404 : OAI221_X1 port map( B1 => n574, B2 => n2025, C1 => n1869, C2 => n2017
                           , A => n774, ZN => n1597);
   U405 : AOI222_X1 port map( A1 => n2013, A2 => n48, B1 => n2007, B2 => n176, 
                           C1 => n2001, C2 => n576, ZN => n774);
   U406 : OAI221_X1 port map( B1 => n577, B2 => n2025, C1 => n1868, C2 => n2017
                           , A => n776, ZN => n1595);
   U407 : AOI222_X1 port map( A1 => n2013, A2 => n47, B1 => n2007, B2 => n175, 
                           C1 => n2001, C2 => n579, ZN => n776);
   U408 : OAI221_X1 port map( B1 => n580, B2 => n2025, C1 => n1867, C2 => n2017
                           , A => n778, ZN => n1593);
   U409 : AOI222_X1 port map( A1 => n2013, A2 => n46, B1 => n2007, B2 => n174, 
                           C1 => n2001, C2 => n582, ZN => n778);
   U410 : OAI221_X1 port map( B1 => n2051, B2 => n716, C1 => n1890, C2 => n2050
                           , A => n717, ZN => n1634);
   U411 : AOI222_X1 port map( A1 => n5, A2 => n2043, B1 => n2038, B2 => n718, 
                           C1 => n69, C2 => n2028, ZN => n717);
   U412 : OAI221_X1 port map( B1 => n2051, B2 => n722, C1 => n1888, C2 => n2050
                           , A => n723, ZN => n1632);
   U413 : AOI222_X1 port map( A1 => n3, A2 => n2043, B1 => n2038, B2 => n724, 
                           C1 => n67, C2 => n2028, ZN => n723);
   U414 : OAI221_X1 port map( B1 => n2051, B2 => n725, C1 => n1887, C2 => n2050
                           , A => n726, ZN => n1631);
   U415 : AOI222_X1 port map( A1 => n2, A2 => n2043, B1 => n2038, B2 => n727, 
                           C1 => n66, C2 => n2028, ZN => n726);
   U416 : OAI221_X1 port map( B1 => n2051, B2 => n728, C1 => n1886, C2 => n2050
                           , A => n729, ZN => n1630);
   U417 : AOI222_X1 port map( A1 => n2044, A2 => n730, B1 => n2036, B2 => n731,
                           C1 => n65, C2 => n2028, ZN => n729);
   U418 : OAI221_X1 port map( B1 => n623, B2 => n2024, C1 => n1856, C2 => n2018
                           , A => n800, ZN => n1571);
   U419 : AOI222_X1 port map( A1 => n2012, A2 => n35, B1 => n2006, B2 => n625, 
                           C1 => n2000, C2 => n99, ZN => n800);
   U420 : OAI221_X1 port map( B1 => n626, B2 => n2024, C1 => n1855, C2 => n2018
                           , A => n802, ZN => n1569);
   U421 : AOI222_X1 port map( A1 => n2012, A2 => n34, B1 => n2006, B2 => n628, 
                           C1 => n2000, C2 => n98, ZN => n802);
   U422 : OAI221_X1 port map( B1 => n629, B2 => n2024, C1 => n1854, C2 => n2018
                           , A => n804, ZN => n1567);
   U423 : AOI222_X1 port map( A1 => n2012, A2 => n33, B1 => n2006, B2 => n631, 
                           C1 => n2000, C2 => n97, ZN => n804);
   U424 : OAI221_X1 port map( B1 => n632, B2 => n2024, C1 => n1853, C2 => n2018
                           , A => n806, ZN => n1565);
   U425 : AOI222_X1 port map( A1 => n2012, A2 => n32, B1 => n2006, B2 => n634, 
                           C1 => n2000, C2 => n96, ZN => n806);
   U426 : OAI221_X1 port map( B1 => n635, B2 => n2024, C1 => n1852, C2 => n2018
                           , A => n808, ZN => n1563);
   U427 : AOI222_X1 port map( A1 => n2012, A2 => n31, B1 => n2006, B2 => n637, 
                           C1 => n2000, C2 => n95, ZN => n808);
   U428 : OAI221_X1 port map( B1 => n638, B2 => n2024, C1 => n1851, C2 => n2018
                           , A => n810, ZN => n1561);
   U429 : AOI222_X1 port map( A1 => n2012, A2 => n30, B1 => n2006, B2 => n640, 
                           C1 => n2000, C2 => n94, ZN => n810);
   U430 : OAI221_X1 port map( B1 => n641, B2 => n2024, C1 => n1850, C2 => n2018
                           , A => n812, ZN => n1559);
   U431 : AOI222_X1 port map( A1 => n2012, A2 => n29, B1 => n2006, B2 => n643, 
                           C1 => n2000, C2 => n93, ZN => n812);
   U432 : OAI221_X1 port map( B1 => n644, B2 => n2024, C1 => n1849, C2 => n2019
                           , A => n814, ZN => n1557);
   U433 : AOI222_X1 port map( A1 => n2012, A2 => n28, B1 => n2006, B2 => n646, 
                           C1 => n2000, C2 => n92, ZN => n814);
   U434 : OAI221_X1 port map( B1 => n647, B2 => n2024, C1 => n1848, C2 => n2019
                           , A => n816, ZN => n1555);
   U435 : AOI222_X1 port map( A1 => n2012, A2 => n27, B1 => n2006, B2 => n649, 
                           C1 => n2000, C2 => n91, ZN => n816);
   U436 : OAI221_X1 port map( B1 => n650, B2 => n2024, C1 => n1847, C2 => n2019
                           , A => n818, ZN => n1553);
   U437 : AOI222_X1 port map( A1 => n2012, A2 => n26, B1 => n2006, B2 => n652, 
                           C1 => n2000, C2 => n90, ZN => n818);
   U438 : OAI221_X1 port map( B1 => n653, B2 => n2024, C1 => n1846, C2 => n2019
                           , A => n820, ZN => n1551);
   U439 : AOI222_X1 port map( A1 => n2012, A2 => n25, B1 => n2006, B2 => n655, 
                           C1 => n2000, C2 => n89, ZN => n820);
   U440 : OAI221_X1 port map( B1 => n656, B2 => n2023, C1 => n1845, C2 => n2019
                           , A => n822, ZN => n1549);
   U441 : AOI222_X1 port map( A1 => n2011, A2 => n24, B1 => n2005, B2 => n658, 
                           C1 => n1999, C2 => n88, ZN => n822);
   U442 : OAI221_X1 port map( B1 => n659, B2 => n2023, C1 => n1844, C2 => n2019
                           , A => n824, ZN => n1547);
   U443 : AOI222_X1 port map( A1 => n2011, A2 => n23, B1 => n2005, B2 => n661, 
                           C1 => n1999, C2 => n87, ZN => n824);
   U444 : OAI221_X1 port map( B1 => n662, B2 => n2023, C1 => n1843, C2 => n2019
                           , A => n826, ZN => n1545);
   U445 : AOI222_X1 port map( A1 => n2011, A2 => n22, B1 => n2005, B2 => n664, 
                           C1 => n1999, C2 => n86, ZN => n826);
   U446 : OAI221_X1 port map( B1 => n665, B2 => n2023, C1 => n1842, C2 => n2019
                           , A => n828, ZN => n1543);
   U447 : AOI222_X1 port map( A1 => n2011, A2 => n21, B1 => n2005, B2 => n667, 
                           C1 => n1999, C2 => n85, ZN => n828);
   U448 : OAI221_X1 port map( B1 => n668, B2 => n2023, C1 => n1841, C2 => n2019
                           , A => n830, ZN => n1541);
   U449 : AOI222_X1 port map( A1 => n2011, A2 => n20, B1 => n2005, B2 => n670, 
                           C1 => n1999, C2 => n84, ZN => n830);
   U450 : OAI221_X1 port map( B1 => n671, B2 => n2023, C1 => n1840, C2 => n2019
                           , A => n832, ZN => n1539);
   U451 : AOI222_X1 port map( A1 => n2011, A2 => n19, B1 => n2005, B2 => n673, 
                           C1 => n1999, C2 => n83, ZN => n832);
   U452 : OAI221_X1 port map( B1 => n674, B2 => n2023, C1 => n1839, C2 => n2019
                           , A => n834, ZN => n1537);
   U453 : AOI222_X1 port map( A1 => n2011, A2 => n18, B1 => n2005, B2 => n676, 
                           C1 => n1999, C2 => n82, ZN => n834);
   U454 : OAI221_X1 port map( B1 => n677, B2 => n2023, C1 => n1838, C2 => n2019
                           , A => n836, ZN => n1535);
   U455 : AOI222_X1 port map( A1 => n2011, A2 => n17, B1 => n2005, B2 => n679, 
                           C1 => n1999, C2 => n81, ZN => n836);
   U456 : OAI221_X1 port map( B1 => n680, B2 => n2023, C1 => n1837, C2 => n2020
                           , A => n838, ZN => n1533);
   U457 : AOI222_X1 port map( A1 => n2011, A2 => n16, B1 => n2005, B2 => n682, 
                           C1 => n1999, C2 => n80, ZN => n838);
   U458 : OAI221_X1 port map( B1 => n683, B2 => n2023, C1 => n1836, C2 => n2020
                           , A => n840, ZN => n1531);
   U459 : AOI222_X1 port map( A1 => n2011, A2 => n15, B1 => n2005, B2 => n685, 
                           C1 => n1999, C2 => n79, ZN => n840);
   U460 : OAI221_X1 port map( B1 => n686, B2 => n2023, C1 => n1835, C2 => n2020
                           , A => n842, ZN => n1529);
   U461 : AOI222_X1 port map( A1 => n2011, A2 => n14, B1 => n2005, B2 => n688, 
                           C1 => n1999, C2 => n78, ZN => n842);
   U462 : OAI221_X1 port map( B1 => n689, B2 => n2023, C1 => n1834, C2 => n2020
                           , A => n844, ZN => n1527);
   U463 : AOI222_X1 port map( A1 => n2011, A2 => n13, B1 => n2005, B2 => n691, 
                           C1 => n1999, C2 => n77, ZN => n844);
   U464 : OAI221_X1 port map( B1 => n692, B2 => n2022, C1 => n1833, C2 => n2020
                           , A => n846, ZN => n1525);
   U465 : AOI222_X1 port map( A1 => n2010, A2 => n694, B1 => n2004, B2 => n695,
                           C1 => n1998, C2 => n76, ZN => n846);
   U466 : OAI221_X1 port map( B1 => n696, B2 => n2022, C1 => n1832, C2 => n2020
                           , A => n848, ZN => n1523);
   U467 : AOI222_X1 port map( A1 => n2010, A2 => n698, B1 => n2004, B2 => n699,
                           C1 => n1998, C2 => n75, ZN => n848);
   U468 : OAI221_X1 port map( B1 => n700, B2 => n2022, C1 => n1831, C2 => n2020
                           , A => n850, ZN => n1521);
   U469 : AOI222_X1 port map( A1 => n2010, A2 => n702, B1 => n2004, B2 => n703,
                           C1 => n1998, C2 => n74, ZN => n850);
   U470 : OAI221_X1 port map( B1 => n704, B2 => n2022, C1 => n1830, C2 => n2020
                           , A => n852, ZN => n1519);
   U471 : AOI222_X1 port map( A1 => n2010, A2 => n9, B1 => n2004, B2 => n706, 
                           C1 => n1998, C2 => n73, ZN => n852);
   U472 : OAI221_X1 port map( B1 => n707, B2 => n2022, C1 => n1829, C2 => n2020
                           , A => n854, ZN => n1517);
   U473 : AOI222_X1 port map( A1 => n2010, A2 => n8, B1 => n2004, B2 => n709, 
                           C1 => n1998, C2 => n72, ZN => n854);
   U474 : OAI221_X1 port map( B1 => n710, B2 => n2022, C1 => n1828, C2 => n2020
                           , A => n856, ZN => n1515);
   U475 : AOI222_X1 port map( A1 => n2010, A2 => n7, B1 => n2004, B2 => n712, 
                           C1 => n1998, C2 => n71, ZN => n856);
   U476 : OAI221_X1 port map( B1 => n713, B2 => n2022, C1 => n1827, C2 => n2020
                           , A => n858, ZN => n1513);
   U477 : AOI222_X1 port map( A1 => n2010, A2 => n6, B1 => n2004, B2 => n715, 
                           C1 => n1998, C2 => n70, ZN => n858);
   U478 : OAI221_X1 port map( B1 => n716, B2 => n2022, C1 => n1826, C2 => n2021
                           , A => n860, ZN => n1511);
   U479 : AOI222_X1 port map( A1 => n2010, A2 => n5, B1 => n2004, B2 => n718, 
                           C1 => n1998, C2 => n69, ZN => n860);
   U480 : OAI221_X1 port map( B1 => n719, B2 => n2022, C1 => n1825, C2 => n2020
                           , A => n862, ZN => n1509);
   U481 : AOI222_X1 port map( A1 => n2010, A2 => n4, B1 => n2004, B2 => n721, 
                           C1 => n1998, C2 => n68, ZN => n862);
   U482 : OAI221_X1 port map( B1 => n722, B2 => n2022, C1 => n1824, C2 => n2021
                           , A => n864, ZN => n1507);
   U483 : AOI222_X1 port map( A1 => n2010, A2 => n3, B1 => n2004, B2 => n724, 
                           C1 => n1998, C2 => n67, ZN => n864);
   U484 : OAI221_X1 port map( B1 => n725, B2 => n2022, C1 => n1823, C2 => n2021
                           , A => n866, ZN => n1505);
   U485 : AOI222_X1 port map( A1 => n2010, A2 => n2, B1 => n2004, B2 => n727, 
                           C1 => n1998, C2 => n66, ZN => n866);
   U486 : OAI221_X1 port map( B1 => n728, B2 => n2022, C1 => n1822, C2 => n2021
                           , A => n868, ZN => n1503);
   U487 : AOI222_X1 port map( A1 => n2010, A2 => n730, B1 => n2004, B2 => n731,
                           C1 => n1998, C2 => n65, ZN => n868);
   U488 : INV_X1 port map( A => RESET, ZN => n734);
   U489 : OAI221_X1 port map( B1 => n2056, B2 => n522, C1 => n1949, C2 => n2045
                           , A => n524, ZN => n1693);
   U490 : AOI222_X1 port map( A1 => n64, A2 => n2041, B1 => n192, B2 => n2034, 
                           C1 => n2033, C2 => n528, ZN => n524);
   U491 : OAI221_X1 port map( B1 => n2056, B2 => n529, C1 => n1948, C2 => n2045
                           , A => n530, ZN => n1692);
   U492 : AOI222_X1 port map( A1 => n63, A2 => n2039, B1 => n191, B2 => n2034, 
                           C1 => n2033, C2 => n531, ZN => n530);
   U493 : OAI221_X1 port map( B1 => n2056, B2 => n532, C1 => n1947, C2 => n2045
                           , A => n533, ZN => n1691);
   U494 : AOI222_X1 port map( A1 => n62, A2 => n2039, B1 => n190, B2 => n2034, 
                           C1 => n2032, C2 => n534, ZN => n533);
   U495 : OAI221_X1 port map( B1 => n2056, B2 => n535, C1 => n1946, C2 => n2045
                           , A => n536, ZN => n1690);
   U496 : AOI222_X1 port map( A1 => n61, A2 => n2039, B1 => n189, B2 => n2034, 
                           C1 => n2032, C2 => n537, ZN => n536);
   U497 : OAI221_X1 port map( B1 => n2053, B2 => n619, C1 => n1921, C2 => n2047
                           , A => n620, ZN => n1665);
   U498 : AOI222_X1 port map( A1 => n36, A2 => n2041, B1 => n2036, B2 => n621, 
                           C1 => n2030, C2 => n622, ZN => n620);
   U499 : OAI221_X1 port map( B1 => n2053, B2 => n623, C1 => n1920, C2 => n2047
                           , A => n624, ZN => n1664);
   U500 : AOI222_X1 port map( A1 => n35, A2 => n2041, B1 => n2036, B2 => n625, 
                           C1 => n99, C2 => n2030, ZN => n624);
   U501 : OAI221_X1 port map( B1 => n2053, B2 => n626, C1 => n1919, C2 => n2047
                           , A => n627, ZN => n1663);
   U502 : AOI222_X1 port map( A1 => n34, A2 => n2041, B1 => n2036, B2 => n628, 
                           C1 => n98, C2 => n2030, ZN => n627);
   U503 : OAI221_X1 port map( B1 => n2053, B2 => n629, C1 => n1918, C2 => n2047
                           , A => n630, ZN => n1662);
   U504 : AOI222_X1 port map( A1 => n33, A2 => n2041, B1 => n2036, B2 => n631, 
                           C1 => n97, C2 => n2030, ZN => n630);
   U505 : OAI221_X1 port map( B1 => n2053, B2 => n632, C1 => n1917, C2 => n2047
                           , A => n633, ZN => n1661);
   U506 : AOI222_X1 port map( A1 => n32, A2 => n2041, B1 => n2036, B2 => n634, 
                           C1 => n96, C2 => n2030, ZN => n633);
   U507 : OAI221_X1 port map( B1 => n2053, B2 => n635, C1 => n1916, C2 => n2047
                           , A => n636, ZN => n1660);
   U508 : AOI222_X1 port map( A1 => n31, A2 => n2041, B1 => n2036, B2 => n637, 
                           C1 => n95, C2 => n2030, ZN => n636);
   U509 : OAI221_X1 port map( B1 => n2053, B2 => n638, C1 => n1915, C2 => n2047
                           , A => n639, ZN => n1659);
   U510 : AOI222_X1 port map( A1 => n30, A2 => n2041, B1 => n2036, B2 => n640, 
                           C1 => n94, C2 => n2030, ZN => n639);
   U511 : OAI221_X1 port map( B1 => n2053, B2 => n641, C1 => n1914, C2 => n2047
                           , A => n642, ZN => n1658);
   U512 : AOI222_X1 port map( A1 => n29, A2 => n2041, B1 => n2036, B2 => n643, 
                           C1 => n93, C2 => n2030, ZN => n642);
   U513 : OAI221_X1 port map( B1 => n2053, B2 => n644, C1 => n1913, C2 => n2048
                           , A => n645, ZN => n1657);
   U514 : AOI222_X1 port map( A1 => n28, A2 => n2042, B1 => n2036, B2 => n646, 
                           C1 => n92, C2 => n2030, ZN => n645);
   U515 : OAI221_X1 port map( B1 => n2053, B2 => n647, C1 => n1912, C2 => n2048
                           , A => n648, ZN => n1656);
   U516 : AOI222_X1 port map( A1 => n27, A2 => n2042, B1 => n2037, B2 => n649, 
                           C1 => n91, C2 => n2030, ZN => n648);
   U517 : OAI221_X1 port map( B1 => n2053, B2 => n650, C1 => n1911, C2 => n2048
                           , A => n651, ZN => n1655);
   U518 : AOI222_X1 port map( A1 => n26, A2 => n2042, B1 => n2037, B2 => n652, 
                           C1 => n90, C2 => n2030, ZN => n651);
   U519 : OAI221_X1 port map( B1 => n2053, B2 => n653, C1 => n1910, C2 => n2048
                           , A => n654, ZN => n1654);
   U520 : AOI222_X1 port map( A1 => n25, A2 => n2042, B1 => n2037, B2 => n655, 
                           C1 => n89, C2 => n2030, ZN => n654);
   U521 : OAI221_X1 port map( B1 => n2052, B2 => n656, C1 => n1909, C2 => n2048
                           , A => n657, ZN => n1653);
   U522 : AOI222_X1 port map( A1 => n24, A2 => n2042, B1 => n2037, B2 => n658, 
                           C1 => n88, C2 => n2029, ZN => n657);
   U523 : OAI221_X1 port map( B1 => n2052, B2 => n659, C1 => n1908, C2 => n2048
                           , A => n660, ZN => n1652);
   U524 : AOI222_X1 port map( A1 => n23, A2 => n2042, B1 => n2037, B2 => n661, 
                           C1 => n87, C2 => n2029, ZN => n660);
   U525 : OAI221_X1 port map( B1 => n2052, B2 => n662, C1 => n1907, C2 => n2048
                           , A => n663, ZN => n1651);
   U526 : AOI222_X1 port map( A1 => n22, A2 => n2042, B1 => n2037, B2 => n664, 
                           C1 => n86, C2 => n2029, ZN => n663);
   U527 : OAI221_X1 port map( B1 => n2052, B2 => n665, C1 => n1906, C2 => n2048
                           , A => n666, ZN => n1650);
   U528 : AOI222_X1 port map( A1 => n21, A2 => n2042, B1 => n2037, B2 => n667, 
                           C1 => n85, C2 => n2029, ZN => n666);
   U529 : OAI221_X1 port map( B1 => n2052, B2 => n668, C1 => n1905, C2 => n2048
                           , A => n669, ZN => n1649);
   U530 : AOI222_X1 port map( A1 => n20, A2 => n2042, B1 => n2037, B2 => n670, 
                           C1 => n84, C2 => n2029, ZN => n669);
   U531 : OAI221_X1 port map( B1 => n2052, B2 => n671, C1 => n1904, C2 => n2048
                           , A => n672, ZN => n1648);
   U532 : AOI222_X1 port map( A1 => n19, A2 => n2042, B1 => n2037, B2 => n673, 
                           C1 => n83, C2 => n2029, ZN => n672);
   U533 : OAI221_X1 port map( B1 => n2052, B2 => n674, C1 => n1903, C2 => n2048
                           , A => n675, ZN => n1647);
   U534 : AOI222_X1 port map( A1 => n18, A2 => n2042, B1 => n2037, B2 => n676, 
                           C1 => n82, C2 => n2029, ZN => n675);
   U535 : OAI221_X1 port map( B1 => n2052, B2 => n677, C1 => n1902, C2 => n2048
                           , A => n678, ZN => n1646);
   U536 : AOI222_X1 port map( A1 => n17, A2 => n2042, B1 => n2037, B2 => n679, 
                           C1 => n81, C2 => n2029, ZN => n678);
   U537 : OAI221_X1 port map( B1 => n2052, B2 => n680, C1 => n1901, C2 => n2049
                           , A => n681, ZN => n1645);
   U538 : AOI222_X1 port map( A1 => n16, A2 => n2043, B1 => n2037, B2 => n682, 
                           C1 => n80, C2 => n2029, ZN => n681);
   U539 : OAI221_X1 port map( B1 => n2052, B2 => n683, C1 => n1900, C2 => n2049
                           , A => n684, ZN => n1644);
   U540 : AOI222_X1 port map( A1 => n15, A2 => n2043, B1 => n2037, B2 => n685, 
                           C1 => n79, C2 => n2029, ZN => n684);
   U541 : OAI221_X1 port map( B1 => n2052, B2 => n686, C1 => n1899, C2 => n2049
                           , A => n687, ZN => n1643);
   U542 : AOI222_X1 port map( A1 => n14, A2 => n2043, B1 => n2038, B2 => n688, 
                           C1 => n78, C2 => n2029, ZN => n687);
   U543 : OAI221_X1 port map( B1 => n2052, B2 => n689, C1 => n1898, C2 => n2049
                           , A => n690, ZN => n1642);
   U544 : AOI222_X1 port map( A1 => n13, A2 => n2043, B1 => n2038, B2 => n691, 
                           C1 => n77, C2 => n2029, ZN => n690);
   U545 : OAI221_X1 port map( B1 => n2051, B2 => n692, C1 => n1897, C2 => n2049
                           , A => n693, ZN => n1641);
   U546 : AOI222_X1 port map( A1 => n2044, A2 => n694, B1 => n2038, B2 => n695,
                           C1 => n76, C2 => n2028, ZN => n693);
   U547 : OAI221_X1 port map( B1 => n2051, B2 => n696, C1 => n1896, C2 => n2049
                           , A => n697, ZN => n1640);
   U548 : AOI222_X1 port map( A1 => n2044, A2 => n698, B1 => n2038, B2 => n699,
                           C1 => n75, C2 => n2028, ZN => n697);
   U549 : OAI221_X1 port map( B1 => n2051, B2 => n700, C1 => n1895, C2 => n2049
                           , A => n701, ZN => n1639);
   U550 : AOI222_X1 port map( A1 => n2044, A2 => n702, B1 => n2038, B2 => n703,
                           C1 => n74, C2 => n2028, ZN => n701);
   U551 : OAI221_X1 port map( B1 => n2051, B2 => n704, C1 => n1894, C2 => n2049
                           , A => n705, ZN => n1638);
   U552 : AOI222_X1 port map( A1 => n9, A2 => n2043, B1 => n2038, B2 => n706, 
                           C1 => n73, C2 => n2028, ZN => n705);
   U553 : OAI221_X1 port map( B1 => n2051, B2 => n707, C1 => n1893, C2 => n2049
                           , A => n708, ZN => n1637);
   U554 : AOI222_X1 port map( A1 => n8, A2 => n2043, B1 => n2038, B2 => n709, 
                           C1 => n72, C2 => n2028, ZN => n708);
   U555 : OAI221_X1 port map( B1 => n2051, B2 => n710, C1 => n1892, C2 => n2049
                           , A => n711, ZN => n1636);
   U556 : AOI222_X1 port map( A1 => n7, A2 => n2043, B1 => n2038, B2 => n712, 
                           C1 => n71, C2 => n2028, ZN => n711);
   U557 : OAI221_X1 port map( B1 => n2051, B2 => n713, C1 => n1891, C2 => n2049
                           , A => n714, ZN => n1635);
   U558 : AOI222_X1 port map( A1 => n6, A2 => n2043, B1 => n2038, B2 => n715, 
                           C1 => n70, C2 => n2028, ZN => n714);
   U559 : OAI221_X1 port map( B1 => n2051, B2 => n719, C1 => n1889, C2 => n2049
                           , A => n720, ZN => n1633);
   U560 : AOI222_X1 port map( A1 => n4, A2 => n2043, B1 => n2038, B2 => n721, 
                           C1 => n68, C2 => n2028, ZN => n720);
   U561 : OAI221_X1 port map( B1 => n522, B2 => n2027, C1 => n1885, C2 => n2016
                           , A => n737, ZN => n1629);
   U562 : AOI222_X1 port map( A1 => n2015, A2 => n64, B1 => n2009, B2 => n192, 
                           C1 => n2003, C2 => n528, ZN => n737);
   U563 : OAI221_X1 port map( B1 => n529, B2 => n2027, C1 => n1884, C2 => n2016
                           , A => n744, ZN => n1627);
   U564 : AOI222_X1 port map( A1 => n2015, A2 => n63, B1 => n2009, B2 => n191, 
                           C1 => n2003, C2 => n531, ZN => n744);
   U565 : OAI221_X1 port map( B1 => n532, B2 => n2027, C1 => n1883, C2 => n2016
                           , A => n746, ZN => n1625);
   U566 : AOI222_X1 port map( A1 => n2015, A2 => n62, B1 => n2009, B2 => n190, 
                           C1 => n2003, C2 => n534, ZN => n746);
   U567 : OAI221_X1 port map( B1 => n535, B2 => n2027, C1 => n1882, C2 => n2016
                           , A => n748, ZN => n1623);
   U568 : AOI222_X1 port map( A1 => n2015, A2 => n61, B1 => n2009, B2 => n189, 
                           C1 => n2003, C2 => n537, ZN => n748);
   U569 : OAI221_X1 port map( B1 => n583, B2 => n2025, C1 => n1866, C2 => n2017
                           , A => n780, ZN => n1591);
   U570 : AOI222_X1 port map( A1 => n2013, A2 => n45, B1 => n2007, B2 => n585, 
                           C1 => n2001, C2 => n586, ZN => n780);
   U571 : OAI221_X1 port map( B1 => n587, B2 => n2025, C1 => n1865, C2 => n2017
                           , A => n782, ZN => n1589);
   U572 : AOI222_X1 port map( A1 => n2013, A2 => n44, B1 => n2007, B2 => n589, 
                           C1 => n2001, C2 => n590, ZN => n782);
   U573 : OAI221_X1 port map( B1 => n591, B2 => n2025, C1 => n1864, C2 => n2017
                           , A => n784, ZN => n1587);
   U574 : AOI222_X1 port map( A1 => n2013, A2 => n43, B1 => n2007, B2 => n593, 
                           C1 => n2001, C2 => n594, ZN => n784);
   U575 : OAI221_X1 port map( B1 => n595, B2 => n2025, C1 => n1863, C2 => n2017
                           , A => n786, ZN => n1585);
   U576 : AOI222_X1 port map( A1 => n2013, A2 => n42, B1 => n2007, B2 => n597, 
                           C1 => n2001, C2 => n598, ZN => n786);
   U577 : OAI221_X1 port map( B1 => n599, B2 => n2025, C1 => n1862, C2 => n2017
                           , A => n788, ZN => n1583);
   U578 : AOI222_X1 port map( A1 => n2013, A2 => n41, B1 => n2007, B2 => n601, 
                           C1 => n2001, C2 => n602, ZN => n788);
   U579 : OAI221_X1 port map( B1 => n603, B2 => n2025, C1 => n1861, C2 => n2017
                           , A => n790, ZN => n1581);
   U580 : AOI222_X1 port map( A1 => n2013, A2 => n40, B1 => n2007, B2 => n605, 
                           C1 => n2001, C2 => n606, ZN => n790);
   U581 : OAI221_X1 port map( B1 => n607, B2 => n2025, C1 => n1860, C2 => n2018
                           , A => n792, ZN => n1579);
   U582 : AOI222_X1 port map( A1 => n2013, A2 => n39, B1 => n2007, B2 => n609, 
                           C1 => n2001, C2 => n610, ZN => n792);
   U583 : OAI221_X1 port map( B1 => n611, B2 => n2025, C1 => n1859, C2 => n2018
                           , A => n794, ZN => n1577);
   U584 : AOI222_X1 port map( A1 => n2013, A2 => n38, B1 => n2007, B2 => n613, 
                           C1 => n2001, C2 => n614, ZN => n794);
   U585 : OAI221_X1 port map( B1 => n615, B2 => n2025, C1 => n1858, C2 => n2018
                           , A => n796, ZN => n1575);
   U586 : AOI222_X1 port map( A1 => n2013, A2 => n37, B1 => n2007, B2 => n617, 
                           C1 => n2001, C2 => n618, ZN => n796);
   U587 : OAI221_X1 port map( B1 => n619, B2 => n2024, C1 => n1857, C2 => n2018
                           , A => n798, ZN => n1573);
   U588 : AOI222_X1 port map( A1 => n2012, A2 => n36, B1 => n2006, B2 => n621, 
                           C1 => n2000, C2 => n622, ZN => n798);
   U589 : OAI221_X1 port map( B1 => n2055, B2 => n538, C1 => n1945, C2 => n2045
                           , A => n539, ZN => n1689);
   U590 : AOI222_X1 port map( A1 => n60, A2 => n2039, B1 => n188, B2 => n2034, 
                           C1 => n2032, C2 => n540, ZN => n539);
   U591 : OAI221_X1 port map( B1 => n2055, B2 => n541, C1 => n1944, C2 => n2045
                           , A => n542, ZN => n1688);
   U592 : AOI222_X1 port map( A1 => n59, A2 => n2039, B1 => n187, B2 => n2034, 
                           C1 => n2032, C2 => n543, ZN => n542);
   U593 : OAI221_X1 port map( B1 => n2055, B2 => n544, C1 => n1943, C2 => n2045
                           , A => n545, ZN => n1687);
   U594 : AOI222_X1 port map( A1 => n58, A2 => n2039, B1 => n186, B2 => n2034, 
                           C1 => n2032, C2 => n546, ZN => n545);
   U595 : OAI221_X1 port map( B1 => n2055, B2 => n547, C1 => n1942, C2 => n2045
                           , A => n548, ZN => n1686);
   U596 : AOI222_X1 port map( A1 => n57, A2 => n2039, B1 => n185, B2 => n2034, 
                           C1 => n2032, C2 => n549, ZN => n548);
   U597 : OAI221_X1 port map( B1 => n2055, B2 => n550, C1 => n1941, C2 => n2045
                           , A => n551, ZN => n1685);
   U598 : AOI222_X1 port map( A1 => n56, A2 => n2039, B1 => n184, B2 => n2034, 
                           C1 => n2032, C2 => n552, ZN => n551);
   U599 : OAI221_X1 port map( B1 => n2055, B2 => n553, C1 => n1940, C2 => n2045
                           , A => n554, ZN => n1684);
   U600 : AOI222_X1 port map( A1 => n55, A2 => n2039, B1 => n183, B2 => n2034, 
                           C1 => n2032, C2 => n555, ZN => n554);
   U601 : OAI221_X1 port map( B1 => n2055, B2 => n556, C1 => n1939, C2 => n2045
                           , A => n557, ZN => n1683);
   U602 : AOI222_X1 port map( A1 => n54, A2 => n2039, B1 => n182, B2 => n2034, 
                           C1 => n2032, C2 => n558, ZN => n557);
   U603 : OAI221_X1 port map( B1 => n2055, B2 => n559, C1 => n1938, C2 => n2045
                           , A => n560, ZN => n1682);
   U604 : AOI222_X1 port map( A1 => n53, A2 => n2039, B1 => n181, B2 => n2034, 
                           C1 => n2032, C2 => n561, ZN => n560);
   U605 : OAI221_X1 port map( B1 => n2054, B2 => n583, C1 => n1930, C2 => n2046
                           , A => n584, ZN => n1674);
   U606 : AOI222_X1 port map( A1 => n45, A2 => n2040, B1 => n2035, B2 => n585, 
                           C1 => n2031, C2 => n586, ZN => n584);
   U607 : OAI221_X1 port map( B1 => n2054, B2 => n587, C1 => n1929, C2 => n2046
                           , A => n588, ZN => n1673);
   U608 : AOI222_X1 port map( A1 => n44, A2 => n2040, B1 => n2035, B2 => n589, 
                           C1 => n2031, C2 => n590, ZN => n588);
   U609 : OAI221_X1 port map( B1 => n2054, B2 => n591, C1 => n1928, C2 => n2046
                           , A => n592, ZN => n1672);
   U610 : AOI222_X1 port map( A1 => n43, A2 => n2040, B1 => n2035, B2 => n593, 
                           C1 => n2031, C2 => n594, ZN => n592);
   U611 : OAI221_X1 port map( B1 => n2054, B2 => n595, C1 => n1927, C2 => n2046
                           , A => n596, ZN => n1671);
   U612 : AOI222_X1 port map( A1 => n42, A2 => n2040, B1 => n2035, B2 => n597, 
                           C1 => n2031, C2 => n598, ZN => n596);
   U613 : OAI221_X1 port map( B1 => n2054, B2 => n599, C1 => n1926, C2 => n2046
                           , A => n600, ZN => n1670);
   U614 : AOI222_X1 port map( A1 => n41, A2 => n2040, B1 => n2035, B2 => n601, 
                           C1 => n2031, C2 => n602, ZN => n600);
   U615 : OAI221_X1 port map( B1 => n2054, B2 => n603, C1 => n1925, C2 => n2046
                           , A => n604, ZN => n1669);
   U616 : AOI222_X1 port map( A1 => n40, A2 => n2040, B1 => n2036, B2 => n605, 
                           C1 => n2031, C2 => n606, ZN => n604);
   U617 : OAI221_X1 port map( B1 => n2054, B2 => n607, C1 => n1924, C2 => n2047
                           , A => n608, ZN => n1668);
   U618 : AOI222_X1 port map( A1 => n39, A2 => n2041, B1 => n2036, B2 => n609, 
                           C1 => n2031, C2 => n610, ZN => n608);
   U619 : OAI221_X1 port map( B1 => n2054, B2 => n611, C1 => n1923, C2 => n2047
                           , A => n612, ZN => n1667);
   U620 : AOI222_X1 port map( A1 => n38, A2 => n2041, B1 => n2036, B2 => n613, 
                           C1 => n2031, C2 => n614, ZN => n612);
   U621 : OAI221_X1 port map( B1 => n2054, B2 => n615, C1 => n1922, C2 => n2047
                           , A => n616, ZN => n1666);
   U622 : AOI222_X1 port map( A1 => n37, A2 => n2041, B1 => n2036, B2 => n617, 
                           C1 => n2031, C2 => n618, ZN => n616);
   U623 : INV_X1 port map( A => DATAIN(0), ZN => n743);
   U624 : INV_X1 port map( A => DATAIN(1), ZN => n745);
   U625 : INV_X1 port map( A => DATAIN(2), ZN => n747);
   U626 : INV_X1 port map( A => DATAIN(3), ZN => n749);
   U627 : INV_X1 port map( A => DATAIN(4), ZN => n751);
   U628 : INV_X1 port map( A => DATAIN(5), ZN => n753);
   U629 : INV_X1 port map( A => DATAIN(6), ZN => n755);
   U630 : INV_X1 port map( A => DATAIN(7), ZN => n757);
   U631 : INV_X1 port map( A => DATAIN(8), ZN => n759);
   U632 : INV_X1 port map( A => DATAIN(9), ZN => n761);
   U633 : INV_X1 port map( A => DATAIN(10), ZN => n763);
   U634 : INV_X1 port map( A => DATAIN(11), ZN => n765);
   U635 : INV_X1 port map( A => DATAIN(12), ZN => n767);
   U636 : INV_X1 port map( A => DATAIN(13), ZN => n769);
   U637 : INV_X1 port map( A => DATAIN(14), ZN => n771);
   U638 : INV_X1 port map( A => DATAIN(15), ZN => n773);
   U639 : INV_X1 port map( A => DATAIN(16), ZN => n775);
   U640 : INV_X1 port map( A => DATAIN(17), ZN => n777);
   U641 : INV_X1 port map( A => DATAIN(18), ZN => n779);
   U642 : INV_X1 port map( A => DATAIN(19), ZN => n781);
   U643 : INV_X1 port map( A => DATAIN(20), ZN => n783);
   U644 : INV_X1 port map( A => DATAIN(21), ZN => n785);
   U645 : INV_X1 port map( A => DATAIN(22), ZN => n787);
   U646 : INV_X1 port map( A => DATAIN(23), ZN => n789);
   U647 : INV_X1 port map( A => DATAIN(24), ZN => n791);
   U648 : INV_X1 port map( A => DATAIN(25), ZN => n793);
   U649 : INV_X1 port map( A => DATAIN(26), ZN => n795);
   U650 : INV_X1 port map( A => DATAIN(27), ZN => n797);
   U651 : INV_X1 port map( A => DATAIN(28), ZN => n799);
   U652 : INV_X1 port map( A => DATAIN(29), ZN => n801);
   U653 : INV_X1 port map( A => DATAIN(30), ZN => n803);
   U654 : INV_X1 port map( A => DATAIN(31), ZN => n805);
   U655 : INV_X1 port map( A => DATAIN(32), ZN => n807);
   U656 : INV_X1 port map( A => DATAIN(33), ZN => n809);
   U657 : INV_X1 port map( A => DATAIN(34), ZN => n811);
   U658 : INV_X1 port map( A => DATAIN(35), ZN => n813);
   U659 : INV_X1 port map( A => DATAIN(36), ZN => n815);
   U660 : INV_X1 port map( A => DATAIN(37), ZN => n817);
   U661 : INV_X1 port map( A => DATAIN(38), ZN => n819);
   U662 : INV_X1 port map( A => DATAIN(39), ZN => n821);
   U663 : INV_X1 port map( A => DATAIN(40), ZN => n823);
   U664 : INV_X1 port map( A => DATAIN(41), ZN => n825);
   U665 : INV_X1 port map( A => DATAIN(42), ZN => n827);
   U666 : INV_X1 port map( A => DATAIN(43), ZN => n829);
   U667 : INV_X1 port map( A => DATAIN(44), ZN => n831);
   U668 : INV_X1 port map( A => DATAIN(45), ZN => n833);
   U669 : INV_X1 port map( A => DATAIN(46), ZN => n835);
   U670 : INV_X1 port map( A => DATAIN(47), ZN => n837);
   U671 : INV_X1 port map( A => DATAIN(48), ZN => n839);
   U672 : INV_X1 port map( A => DATAIN(49), ZN => n841);
   U673 : INV_X1 port map( A => DATAIN(50), ZN => n843);
   U674 : INV_X1 port map( A => DATAIN(51), ZN => n845);
   U675 : INV_X1 port map( A => DATAIN(52), ZN => n847);
   U676 : INV_X1 port map( A => DATAIN(53), ZN => n849);
   U677 : INV_X1 port map( A => DATAIN(54), ZN => n851);
   U678 : INV_X1 port map( A => DATAIN(55), ZN => n853);
   U679 : INV_X1 port map( A => DATAIN(56), ZN => n855);
   U680 : INV_X1 port map( A => DATAIN(57), ZN => n857);
   U681 : INV_X1 port map( A => DATAIN(58), ZN => n859);
   U682 : INV_X1 port map( A => DATAIN(59), ZN => n861);
   U683 : INV_X1 port map( A => DATAIN(60), ZN => n863);
   U684 : INV_X1 port map( A => DATAIN(61), ZN => n865);
   U685 : INV_X1 port map( A => DATAIN(62), ZN => n867);
   U686 : INV_X1 port map( A => DATAIN(63), ZN => n871);
   U687 : CLKBUF_X1 port map( A => n979, Z => n1955);
   U688 : CLKBUF_X1 port map( A => n978, Z => n1961);
   U689 : CLKBUF_X1 port map( A => n939, Z => n1967);
   U690 : CLKBUF_X1 port map( A => n938, Z => n1973);
   U691 : CLKBUF_X1 port map( A => n876, Z => n1979);
   U692 : CLKBUF_X1 port map( A => n875, Z => n1985);
   U693 : CLKBUF_X1 port map( A => n742, Z => n1991);
   U694 : CLKBUF_X1 port map( A => n741, Z => n1997);
   U695 : CLKBUF_X1 port map( A => n740, Z => n2003);
   U696 : CLKBUF_X1 port map( A => n739, Z => n2009);
   U697 : CLKBUF_X1 port map( A => n738, Z => n2015);
   U698 : CLKBUF_X1 port map( A => n736, Z => n2021);
   U699 : CLKBUF_X1 port map( A => n735, Z => n2027);
   U700 : CLKBUF_X1 port map( A => n527, Z => n2033);
   U701 : CLKBUF_X1 port map( A => n525, Z => n2044);
   U702 : CLKBUF_X1 port map( A => n523, Z => n2050);
   U703 : CLKBUF_X1 port map( A => n521, Z => n2056);
   U704 : INV_X1 port map( A => ADD_RD2(0), ZN => n2057);
   U705 : INV_X1 port map( A => ADD_RD2(1), ZN => n2058);
   U706 : INV_X1 port map( A => ADD_RD1(0), ZN => n2059);
   U707 : INV_X1 port map( A => ADD_RD1(1), ZN => n2060);
   U708 : INV_X1 port map( A => ADD_WR(0), ZN => n2061);
   U709 : INV_X1 port map( A => ADD_WR(1), ZN => n2062);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4.all;

entity register_file_reg_size64_file_size4_3 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_reg_size64_file_size4_3;

architecture SYN_BEHAVIORAL of register_file_reg_size64_file_size4_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n415, n1200, n1202, n1204, n1310, n1311, n1312, n1313, n1314, n1315
      , n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n871, n872, 
      n873, n875, n876, n936, n938, n939, n975, n978, n979, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176 : std_logic
      ;

begin
   
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => n174,
                           QN => n2028);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => n175,
                           QN => n2027);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => n176,
                           QN => n2026);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => n177,
                           QN => n2025);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => n178,
                           QN => n2024);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => n179,
                           QN => n2023);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => n180,
                           QN => n2022);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => n181,
                           QN => n2021);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => n182,
                           QN => n2020);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => n183, 
                           QN => n2019);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => n184, 
                           QN => n2018);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => n185, 
                           QN => n2017);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => n186, 
                           QN => n2016);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => n187, 
                           QN => n2015);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => n188, 
                           QN => n2014);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => n189, 
                           QN => n2013);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => n190, 
                           QN => n2012);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => n191, 
                           QN => n2011);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => n192, 
                           QN => n2010);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => n65, 
                           QN => n2063);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => n66, 
                           QN => n2062);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n67, 
                           QN => n2061);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => n68, 
                           QN => n2060);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => n69, 
                           QN => n2059);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => n70, 
                           QN => n2058);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => n71, 
                           QN => n2057);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => n72, 
                           QN => n2056);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => n73, 
                           QN => n2055);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => n74, 
                           QN => n2054);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => n75, 
                           QN => n2053);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => n76, 
                           QN => n2052);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => n77, 
                           QN => n2051);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => n78, 
                           QN => n2050);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => n79, 
                           QN => n2049);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => n80, 
                           QN => n2048);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => n81, 
                           QN => n2047);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => n82, 
                           QN => n2046);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => n83, 
                           QN => n2045);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => n84, 
                           QN => n2044);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => n85, 
                           QN => n2043);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => n86, 
                           QN => n2042);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => n87, 
                           QN => n2041);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => n88, 
                           QN => n2040);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => n89, 
                           QN => n2039);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => n90, 
                           QN => n2038);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => n91, 
                           QN => n2037);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => n92, 
                           QN => n2036);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => n93, 
                           QN => n2035);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => n94, 
                           QN => n2034);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => n95, 
                           QN => n2033);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => n96, 
                           QN => n2032);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => n97, 
                           QN => n2031);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => n98, 
                           QN => n2030);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => n99, 
                           QN => n2029);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => n2, 
                           QN => n2009);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => n3, 
                           QN => n2008);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => n4, 
                           QN => n2007);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => n5, 
                           QN => n2006);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => n6, 
                           QN => n2005);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => n7, 
                           QN => n2004);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => n8, 
                           QN => n2003);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => n9, 
                           QN => n2002);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => n13, 
                           QN => n2001);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => n14, 
                           QN => n2000);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => n15, 
                           QN => n1999);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => n16, 
                           QN => n1998);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => n17, 
                           QN => n1997);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => n18, 
                           QN => n1996);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => n19, 
                           QN => n1995);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => n20, 
                           QN => n1994);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => n21, 
                           QN => n1993);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => n22, 
                           QN => n1992);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => n23, 
                           QN => n1991);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => n24, 
                           QN => n1990);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => n25, 
                           QN => n1989);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => n26, 
                           QN => n1988);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n27, 
                           QN => n1987);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => n28, 
                           QN => n1986);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n29, 
                           QN => n1985);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => n30, 
                           QN => n1984);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n31, 
                           QN => n1983);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => n32, 
                           QN => n1982);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n33, 
                           QN => n1981);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => n34, 
                           QN => n1980);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n35, 
                           QN => n1979);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => n36, 
                           QN => n1978);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => n37, 
                           QN => n1977);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => n38, 
                           QN => n1976);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => n39, 
                           QN => n1975);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => n40, 
                           QN => n1974);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => n41, 
                           QN => n1973);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => n42, 
                           QN => n1972);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => n43, 
                           QN => n1971);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => n44, 
                           QN => n1970);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => n45, 
                           QN => n1969);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => n46, 
                           QN => n1968);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => n47, 
                           QN => n1967);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => n48, 
                           QN => n1966);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => n49, 
                           QN => n1965);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => n50, 
                           QN => n1964);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => n51, 
                           QN => n1963);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => n52, 
                           QN => n1962);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => n53, 
                           QN => n1961);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => n54, 
                           QN => n1960);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n55, 
                           QN => n1959);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => n56, 
                           QN => n1958);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n57, 
                           QN => n1957);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => n58, 
                           QN => n1956);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n59, 
                           QN => n1955);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => n60, 
                           QN => n1954);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n61, 
                           QN => n1953);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => n62, 
                           QN => n1952);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n63, 
                           QN => n1951);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => n64, 
                           QN => n1950);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n999,
                           QN => n728);
   OUT2_reg_63_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => OUT2(63), QN
                           => n1822);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n1000
                           , QN => n725);
   OUT2_reg_62_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => OUT2(62), QN
                           => n1823);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n1001
                           , QN => n722);
   OUT2_reg_61_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => OUT2(61), QN
                           => n1824);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n1002
                           , QN => n719);
   OUT2_reg_60_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => OUT2(60), QN
                           => n1825);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n1003
                           , QN => n716);
   OUT2_reg_59_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => OUT2(59), QN
                           => n1826);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n1004
                           , QN => n713);
   OUT2_reg_58_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => OUT2(58), QN
                           => n1827);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n1005
                           , QN => n710);
   OUT2_reg_57_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => OUT2(57), QN
                           => n1828);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n1006
                           , QN => n707);
   OUT2_reg_56_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => OUT2(56), QN
                           => n1829);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n1007
                           , QN => n704);
   OUT2_reg_55_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => OUT2(55), QN
                           => n1830);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n1008
                           , QN => n700);
   OUT2_reg_54_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => OUT2(54), QN
                           => n1831);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n1009
                           , QN => n696);
   OUT2_reg_53_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => OUT2(53), QN
                           => n1832);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n1010
                           , QN => n692);
   OUT2_reg_52_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => OUT2(52), QN
                           => n1833);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n1011
                           , QN => n689);
   OUT2_reg_51_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => OUT2(51), QN
                           => n1834);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n1012
                           , QN => n686);
   OUT2_reg_50_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => OUT2(50), QN
                           => n1835);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n1013
                           , QN => n683);
   OUT2_reg_49_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => OUT2(49), QN
                           => n1836);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n1014
                           , QN => n680);
   OUT2_reg_48_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => OUT2(48), QN
                           => n1837);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n1015
                           , QN => n677);
   OUT2_reg_47_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => OUT2(47), QN
                           => n1838);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n1016
                           , QN => n674);
   OUT2_reg_46_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => OUT2(46), QN
                           => n1839);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n1017
                           , QN => n671);
   OUT2_reg_45_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => OUT2(45), QN
                           => n1840);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n1018
                           , QN => n668);
   OUT2_reg_44_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => OUT2(44), QN
                           => n1841);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n1019
                           , QN => n665);
   OUT2_reg_43_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => OUT2(43), QN
                           => n1842);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n1020
                           , QN => n662);
   OUT2_reg_42_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => OUT2(42), QN
                           => n1843);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n1021
                           , QN => n659);
   OUT2_reg_41_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => OUT2(41), QN
                           => n1844);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n1022
                           , QN => n656);
   OUT2_reg_40_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => OUT2(40), QN
                           => n1845);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n1023
                           , QN => n653);
   OUT2_reg_39_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => OUT2(39), QN
                           => n1846);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n1024
                           , QN => n650);
   OUT2_reg_38_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => OUT2(38), QN
                           => n1847);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n1025
                           , QN => n647);
   OUT2_reg_37_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => OUT2(37), QN
                           => n1848);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n1026
                           , QN => n644);
   OUT2_reg_36_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => OUT2(36), QN
                           => n1849);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n1027
                           , QN => n641);
   OUT2_reg_35_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => OUT2(35), QN
                           => n1850);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n1028
                           , QN => n638);
   OUT2_reg_34_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => OUT2(34), QN
                           => n1851);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n1029
                           , QN => n635);
   OUT2_reg_33_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => OUT2(33), QN
                           => n1852);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n1030
                           , QN => n632);
   OUT2_reg_32_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => OUT2(32), QN
                           => n1853);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n1031
                           , QN => n629);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => OUT2(31), QN
                           => n1854);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n1032
                           , QN => n626);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => OUT2(30), QN
                           => n1855);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n1033
                           , QN => n623);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => OUT2(29), QN
                           => n1856);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n1034
                           , QN => n619);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => OUT2(28), QN
                           => n1857);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n1035
                           , QN => n615);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => OUT2(27), QN
                           => n1858);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n1036
                           , QN => n611);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => OUT2(26), QN
                           => n1859);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n1037
                           , QN => n607);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => OUT2(25), QN
                           => n1860);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n1038
                           , QN => n603);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => OUT2(24), QN
                           => n1861);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n1039
                           , QN => n599);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => OUT2(23), QN
                           => n1862);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n1040
                           , QN => n595);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => OUT2(22), QN
                           => n1863);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n1041
                           , QN => n591);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => OUT2(21), QN
                           => n1864);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n1042
                           , QN => n587);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => OUT2(20), QN
                           => n1865);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n1043
                           , QN => n583);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => OUT2(19), QN
                           => n1866);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n1044
                           , QN => n580);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => OUT2(18), QN
                           => n1867);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n1045
                           , QN => n577);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => OUT2(17), QN
                           => n1868);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n1046
                           , QN => n574);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => OUT2(16), QN
                           => n1869);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n1047
                           , QN => n571);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => OUT2(15), QN
                           => n1870);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n1048
                           , QN => n568);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => OUT2(14), QN
                           => n1871);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n1049
                           , QN => n565);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => OUT2(13), QN
                           => n1872);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n1050
                           , QN => n562);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => OUT2(12), QN
                           => n1873);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n1051
                           , QN => n559);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => OUT2(11), QN
                           => n1874);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n1052
                           , QN => n556);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => OUT2(10), QN
                           => n1875);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n1053,
                           QN => n553);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => OUT2(9), QN 
                           => n1876);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => n1054,
                           QN => n550);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => OUT2(8), QN 
                           => n1877);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => n1055,
                           QN => n547);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => OUT2(7), QN 
                           => n1878);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => n1056,
                           QN => n544);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => OUT2(6), QN 
                           => n1879);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => n1057,
                           QN => n541);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => OUT2(5), QN 
                           => n1880);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => n1058,
                           QN => n538);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => OUT2(4), QN 
                           => n1881);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => n1059,
                           QN => n535);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => OUT2(3), QN 
                           => n1882);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n1060,
                           QN => n532);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => OUT2(2), QN 
                           => n1883);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n1061,
                           QN => n529);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => OUT2(1), QN 
                           => n1884);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n1062,
                           QN => n522);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => OUT2(0), QN 
                           => n1885);
   OUT1_reg_63_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => OUT1(63), QN
                           => n1886);
   OUT1_reg_62_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => OUT1(62), QN
                           => n1887);
   OUT1_reg_61_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => OUT1(61), QN
                           => n1888);
   OUT1_reg_60_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => OUT1(60), QN
                           => n1889);
   OUT1_reg_59_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => OUT1(59), QN
                           => n1890);
   OUT1_reg_58_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => OUT1(58), QN
                           => n1891);
   OUT1_reg_57_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => OUT1(57), QN
                           => n1892);
   OUT1_reg_56_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => OUT1(56), QN
                           => n1893);
   OUT1_reg_55_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => OUT1(55), QN
                           => n1894);
   OUT1_reg_54_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => OUT1(54), QN
                           => n1895);
   OUT1_reg_53_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => OUT1(53), QN
                           => n1896);
   OUT1_reg_52_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => OUT1(52), QN
                           => n1897);
   OUT1_reg_51_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => OUT1(51), QN
                           => n1898);
   OUT1_reg_50_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => OUT1(50), QN
                           => n1899);
   OUT1_reg_49_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => OUT1(49), QN
                           => n1900);
   OUT1_reg_48_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => OUT1(48), QN
                           => n1901);
   OUT1_reg_47_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => OUT1(47), QN
                           => n1902);
   OUT1_reg_46_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => OUT1(46), QN
                           => n1903);
   OUT1_reg_45_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => OUT1(45), QN
                           => n1904);
   OUT1_reg_44_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => OUT1(44), QN
                           => n1905);
   OUT1_reg_43_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => OUT1(43), QN
                           => n1906);
   OUT1_reg_42_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => OUT1(42), QN
                           => n1907);
   OUT1_reg_41_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => OUT1(41), QN
                           => n1908);
   OUT1_reg_40_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => OUT1(40), QN
                           => n1909);
   OUT1_reg_39_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => OUT1(39), QN
                           => n1910);
   OUT1_reg_38_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => OUT1(38), QN
                           => n1911);
   OUT1_reg_37_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => OUT1(37), QN
                           => n1912);
   OUT1_reg_36_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => OUT1(36), QN
                           => n1913);
   OUT1_reg_35_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => OUT1(35), QN
                           => n1914);
   OUT1_reg_34_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => OUT1(34), QN
                           => n1915);
   OUT1_reg_33_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => OUT1(33), QN
                           => n1916);
   OUT1_reg_32_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => OUT1(32), QN
                           => n1917);
   OUT1_reg_31_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => OUT1(31), QN
                           => n1918);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => OUT1(30), QN
                           => n1919);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => OUT1(29), QN
                           => n1920);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => OUT1(28), QN
                           => n1921);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => OUT1(27), QN
                           => n1922);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => OUT1(26), QN
                           => n1923);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => OUT1(25), QN
                           => n1924);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => OUT1(24), QN
                           => n1925);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => OUT1(23), QN
                           => n1926);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => OUT1(22), QN
                           => n1927);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => OUT1(21), QN
                           => n1928);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => OUT1(20), QN
                           => n1929);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => OUT1(19), QN
                           => n1930);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => OUT1(18), QN
                           => n1931);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => OUT1(17), QN
                           => n1932);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => OUT1(16), QN
                           => n1933);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => OUT1(15), QN
                           => n1934);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => OUT1(14), QN
                           => n1935);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => OUT1(13), QN
                           => n1936);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => OUT1(12), QN
                           => n1937);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => OUT1(11), QN
                           => n1938);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => OUT1(10), QN
                           => n1939);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => OUT1(9), QN 
                           => n1940);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => OUT1(8), QN 
                           => n1941);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => OUT1(7), QN 
                           => n1942);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => OUT1(6), QN 
                           => n1943);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => OUT1(5), QN 
                           => n1944);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => OUT1(4), QN 
                           => n1945);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => OUT1(3), QN 
                           => n1946);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => OUT1(2), QN 
                           => n1947);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => OUT1(1), QN 
                           => n1948);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => OUT1(0), QN 
                           => n1949);
   U859 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n2164, A3 => ADD_RD1(1), 
                           ZN => n521);
   U860 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n2135, A3 => ADD_RD2(1), 
                           ZN => n735);
   U861 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n873, A3 => ADD_WR(1), ZN 
                           => n872);
   U862 : NAND3_X1 port map( A1 => n873, A2 => n2175, A3 => ADD_WR(1), ZN => 
                           n936);
   U863 : NAND3_X1 port map( A1 => n873, A2 => n2176, A3 => ADD_WR(0), ZN => 
                           n975);
   U864 : NAND3_X1 port map( A1 => n2175, A2 => n2176, A3 => n873, ZN => n998);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => n537, 
                           QN => n1818);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => n534, 
                           QN => n1819);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => n531, 
                           QN => n1820);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => n528, 
                           QN => n1821);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => n730,
                           QN => n415);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => n702,
                           QN => n1200);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => n698,
                           QN => n1202);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => n694,
                           QN => n1204);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => n622,
                           QN => n1793);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => n618,
                           QN => n1794);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => n614,
                           QN => n1795);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => n610,
                           QN => n1796);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => n606,
                           QN => n1797);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => n602,
                           QN => n1798);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => n598,
                           QN => n1799);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => n594,
                           QN => n1800);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => n590,
                           QN => n1801);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => n586,
                           QN => n1802);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => n582,
                           QN => n1803);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => n579,
                           QN => n1804);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => n576,
                           QN => n1805);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => n573,
                           QN => n1806);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => n570,
                           QN => n1807);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => n567,
                           QN => n1808);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => n564,
                           QN => n1809);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => n561,
                           QN => n1810);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => n558,
                           QN => n1811);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => n555, 
                           QN => n1812);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => n552, 
                           QN => n1813);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => n549, 
                           QN => n1814);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => n546, 
                           QN => n1815);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => n543, 
                           QN => n1816);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => n540, 
                           QN => n1817);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => n731,
                           QN => n1694);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => n727,
                           QN => n1695);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => n724,
                           QN => n1696);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => n721,
                           QN => n1697);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => n718,
                           QN => n1698);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => n715,
                           QN => n1699);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => n712,
                           QN => n1700);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => n709,
                           QN => n1701);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => n706,
                           QN => n1702);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => n703,
                           QN => n1703);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => n699,
                           QN => n1704);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => n695,
                           QN => n1705);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => n691,
                           QN => n1706);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => n688,
                           QN => n1707);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => n685,
                           QN => n1708);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => n682,
                           QN => n1709);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => n679,
                           QN => n1710);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => n676,
                           QN => n1711);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => n673,
                           QN => n1712);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => n670,
                           QN => n1713);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => n667,
                           QN => n1714);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => n664,
                           QN => n1715);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => n661,
                           QN => n1716);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => n658,
                           QN => n1717);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => n655,
                           QN => n1718);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => n652,
                           QN => n1719);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => n649,
                           QN => n1720);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => n646,
                           QN => n1721);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => n643,
                           QN => n1722);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => n640,
                           QN => n1723);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => n637,
                           QN => n1724);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => n634,
                           QN => n1725);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => n631,
                           QN => n1726);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => n628,
                           QN => n1727);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n625,
                           QN => n1728);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => n621,
                           QN => n1729);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => n617,
                           QN => n1730);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => n613,
                           QN => n1731);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => n609,
                           QN => n1732);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => n605,
                           QN => n1733);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => n601,
                           QN => n1734);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => n597,
                           QN => n1735);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => n593,
                           QN => n1736);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => n589,
                           QN => n1737);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => n585,
                           QN => n1738);
   U3 : BUF_X1 port map( A => n521, Z => n2167);
   U4 : BUF_X1 port map( A => n521, Z => n2166);
   U5 : BUF_X1 port map( A => n521, Z => n2165);
   U6 : BUF_X1 port map( A => n735, Z => n2139);
   U7 : BUF_X1 port map( A => n735, Z => n2138);
   U8 : BUF_X1 port map( A => n735, Z => n2137);
   U9 : BUF_X1 port map( A => n735, Z => n2136);
   U10 : BUF_X1 port map( A => n521, Z => n2169);
   U11 : BUF_X1 port map( A => n521, Z => n2168);
   U12 : BUF_X1 port map( A => n735, Z => n2140);
   U13 : BUF_X1 port map( A => n526, Z => n2151);
   U14 : BUF_X1 port map( A => n526, Z => n2152);
   U15 : BUF_X1 port map( A => n527, Z => n2144);
   U16 : BUF_X1 port map( A => n527, Z => n2146);
   U17 : BUF_X1 port map( A => n527, Z => n2145);
   U18 : BUF_X1 port map( A => n523, Z => n2159);
   U19 : BUF_X1 port map( A => n523, Z => n2160);
   U20 : BUF_X1 port map( A => n523, Z => n2161);
   U21 : BUF_X1 port map( A => n523, Z => n2162);
   U22 : BUF_X1 port map( A => n523, Z => n2163);
   U23 : BUF_X1 port map( A => n736, Z => n2130);
   U24 : BUF_X1 port map( A => n736, Z => n2131);
   U25 : BUF_X1 port map( A => n736, Z => n2132);
   U26 : BUF_X1 port map( A => n736, Z => n2133);
   U27 : BUF_X1 port map( A => n736, Z => n2134);
   U28 : BUF_X1 port map( A => n525, Z => n2154);
   U29 : BUF_X1 port map( A => n525, Z => n2155);
   U30 : BUF_X1 port map( A => n525, Z => n2156);
   U31 : BUF_X1 port map( A => n525, Z => n2157);
   U32 : BUF_X1 port map( A => n738, Z => n2128);
   U33 : BUF_X1 port map( A => n738, Z => n2127);
   U34 : BUF_X1 port map( A => n738, Z => n2126);
   U35 : BUF_X1 port map( A => n738, Z => n2125);
   U36 : BUF_X1 port map( A => n738, Z => n2124);
   U37 : BUF_X1 port map( A => n742, Z => n2104);
   U38 : BUF_X1 port map( A => n742, Z => n2103);
   U39 : BUF_X1 port map( A => n742, Z => n2102);
   U40 : BUF_X1 port map( A => n742, Z => n2101);
   U41 : BUF_X1 port map( A => n739, Z => n2122);
   U42 : BUF_X1 port map( A => n739, Z => n2121);
   U43 : BUF_X1 port map( A => n739, Z => n2120);
   U44 : BUF_X1 port map( A => n739, Z => n2119);
   U45 : BUF_X1 port map( A => n739, Z => n2118);
   U46 : BUF_X1 port map( A => n740, Z => n2116);
   U47 : BUF_X1 port map( A => n740, Z => n2115);
   U48 : BUF_X1 port map( A => n740, Z => n2114);
   U49 : BUF_X1 port map( A => n740, Z => n2113);
   U50 : BUF_X1 port map( A => n740, Z => n2112);
   U51 : BUF_X1 port map( A => n741, Z => n2106);
   U52 : BUF_X1 port map( A => n875, Z => n2094);
   U53 : BUF_X1 port map( A => n938, Z => n2082);
   U54 : BUF_X1 port map( A => n978, Z => n2070);
   U55 : BUF_X1 port map( A => n741, Z => n2110);
   U56 : BUF_X1 port map( A => n741, Z => n2109);
   U57 : BUF_X1 port map( A => n741, Z => n2108);
   U58 : BUF_X1 port map( A => n741, Z => n2107);
   U59 : BUF_X1 port map( A => n875, Z => n2098);
   U60 : BUF_X1 port map( A => n875, Z => n2097);
   U61 : BUF_X1 port map( A => n875, Z => n2096);
   U62 : BUF_X1 port map( A => n875, Z => n2095);
   U63 : BUF_X1 port map( A => n938, Z => n2086);
   U64 : BUF_X1 port map( A => n938, Z => n2085);
   U65 : BUF_X1 port map( A => n938, Z => n2084);
   U66 : BUF_X1 port map( A => n938, Z => n2083);
   U67 : BUF_X1 port map( A => n978, Z => n2074);
   U68 : BUF_X1 port map( A => n978, Z => n2073);
   U69 : BUF_X1 port map( A => n978, Z => n2072);
   U70 : BUF_X1 port map( A => n978, Z => n2071);
   U71 : BUF_X1 port map( A => n526, Z => n2148);
   U72 : BUF_X1 port map( A => n526, Z => n2150);
   U73 : BUF_X1 port map( A => n876, Z => n2092);
   U74 : BUF_X1 port map( A => n876, Z => n2091);
   U75 : BUF_X1 port map( A => n876, Z => n2090);
   U76 : BUF_X1 port map( A => n876, Z => n2089);
   U77 : BUF_X1 port map( A => n876, Z => n2088);
   U78 : BUF_X1 port map( A => n939, Z => n2080);
   U79 : BUF_X1 port map( A => n939, Z => n2079);
   U80 : BUF_X1 port map( A => n939, Z => n2078);
   U81 : BUF_X1 port map( A => n939, Z => n2077);
   U82 : BUF_X1 port map( A => n939, Z => n2076);
   U83 : BUF_X1 port map( A => n979, Z => n2068);
   U84 : BUF_X1 port map( A => n979, Z => n2067);
   U85 : BUF_X1 port map( A => n979, Z => n2066);
   U86 : BUF_X1 port map( A => n979, Z => n2065);
   U87 : BUF_X1 port map( A => n979, Z => n2064);
   U88 : BUF_X1 port map( A => n527, Z => n2143);
   U89 : BUF_X1 port map( A => n527, Z => n2142);
   U90 : BUF_X1 port map( A => n526, Z => n2149);
   U91 : BUF_X1 port map( A => n525, Z => n2153);
   U92 : BUF_X1 port map( A => n742, Z => n2100);
   U93 : NAND2_X1 port map( A1 => n734, A2 => n872, ZN => n741);
   U94 : NAND2_X1 port map( A1 => n734, A2 => n936, ZN => n875);
   U95 : NAND2_X1 port map( A1 => n734, A2 => n2094, ZN => n876);
   U96 : NAND2_X1 port map( A1 => n734, A2 => n975, ZN => n938);
   U97 : NAND2_X1 port map( A1 => n734, A2 => n2082, ZN => n939);
   U98 : NAND2_X1 port map( A1 => n734, A2 => n998, ZN => n978);
   U99 : NAND2_X1 port map( A1 => n734, A2 => n2070, ZN => n979);
   U100 : OAI22_X1 port map( A1 => n538, A2 => n2111, B1 => n2104, B2 => n751, 
                           ZN => n1620);
   U101 : OAI22_X1 port map( A1 => n541, A2 => n2110, B1 => n2104, B2 => n753, 
                           ZN => n1618);
   U102 : OAI22_X1 port map( A1 => n544, A2 => n2110, B1 => n2104, B2 => n755, 
                           ZN => n1616);
   U103 : OAI22_X1 port map( A1 => n547, A2 => n2110, B1 => n2104, B2 => n757, 
                           ZN => n1614);
   U104 : OAI22_X1 port map( A1 => n550, A2 => n2110, B1 => n2104, B2 => n759, 
                           ZN => n1612);
   U105 : OAI22_X1 port map( A1 => n553, A2 => n2110, B1 => n2104, B2 => n761, 
                           ZN => n1610);
   U106 : OAI22_X1 port map( A1 => n556, A2 => n2110, B1 => n2104, B2 => n763, 
                           ZN => n1608);
   U107 : OAI22_X1 port map( A1 => n559, A2 => n2110, B1 => n2104, B2 => n765, 
                           ZN => n1606);
   U108 : OAI22_X1 port map( A1 => n562, A2 => n2110, B1 => n2104, B2 => n767, 
                           ZN => n1604);
   U109 : OAI22_X1 port map( A1 => n565, A2 => n2110, B1 => n2104, B2 => n769, 
                           ZN => n1602);
   U110 : OAI22_X1 port map( A1 => n568, A2 => n2110, B1 => n2104, B2 => n771, 
                           ZN => n1600);
   U111 : OAI22_X1 port map( A1 => n571, A2 => n2110, B1 => n2104, B2 => n773, 
                           ZN => n1598);
   U112 : OAI22_X1 port map( A1 => n574, A2 => n2110, B1 => n2103, B2 => n775, 
                           ZN => n1596);
   U113 : OAI22_X1 port map( A1 => n577, A2 => n2109, B1 => n2103, B2 => n777, 
                           ZN => n1594);
   U114 : OAI22_X1 port map( A1 => n580, A2 => n2109, B1 => n2103, B2 => n779, 
                           ZN => n1592);
   U115 : OAI22_X1 port map( A1 => n583, A2 => n2109, B1 => n2103, B2 => n781, 
                           ZN => n1590);
   U116 : OAI22_X1 port map( A1 => n587, A2 => n2109, B1 => n2103, B2 => n783, 
                           ZN => n1588);
   U117 : OAI22_X1 port map( A1 => n591, A2 => n2109, B1 => n2103, B2 => n785, 
                           ZN => n1586);
   U118 : OAI22_X1 port map( A1 => n595, A2 => n2109, B1 => n2103, B2 => n787, 
                           ZN => n1584);
   U119 : OAI22_X1 port map( A1 => n599, A2 => n2109, B1 => n2103, B2 => n789, 
                           ZN => n1582);
   U120 : OAI22_X1 port map( A1 => n603, A2 => n2109, B1 => n2103, B2 => n791, 
                           ZN => n1580);
   U121 : OAI22_X1 port map( A1 => n607, A2 => n2109, B1 => n2103, B2 => n793, 
                           ZN => n1578);
   U122 : OAI22_X1 port map( A1 => n611, A2 => n2109, B1 => n2103, B2 => n795, 
                           ZN => n1576);
   U123 : OAI22_X1 port map( A1 => n615, A2 => n2109, B1 => n2103, B2 => n797, 
                           ZN => n1574);
   U124 : OAI22_X1 port map( A1 => n619, A2 => n2109, B1 => n2102, B2 => n799, 
                           ZN => n1572);
   U125 : OAI22_X1 port map( A1 => n623, A2 => n2108, B1 => n2102, B2 => n801, 
                           ZN => n1570);
   U126 : OAI22_X1 port map( A1 => n626, A2 => n2108, B1 => n2102, B2 => n803, 
                           ZN => n1568);
   U127 : OAI22_X1 port map( A1 => n629, A2 => n2108, B1 => n2102, B2 => n805, 
                           ZN => n1566);
   U128 : OAI22_X1 port map( A1 => n632, A2 => n2108, B1 => n2102, B2 => n807, 
                           ZN => n1564);
   U129 : OAI22_X1 port map( A1 => n635, A2 => n2108, B1 => n2102, B2 => n809, 
                           ZN => n1562);
   U130 : OAI22_X1 port map( A1 => n638, A2 => n2108, B1 => n2102, B2 => n811, 
                           ZN => n1560);
   U131 : OAI22_X1 port map( A1 => n641, A2 => n2108, B1 => n2102, B2 => n813, 
                           ZN => n1558);
   U132 : OAI22_X1 port map( A1 => n644, A2 => n2108, B1 => n2102, B2 => n815, 
                           ZN => n1556);
   U133 : OAI22_X1 port map( A1 => n647, A2 => n2108, B1 => n2102, B2 => n817, 
                           ZN => n1554);
   U134 : OAI22_X1 port map( A1 => n650, A2 => n2108, B1 => n2102, B2 => n819, 
                           ZN => n1552);
   U135 : OAI22_X1 port map( A1 => n653, A2 => n2108, B1 => n2102, B2 => n821, 
                           ZN => n1550);
   U136 : OAI22_X1 port map( A1 => n656, A2 => n2108, B1 => n2101, B2 => n823, 
                           ZN => n1548);
   U137 : OAI22_X1 port map( A1 => n659, A2 => n2107, B1 => n2101, B2 => n825, 
                           ZN => n1546);
   U138 : OAI22_X1 port map( A1 => n662, A2 => n2107, B1 => n2101, B2 => n827, 
                           ZN => n1544);
   U139 : OAI22_X1 port map( A1 => n665, A2 => n2107, B1 => n2101, B2 => n829, 
                           ZN => n1542);
   U140 : OAI22_X1 port map( A1 => n668, A2 => n2107, B1 => n2101, B2 => n831, 
                           ZN => n1540);
   U141 : OAI22_X1 port map( A1 => n671, A2 => n2107, B1 => n2101, B2 => n833, 
                           ZN => n1538);
   U142 : OAI22_X1 port map( A1 => n674, A2 => n2107, B1 => n2101, B2 => n835, 
                           ZN => n1536);
   U143 : OAI22_X1 port map( A1 => n677, A2 => n2107, B1 => n2101, B2 => n837, 
                           ZN => n1534);
   U144 : OAI22_X1 port map( A1 => n680, A2 => n2107, B1 => n2101, B2 => n839, 
                           ZN => n1532);
   U145 : OAI22_X1 port map( A1 => n683, A2 => n2107, B1 => n2101, B2 => n841, 
                           ZN => n1530);
   U146 : OAI22_X1 port map( A1 => n686, A2 => n2107, B1 => n2101, B2 => n843, 
                           ZN => n1528);
   U147 : OAI22_X1 port map( A1 => n689, A2 => n2107, B1 => n2101, B2 => n845, 
                           ZN => n1526);
   U148 : OAI22_X1 port map( A1 => n522, A2 => n2111, B1 => n2105, B2 => n743, 
                           ZN => n1628);
   U149 : OAI22_X1 port map( A1 => n529, A2 => n2111, B1 => n2105, B2 => n745, 
                           ZN => n1626);
   U150 : OAI22_X1 port map( A1 => n532, A2 => n2111, B1 => n2105, B2 => n747, 
                           ZN => n1624);
   U151 : OAI22_X1 port map( A1 => n535, A2 => n2111, B1 => n2105, B2 => n749, 
                           ZN => n1622);
   U152 : OAI22_X1 port map( A1 => n692, A2 => n2107, B1 => n2100, B2 => n847, 
                           ZN => n1524);
   U153 : OAI22_X1 port map( A1 => n696, A2 => n2106, B1 => n2100, B2 => n849, 
                           ZN => n1522);
   U154 : OAI22_X1 port map( A1 => n700, A2 => n2106, B1 => n2100, B2 => n851, 
                           ZN => n1520);
   U155 : OAI22_X1 port map( A1 => n704, A2 => n2106, B1 => n2100, B2 => n853, 
                           ZN => n1518);
   U156 : OAI22_X1 port map( A1 => n707, A2 => n2106, B1 => n2100, B2 => n855, 
                           ZN => n1516);
   U157 : OAI22_X1 port map( A1 => n710, A2 => n2106, B1 => n2100, B2 => n857, 
                           ZN => n1514);
   U158 : OAI22_X1 port map( A1 => n713, A2 => n2106, B1 => n2100, B2 => n859, 
                           ZN => n1512);
   U159 : OAI22_X1 port map( A1 => n716, A2 => n2106, B1 => n2100, B2 => n861, 
                           ZN => n1510);
   U160 : OAI22_X1 port map( A1 => n719, A2 => n2106, B1 => n2100, B2 => n863, 
                           ZN => n1508);
   U161 : OAI22_X1 port map( A1 => n722, A2 => n2106, B1 => n2100, B2 => n865, 
                           ZN => n1506);
   U162 : OAI22_X1 port map( A1 => n725, A2 => n2106, B1 => n2100, B2 => n867, 
                           ZN => n1504);
   U163 : OAI22_X1 port map( A1 => n728, A2 => n2106, B1 => n2100, B2 => n871, 
                           ZN => n1502);
   U164 : AND3_X1 port map( A1 => n2173, A2 => n2174, A3 => n2164, ZN => n526);
   U165 : AND3_X1 port map( A1 => n2164, A2 => n2174, A3 => ADD_RD1(0), ZN => 
                           n527);
   U166 : AND3_X1 port map( A1 => n2164, A2 => n2173, A3 => ADD_RD1(1), ZN => 
                           n525);
   U167 : NAND2_X1 port map( A1 => n734, A2 => n2106, ZN => n742);
   U168 : AND3_X1 port map( A1 => n2135, A2 => n2172, A3 => ADD_RD2(0), ZN => 
                           n740);
   U169 : AND3_X1 port map( A1 => n2135, A2 => n2171, A3 => ADD_RD2(1), ZN => 
                           n738);
   U170 : AND3_X1 port map( A1 => n2171, A2 => n2172, A3 => n2135, ZN => n739);
   U171 : AND2_X1 port map( A1 => RD1, A2 => n734, ZN => n523);
   U172 : AND2_X1 port map( A1 => RD2, A2 => n734, ZN => n736);
   U173 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n873);
   U174 : OAI221_X1 port map( B1 => n2169, B2 => n562, C1 => n1937, C2 => n2160
                           , A => n563, ZN => n1681);
   U175 : AOI222_X1 port map( A1 => n52, A2 => n2153, B1 => n180, B2 => n2149, 
                           C1 => n2146, C2 => n564, ZN => n563);
   U176 : OAI221_X1 port map( B1 => n2169, B2 => n565, C1 => n1936, C2 => n2160
                           , A => n566, ZN => n1680);
   U177 : AOI222_X1 port map( A1 => n51, A2 => n2154, B1 => n179, B2 => n2149, 
                           C1 => n2146, C2 => n567, ZN => n566);
   U178 : OAI221_X1 port map( B1 => n2169, B2 => n568, C1 => n1935, C2 => n2160
                           , A => n569, ZN => n1679);
   U179 : AOI222_X1 port map( A1 => n50, A2 => n2154, B1 => n178, B2 => n2149, 
                           C1 => n2146, C2 => n570, ZN => n569);
   U180 : OAI221_X1 port map( B1 => n2169, B2 => n571, C1 => n1934, C2 => n2161
                           , A => n572, ZN => n1678);
   U181 : AOI222_X1 port map( A1 => n49, A2 => n2154, B1 => n177, B2 => n2149, 
                           C1 => n2145, C2 => n573, ZN => n572);
   U182 : OAI221_X1 port map( B1 => n2168, B2 => n574, C1 => n1933, C2 => n2160
                           , A => n575, ZN => n1677);
   U183 : AOI222_X1 port map( A1 => n48, A2 => n2154, B1 => n176, B2 => n2149, 
                           C1 => n2145, C2 => n576, ZN => n575);
   U184 : OAI221_X1 port map( B1 => n2168, B2 => n577, C1 => n1932, C2 => n2160
                           , A => n578, ZN => n1676);
   U185 : AOI222_X1 port map( A1 => n47, A2 => n2154, B1 => n175, B2 => n2149, 
                           C1 => n2145, C2 => n579, ZN => n578);
   U186 : OAI221_X1 port map( B1 => n2168, B2 => n580, C1 => n1931, C2 => n2160
                           , A => n581, ZN => n1675);
   U187 : AOI222_X1 port map( A1 => n46, A2 => n2154, B1 => n174, B2 => n2149, 
                           C1 => n2145, C2 => n582, ZN => n581);
   U188 : OAI221_X1 port map( B1 => n538, B2 => n2140, C1 => n1881, C2 => n2130
                           , A => n750, ZN => n1621);
   U189 : AOI222_X1 port map( A1 => n2128, A2 => n60, B1 => n2122, B2 => n188, 
                           C1 => n2116, C2 => n540, ZN => n750);
   U190 : OAI221_X1 port map( B1 => n541, B2 => n2140, C1 => n1880, C2 => n2130
                           , A => n752, ZN => n1619);
   U191 : AOI222_X1 port map( A1 => n2128, A2 => n59, B1 => n2122, B2 => n187, 
                           C1 => n2116, C2 => n543, ZN => n752);
   U192 : OAI221_X1 port map( B1 => n544, B2 => n2140, C1 => n1879, C2 => n2130
                           , A => n754, ZN => n1617);
   U193 : AOI222_X1 port map( A1 => n2128, A2 => n58, B1 => n2122, B2 => n186, 
                           C1 => n2116, C2 => n546, ZN => n754);
   U194 : OAI221_X1 port map( B1 => n547, B2 => n2140, C1 => n1878, C2 => n2130
                           , A => n756, ZN => n1615);
   U195 : AOI222_X1 port map( A1 => n2128, A2 => n57, B1 => n2122, B2 => n185, 
                           C1 => n2116, C2 => n549, ZN => n756);
   U196 : OAI221_X1 port map( B1 => n550, B2 => n2140, C1 => n1877, C2 => n2130
                           , A => n758, ZN => n1613);
   U197 : AOI222_X1 port map( A1 => n2128, A2 => n56, B1 => n2122, B2 => n184, 
                           C1 => n2116, C2 => n552, ZN => n758);
   U198 : OAI221_X1 port map( B1 => n553, B2 => n2140, C1 => n1876, C2 => n2130
                           , A => n760, ZN => n1611);
   U199 : AOI222_X1 port map( A1 => n2128, A2 => n55, B1 => n2122, B2 => n183, 
                           C1 => n2116, C2 => n555, ZN => n760);
   U200 : OAI221_X1 port map( B1 => n556, B2 => n2140, C1 => n1875, C2 => n2130
                           , A => n762, ZN => n1609);
   U201 : AOI222_X1 port map( A1 => n2128, A2 => n54, B1 => n2122, B2 => n182, 
                           C1 => n2116, C2 => n558, ZN => n762);
   U202 : OAI221_X1 port map( B1 => n559, B2 => n2140, C1 => n1874, C2 => n2130
                           , A => n764, ZN => n1607);
   U203 : AOI222_X1 port map( A1 => n2128, A2 => n53, B1 => n2122, B2 => n181, 
                           C1 => n2116, C2 => n561, ZN => n764);
   U204 : OAI221_X1 port map( B1 => n562, B2 => n2140, C1 => n1873, C2 => n2131
                           , A => n766, ZN => n1605);
   U205 : AOI222_X1 port map( A1 => n2128, A2 => n52, B1 => n2122, B2 => n180, 
                           C1 => n2116, C2 => n564, ZN => n766);
   U206 : OAI221_X1 port map( B1 => n565, B2 => n2140, C1 => n1872, C2 => n2131
                           , A => n768, ZN => n1603);
   U207 : AOI222_X1 port map( A1 => n2128, A2 => n51, B1 => n2122, B2 => n179, 
                           C1 => n2116, C2 => n567, ZN => n768);
   U208 : OAI221_X1 port map( B1 => n568, B2 => n2140, C1 => n1871, C2 => n2131
                           , A => n770, ZN => n1601);
   U209 : AOI222_X1 port map( A1 => n2128, A2 => n50, B1 => n2122, B2 => n178, 
                           C1 => n2116, C2 => n570, ZN => n770);
   U210 : OAI221_X1 port map( B1 => n571, B2 => n2140, C1 => n1870, C2 => n2132
                           , A => n772, ZN => n1599);
   U211 : AOI222_X1 port map( A1 => n2128, A2 => n49, B1 => n2122, B2 => n177, 
                           C1 => n2116, C2 => n573, ZN => n772);
   U212 : OAI221_X1 port map( B1 => n574, B2 => n2139, C1 => n1869, C2 => n2131
                           , A => n774, ZN => n1597);
   U213 : AOI222_X1 port map( A1 => n2127, A2 => n48, B1 => n2121, B2 => n176, 
                           C1 => n2115, C2 => n576, ZN => n774);
   U214 : OAI221_X1 port map( B1 => n577, B2 => n2139, C1 => n1868, C2 => n2131
                           , A => n776, ZN => n1595);
   U215 : AOI222_X1 port map( A1 => n2127, A2 => n47, B1 => n2121, B2 => n175, 
                           C1 => n2115, C2 => n579, ZN => n776);
   U216 : OAI221_X1 port map( B1 => n580, B2 => n2139, C1 => n1867, C2 => n2131
                           , A => n778, ZN => n1593);
   U217 : AOI222_X1 port map( A1 => n2127, A2 => n46, B1 => n2121, B2 => n174, 
                           C1 => n2115, C2 => n582, ZN => n778);
   U218 : OAI221_X1 port map( B1 => n2166, B2 => n656, C1 => n1909, C2 => n2162
                           , A => n657, ZN => n1653);
   U219 : AOI222_X1 port map( A1 => n24, A2 => n2156, B1 => n2151, B2 => n658, 
                           C1 => n88, C2 => n2143, ZN => n657);
   U220 : OAI221_X1 port map( B1 => n2166, B2 => n659, C1 => n1908, C2 => n2162
                           , A => n660, ZN => n1652);
   U221 : AOI222_X1 port map( A1 => n23, A2 => n2156, B1 => n2151, B2 => n661, 
                           C1 => n87, C2 => n2143, ZN => n660);
   U222 : OAI221_X1 port map( B1 => n2166, B2 => n662, C1 => n1907, C2 => n2162
                           , A => n663, ZN => n1651);
   U223 : AOI222_X1 port map( A1 => n22, A2 => n2156, B1 => n2151, B2 => n664, 
                           C1 => n86, C2 => n2143, ZN => n663);
   U224 : OAI221_X1 port map( B1 => n2166, B2 => n665, C1 => n1906, C2 => n2162
                           , A => n666, ZN => n1650);
   U225 : AOI222_X1 port map( A1 => n21, A2 => n2156, B1 => n2151, B2 => n667, 
                           C1 => n85, C2 => n2143, ZN => n666);
   U226 : OAI221_X1 port map( B1 => n2166, B2 => n668, C1 => n1905, C2 => n2162
                           , A => n669, ZN => n1649);
   U227 : AOI222_X1 port map( A1 => n20, A2 => n2156, B1 => n2151, B2 => n670, 
                           C1 => n84, C2 => n2143, ZN => n669);
   U228 : OAI221_X1 port map( B1 => n2166, B2 => n671, C1 => n1904, C2 => n2162
                           , A => n672, ZN => n1648);
   U229 : AOI222_X1 port map( A1 => n19, A2 => n2156, B1 => n2151, B2 => n673, 
                           C1 => n83, C2 => n2143, ZN => n672);
   U230 : OAI221_X1 port map( B1 => n2166, B2 => n674, C1 => n1903, C2 => n2162
                           , A => n675, ZN => n1647);
   U231 : AOI222_X1 port map( A1 => n18, A2 => n2156, B1 => n2151, B2 => n676, 
                           C1 => n82, C2 => n2143, ZN => n675);
   U232 : OAI221_X1 port map( B1 => n2166, B2 => n677, C1 => n1902, C2 => n2162
                           , A => n678, ZN => n1646);
   U233 : AOI222_X1 port map( A1 => n17, A2 => n2156, B1 => n2151, B2 => n679, 
                           C1 => n81, C2 => n2143, ZN => n678);
   U234 : OAI221_X1 port map( B1 => n2166, B2 => n680, C1 => n1901, C2 => n2163
                           , A => n681, ZN => n1645);
   U235 : AOI222_X1 port map( A1 => n16, A2 => n2157, B1 => n2151, B2 => n682, 
                           C1 => n80, C2 => n2143, ZN => n681);
   U236 : OAI221_X1 port map( B1 => n2166, B2 => n683, C1 => n1900, C2 => n2163
                           , A => n684, ZN => n1644);
   U237 : AOI222_X1 port map( A1 => n15, A2 => n2157, B1 => n2151, B2 => n685, 
                           C1 => n79, C2 => n2143, ZN => n684);
   U238 : OAI221_X1 port map( B1 => n2166, B2 => n686, C1 => n1899, C2 => n2163
                           , A => n687, ZN => n1643);
   U239 : AOI222_X1 port map( A1 => n14, A2 => n2157, B1 => n2152, B2 => n688, 
                           C1 => n78, C2 => n2143, ZN => n687);
   U240 : OAI221_X1 port map( B1 => n2166, B2 => n689, C1 => n1898, C2 => n2163
                           , A => n690, ZN => n1642);
   U241 : AOI222_X1 port map( A1 => n13, A2 => n2157, B1 => n2152, B2 => n691, 
                           C1 => n77, C2 => n2143, ZN => n690);
   U242 : OAI221_X1 port map( B1 => n2165, B2 => n692, C1 => n1897, C2 => n2163
                           , A => n693, ZN => n1641);
   U243 : AOI222_X1 port map( A1 => n2158, A2 => n694, B1 => n2152, B2 => n695,
                           C1 => n76, C2 => n2142, ZN => n693);
   U244 : OAI221_X1 port map( B1 => n2165, B2 => n696, C1 => n1896, C2 => n2163
                           , A => n697, ZN => n1640);
   U245 : AOI222_X1 port map( A1 => n2158, A2 => n698, B1 => n2152, B2 => n699,
                           C1 => n75, C2 => n2142, ZN => n697);
   U246 : OAI221_X1 port map( B1 => n2165, B2 => n700, C1 => n1895, C2 => n2163
                           , A => n701, ZN => n1639);
   U247 : AOI222_X1 port map( A1 => n2158, A2 => n702, B1 => n2152, B2 => n703,
                           C1 => n74, C2 => n2142, ZN => n701);
   U248 : OAI221_X1 port map( B1 => n2165, B2 => n704, C1 => n1894, C2 => n2163
                           , A => n705, ZN => n1638);
   U249 : AOI222_X1 port map( A1 => n9, A2 => n2157, B1 => n2152, B2 => n706, 
                           C1 => n73, C2 => n2142, ZN => n705);
   U250 : OAI221_X1 port map( B1 => n2165, B2 => n707, C1 => n1893, C2 => n2163
                           , A => n708, ZN => n1637);
   U251 : AOI222_X1 port map( A1 => n8, A2 => n2157, B1 => n2152, B2 => n709, 
                           C1 => n72, C2 => n2142, ZN => n708);
   U252 : OAI221_X1 port map( B1 => n2165, B2 => n710, C1 => n1892, C2 => n2163
                           , A => n711, ZN => n1636);
   U253 : AOI222_X1 port map( A1 => n7, A2 => n2157, B1 => n2152, B2 => n712, 
                           C1 => n71, C2 => n2142, ZN => n711);
   U254 : OAI221_X1 port map( B1 => n2165, B2 => n713, C1 => n1891, C2 => n2163
                           , A => n714, ZN => n1635);
   U255 : AOI222_X1 port map( A1 => n6, A2 => n2157, B1 => n2152, B2 => n715, 
                           C1 => n70, C2 => n2142, ZN => n714);
   U256 : OAI221_X1 port map( B1 => n2165, B2 => n719, C1 => n1889, C2 => n2163
                           , A => n720, ZN => n1633);
   U257 : AOI222_X1 port map( A1 => n4, A2 => n2157, B1 => n2152, B2 => n721, 
                           C1 => n68, C2 => n2142, ZN => n720);
   U258 : OAI221_X1 port map( B1 => n2165, B2 => n728, C1 => n1886, C2 => n2164
                           , A => n729, ZN => n1630);
   U259 : AOI222_X1 port map( A1 => n2158, A2 => n730, B1 => n2148, B2 => n731,
                           C1 => n65, C2 => n2142, ZN => n729);
   U260 : OAI221_X1 port map( B1 => n623, B2 => n2138, C1 => n1856, C2 => n2132
                           , A => n800, ZN => n1571);
   U261 : AOI222_X1 port map( A1 => n2126, A2 => n35, B1 => n2120, B2 => n625, 
                           C1 => n2114, C2 => n99, ZN => n800);
   U262 : OAI221_X1 port map( B1 => n626, B2 => n2138, C1 => n1855, C2 => n2132
                           , A => n802, ZN => n1569);
   U263 : AOI222_X1 port map( A1 => n2126, A2 => n34, B1 => n2120, B2 => n628, 
                           C1 => n2114, C2 => n98, ZN => n802);
   U264 : OAI221_X1 port map( B1 => n629, B2 => n2138, C1 => n1854, C2 => n2132
                           , A => n804, ZN => n1567);
   U265 : AOI222_X1 port map( A1 => n2126, A2 => n33, B1 => n2120, B2 => n631, 
                           C1 => n2114, C2 => n97, ZN => n804);
   U266 : OAI221_X1 port map( B1 => n632, B2 => n2138, C1 => n1853, C2 => n2132
                           , A => n806, ZN => n1565);
   U267 : AOI222_X1 port map( A1 => n2126, A2 => n32, B1 => n2120, B2 => n634, 
                           C1 => n2114, C2 => n96, ZN => n806);
   U268 : OAI221_X1 port map( B1 => n635, B2 => n2138, C1 => n1852, C2 => n2132
                           , A => n808, ZN => n1563);
   U269 : AOI222_X1 port map( A1 => n2126, A2 => n31, B1 => n2120, B2 => n637, 
                           C1 => n2114, C2 => n95, ZN => n808);
   U270 : OAI221_X1 port map( B1 => n638, B2 => n2138, C1 => n1851, C2 => n2132
                           , A => n810, ZN => n1561);
   U271 : AOI222_X1 port map( A1 => n2126, A2 => n30, B1 => n2120, B2 => n640, 
                           C1 => n2114, C2 => n94, ZN => n810);
   U272 : OAI221_X1 port map( B1 => n641, B2 => n2138, C1 => n1850, C2 => n2132
                           , A => n812, ZN => n1559);
   U273 : AOI222_X1 port map( A1 => n2126, A2 => n29, B1 => n2120, B2 => n643, 
                           C1 => n2114, C2 => n93, ZN => n812);
   U274 : OAI221_X1 port map( B1 => n644, B2 => n2138, C1 => n1849, C2 => n2133
                           , A => n814, ZN => n1557);
   U275 : AOI222_X1 port map( A1 => n2126, A2 => n28, B1 => n2120, B2 => n646, 
                           C1 => n2114, C2 => n92, ZN => n814);
   U276 : OAI221_X1 port map( B1 => n647, B2 => n2138, C1 => n1848, C2 => n2133
                           , A => n816, ZN => n1555);
   U277 : AOI222_X1 port map( A1 => n2126, A2 => n27, B1 => n2120, B2 => n649, 
                           C1 => n2114, C2 => n91, ZN => n816);
   U278 : OAI221_X1 port map( B1 => n650, B2 => n2138, C1 => n1847, C2 => n2133
                           , A => n818, ZN => n1553);
   U279 : AOI222_X1 port map( A1 => n2126, A2 => n26, B1 => n2120, B2 => n652, 
                           C1 => n2114, C2 => n90, ZN => n818);
   U280 : OAI221_X1 port map( B1 => n653, B2 => n2138, C1 => n1846, C2 => n2133
                           , A => n820, ZN => n1551);
   U281 : AOI222_X1 port map( A1 => n2126, A2 => n25, B1 => n2120, B2 => n655, 
                           C1 => n2114, C2 => n89, ZN => n820);
   U282 : OAI221_X1 port map( B1 => n656, B2 => n2137, C1 => n1845, C2 => n2133
                           , A => n822, ZN => n1549);
   U283 : AOI222_X1 port map( A1 => n2125, A2 => n24, B1 => n2119, B2 => n658, 
                           C1 => n2113, C2 => n88, ZN => n822);
   U284 : OAI221_X1 port map( B1 => n659, B2 => n2137, C1 => n1844, C2 => n2133
                           , A => n824, ZN => n1547);
   U285 : AOI222_X1 port map( A1 => n2125, A2 => n23, B1 => n2119, B2 => n661, 
                           C1 => n2113, C2 => n87, ZN => n824);
   U286 : OAI221_X1 port map( B1 => n662, B2 => n2137, C1 => n1843, C2 => n2133
                           , A => n826, ZN => n1545);
   U287 : AOI222_X1 port map( A1 => n2125, A2 => n22, B1 => n2119, B2 => n664, 
                           C1 => n2113, C2 => n86, ZN => n826);
   U288 : OAI221_X1 port map( B1 => n665, B2 => n2137, C1 => n1842, C2 => n2133
                           , A => n828, ZN => n1543);
   U289 : AOI222_X1 port map( A1 => n2125, A2 => n21, B1 => n2119, B2 => n667, 
                           C1 => n2113, C2 => n85, ZN => n828);
   U290 : OAI221_X1 port map( B1 => n668, B2 => n2137, C1 => n1841, C2 => n2133
                           , A => n830, ZN => n1541);
   U291 : AOI222_X1 port map( A1 => n2125, A2 => n20, B1 => n2119, B2 => n670, 
                           C1 => n2113, C2 => n84, ZN => n830);
   U292 : OAI221_X1 port map( B1 => n671, B2 => n2137, C1 => n1840, C2 => n2133
                           , A => n832, ZN => n1539);
   U293 : AOI222_X1 port map( A1 => n2125, A2 => n19, B1 => n2119, B2 => n673, 
                           C1 => n2113, C2 => n83, ZN => n832);
   U294 : OAI221_X1 port map( B1 => n674, B2 => n2137, C1 => n1839, C2 => n2133
                           , A => n834, ZN => n1537);
   U295 : AOI222_X1 port map( A1 => n2125, A2 => n18, B1 => n2119, B2 => n676, 
                           C1 => n2113, C2 => n82, ZN => n834);
   U296 : OAI221_X1 port map( B1 => n677, B2 => n2137, C1 => n1838, C2 => n2133
                           , A => n836, ZN => n1535);
   U297 : AOI222_X1 port map( A1 => n2125, A2 => n17, B1 => n2119, B2 => n679, 
                           C1 => n2113, C2 => n81, ZN => n836);
   U298 : OAI221_X1 port map( B1 => n680, B2 => n2137, C1 => n1837, C2 => n2134
                           , A => n838, ZN => n1533);
   U299 : AOI222_X1 port map( A1 => n2125, A2 => n16, B1 => n2119, B2 => n682, 
                           C1 => n2113, C2 => n80, ZN => n838);
   U300 : OAI221_X1 port map( B1 => n683, B2 => n2137, C1 => n1836, C2 => n2134
                           , A => n840, ZN => n1531);
   U301 : AOI222_X1 port map( A1 => n2125, A2 => n15, B1 => n2119, B2 => n685, 
                           C1 => n2113, C2 => n79, ZN => n840);
   U302 : OAI221_X1 port map( B1 => n686, B2 => n2137, C1 => n1835, C2 => n2134
                           , A => n842, ZN => n1529);
   U303 : AOI222_X1 port map( A1 => n2125, A2 => n14, B1 => n2119, B2 => n688, 
                           C1 => n2113, C2 => n78, ZN => n842);
   U304 : OAI221_X1 port map( B1 => n689, B2 => n2137, C1 => n1834, C2 => n2134
                           , A => n844, ZN => n1527);
   U305 : AOI222_X1 port map( A1 => n2125, A2 => n13, B1 => n2119, B2 => n691, 
                           C1 => n2113, C2 => n77, ZN => n844);
   U306 : OAI221_X1 port map( B1 => n692, B2 => n2136, C1 => n1833, C2 => n2134
                           , A => n846, ZN => n1525);
   U307 : AOI222_X1 port map( A1 => n2124, A2 => n694, B1 => n2118, B2 => n695,
                           C1 => n2112, C2 => n76, ZN => n846);
   U308 : OAI221_X1 port map( B1 => n696, B2 => n2136, C1 => n1832, C2 => n2134
                           , A => n848, ZN => n1523);
   U309 : AOI222_X1 port map( A1 => n2124, A2 => n698, B1 => n2118, B2 => n699,
                           C1 => n2112, C2 => n75, ZN => n848);
   U310 : OAI221_X1 port map( B1 => n700, B2 => n2136, C1 => n1831, C2 => n2134
                           , A => n850, ZN => n1521);
   U311 : AOI222_X1 port map( A1 => n2124, A2 => n702, B1 => n2118, B2 => n703,
                           C1 => n2112, C2 => n74, ZN => n850);
   U312 : OAI221_X1 port map( B1 => n704, B2 => n2136, C1 => n1830, C2 => n2134
                           , A => n852, ZN => n1519);
   U313 : AOI222_X1 port map( A1 => n2124, A2 => n9, B1 => n2118, B2 => n706, 
                           C1 => n2112, C2 => n73, ZN => n852);
   U314 : OAI221_X1 port map( B1 => n707, B2 => n2136, C1 => n1829, C2 => n2134
                           , A => n854, ZN => n1517);
   U315 : AOI222_X1 port map( A1 => n2124, A2 => n8, B1 => n2118, B2 => n709, 
                           C1 => n2112, C2 => n72, ZN => n854);
   U316 : OAI221_X1 port map( B1 => n710, B2 => n2136, C1 => n1828, C2 => n2134
                           , A => n856, ZN => n1515);
   U317 : AOI222_X1 port map( A1 => n2124, A2 => n7, B1 => n2118, B2 => n712, 
                           C1 => n2112, C2 => n71, ZN => n856);
   U318 : OAI221_X1 port map( B1 => n713, B2 => n2136, C1 => n1827, C2 => n2134
                           , A => n858, ZN => n1513);
   U319 : AOI222_X1 port map( A1 => n2124, A2 => n6, B1 => n2118, B2 => n715, 
                           C1 => n2112, C2 => n70, ZN => n858);
   U320 : OAI221_X1 port map( B1 => n716, B2 => n2136, C1 => n1826, C2 => n2135
                           , A => n860, ZN => n1511);
   U321 : AOI222_X1 port map( A1 => n2124, A2 => n5, B1 => n2118, B2 => n718, 
                           C1 => n2112, C2 => n69, ZN => n860);
   U322 : OAI221_X1 port map( B1 => n719, B2 => n2136, C1 => n1825, C2 => n2134
                           , A => n862, ZN => n1509);
   U323 : AOI222_X1 port map( A1 => n2124, A2 => n4, B1 => n2118, B2 => n721, 
                           C1 => n2112, C2 => n68, ZN => n862);
   U324 : OAI221_X1 port map( B1 => n722, B2 => n2136, C1 => n1824, C2 => n2135
                           , A => n864, ZN => n1507);
   U325 : AOI222_X1 port map( A1 => n2124, A2 => n3, B1 => n2118, B2 => n724, 
                           C1 => n2112, C2 => n67, ZN => n864);
   U326 : OAI221_X1 port map( B1 => n725, B2 => n2136, C1 => n1823, C2 => n2135
                           , A => n866, ZN => n1505);
   U327 : AOI222_X1 port map( A1 => n2124, A2 => n2, B1 => n2118, B2 => n727, 
                           C1 => n2112, C2 => n66, ZN => n866);
   U328 : OAI221_X1 port map( B1 => n728, B2 => n2136, C1 => n1822, C2 => n2135
                           , A => n868, ZN => n1503);
   U329 : AOI222_X1 port map( A1 => n2124, A2 => n730, B1 => n2118, B2 => n731,
                           C1 => n2112, C2 => n65, ZN => n868);
   U330 : INV_X1 port map( A => RESET, ZN => n734);
   U331 : OAI221_X1 port map( B1 => n2170, B2 => n522, C1 => n1949, C2 => n2159
                           , A => n524, ZN => n1693);
   U332 : AOI222_X1 port map( A1 => n64, A2 => n2155, B1 => n192, B2 => n2148, 
                           C1 => n2147, C2 => n528, ZN => n524);
   U333 : OAI221_X1 port map( B1 => n2170, B2 => n529, C1 => n1948, C2 => n2159
                           , A => n530, ZN => n1692);
   U334 : AOI222_X1 port map( A1 => n63, A2 => n2153, B1 => n191, B2 => n2148, 
                           C1 => n2147, C2 => n531, ZN => n530);
   U335 : OAI221_X1 port map( B1 => n2170, B2 => n532, C1 => n1947, C2 => n2159
                           , A => n533, ZN => n1691);
   U336 : AOI222_X1 port map( A1 => n62, A2 => n2153, B1 => n190, B2 => n2148, 
                           C1 => n2146, C2 => n534, ZN => n533);
   U337 : OAI221_X1 port map( B1 => n2170, B2 => n535, C1 => n1946, C2 => n2159
                           , A => n536, ZN => n1690);
   U338 : AOI222_X1 port map( A1 => n61, A2 => n2153, B1 => n189, B2 => n2148, 
                           C1 => n2146, C2 => n537, ZN => n536);
   U339 : OAI221_X1 port map( B1 => n2167, B2 => n619, C1 => n1921, C2 => n2161
                           , A => n620, ZN => n1665);
   U340 : AOI222_X1 port map( A1 => n36, A2 => n2155, B1 => n2150, B2 => n621, 
                           C1 => n2144, C2 => n622, ZN => n620);
   U341 : OAI221_X1 port map( B1 => n2167, B2 => n623, C1 => n1920, C2 => n2161
                           , A => n624, ZN => n1664);
   U342 : AOI222_X1 port map( A1 => n35, A2 => n2155, B1 => n2150, B2 => n625, 
                           C1 => n99, C2 => n2144, ZN => n624);
   U343 : OAI221_X1 port map( B1 => n2167, B2 => n626, C1 => n1919, C2 => n2161
                           , A => n627, ZN => n1663);
   U344 : AOI222_X1 port map( A1 => n34, A2 => n2155, B1 => n2150, B2 => n628, 
                           C1 => n98, C2 => n2144, ZN => n627);
   U345 : OAI221_X1 port map( B1 => n2167, B2 => n629, C1 => n1918, C2 => n2161
                           , A => n630, ZN => n1662);
   U346 : AOI222_X1 port map( A1 => n33, A2 => n2155, B1 => n2150, B2 => n631, 
                           C1 => n97, C2 => n2144, ZN => n630);
   U347 : OAI221_X1 port map( B1 => n2167, B2 => n632, C1 => n1917, C2 => n2161
                           , A => n633, ZN => n1661);
   U348 : AOI222_X1 port map( A1 => n32, A2 => n2155, B1 => n2150, B2 => n634, 
                           C1 => n96, C2 => n2144, ZN => n633);
   U349 : OAI221_X1 port map( B1 => n2167, B2 => n635, C1 => n1916, C2 => n2161
                           , A => n636, ZN => n1660);
   U350 : AOI222_X1 port map( A1 => n31, A2 => n2155, B1 => n2150, B2 => n637, 
                           C1 => n95, C2 => n2144, ZN => n636);
   U351 : OAI221_X1 port map( B1 => n2167, B2 => n638, C1 => n1915, C2 => n2161
                           , A => n639, ZN => n1659);
   U352 : AOI222_X1 port map( A1 => n30, A2 => n2155, B1 => n2150, B2 => n640, 
                           C1 => n94, C2 => n2144, ZN => n639);
   U353 : OAI221_X1 port map( B1 => n2167, B2 => n641, C1 => n1914, C2 => n2161
                           , A => n642, ZN => n1658);
   U354 : AOI222_X1 port map( A1 => n29, A2 => n2155, B1 => n2150, B2 => n643, 
                           C1 => n93, C2 => n2144, ZN => n642);
   U355 : OAI221_X1 port map( B1 => n2167, B2 => n644, C1 => n1913, C2 => n2162
                           , A => n645, ZN => n1657);
   U356 : AOI222_X1 port map( A1 => n28, A2 => n2156, B1 => n2150, B2 => n646, 
                           C1 => n92, C2 => n2144, ZN => n645);
   U357 : OAI221_X1 port map( B1 => n2167, B2 => n647, C1 => n1912, C2 => n2162
                           , A => n648, ZN => n1656);
   U358 : AOI222_X1 port map( A1 => n27, A2 => n2156, B1 => n2151, B2 => n649, 
                           C1 => n91, C2 => n2144, ZN => n648);
   U359 : OAI221_X1 port map( B1 => n2167, B2 => n650, C1 => n1911, C2 => n2162
                           , A => n651, ZN => n1655);
   U360 : AOI222_X1 port map( A1 => n26, A2 => n2156, B1 => n2151, B2 => n652, 
                           C1 => n90, C2 => n2144, ZN => n651);
   U361 : OAI221_X1 port map( B1 => n2167, B2 => n653, C1 => n1910, C2 => n2162
                           , A => n654, ZN => n1654);
   U362 : AOI222_X1 port map( A1 => n25, A2 => n2156, B1 => n2151, B2 => n655, 
                           C1 => n89, C2 => n2144, ZN => n654);
   U363 : OAI221_X1 port map( B1 => n2165, B2 => n716, C1 => n1890, C2 => n2164
                           , A => n717, ZN => n1634);
   U364 : AOI222_X1 port map( A1 => n5, A2 => n2157, B1 => n2152, B2 => n718, 
                           C1 => n69, C2 => n2142, ZN => n717);
   U365 : OAI221_X1 port map( B1 => n2165, B2 => n722, C1 => n1888, C2 => n2164
                           , A => n723, ZN => n1632);
   U366 : AOI222_X1 port map( A1 => n3, A2 => n2157, B1 => n2152, B2 => n724, 
                           C1 => n67, C2 => n2142, ZN => n723);
   U367 : OAI221_X1 port map( B1 => n2165, B2 => n725, C1 => n1887, C2 => n2164
                           , A => n726, ZN => n1631);
   U368 : AOI222_X1 port map( A1 => n2, A2 => n2157, B1 => n2152, B2 => n727, 
                           C1 => n66, C2 => n2142, ZN => n726);
   U369 : OAI221_X1 port map( B1 => n522, B2 => n2141, C1 => n1885, C2 => n2130
                           , A => n737, ZN => n1629);
   U370 : AOI222_X1 port map( A1 => n2129, A2 => n64, B1 => n2123, B2 => n192, 
                           C1 => n2117, C2 => n528, ZN => n737);
   U371 : OAI221_X1 port map( B1 => n529, B2 => n2141, C1 => n1884, C2 => n2130
                           , A => n744, ZN => n1627);
   U372 : AOI222_X1 port map( A1 => n2129, A2 => n63, B1 => n2123, B2 => n191, 
                           C1 => n2117, C2 => n531, ZN => n744);
   U373 : OAI221_X1 port map( B1 => n532, B2 => n2141, C1 => n1883, C2 => n2130
                           , A => n746, ZN => n1625);
   U374 : AOI222_X1 port map( A1 => n2129, A2 => n62, B1 => n2123, B2 => n190, 
                           C1 => n2117, C2 => n534, ZN => n746);
   U375 : OAI221_X1 port map( B1 => n535, B2 => n2141, C1 => n1882, C2 => n2130
                           , A => n748, ZN => n1623);
   U376 : AOI222_X1 port map( A1 => n2129, A2 => n61, B1 => n2123, B2 => n189, 
                           C1 => n2117, C2 => n537, ZN => n748);
   U377 : OAI221_X1 port map( B1 => n583, B2 => n2139, C1 => n1866, C2 => n2131
                           , A => n780, ZN => n1591);
   U378 : AOI222_X1 port map( A1 => n2127, A2 => n45, B1 => n2121, B2 => n585, 
                           C1 => n2115, C2 => n586, ZN => n780);
   U379 : OAI221_X1 port map( B1 => n587, B2 => n2139, C1 => n1865, C2 => n2131
                           , A => n782, ZN => n1589);
   U380 : AOI222_X1 port map( A1 => n2127, A2 => n44, B1 => n2121, B2 => n589, 
                           C1 => n2115, C2 => n590, ZN => n782);
   U381 : OAI221_X1 port map( B1 => n591, B2 => n2139, C1 => n1864, C2 => n2131
                           , A => n784, ZN => n1587);
   U382 : AOI222_X1 port map( A1 => n2127, A2 => n43, B1 => n2121, B2 => n593, 
                           C1 => n2115, C2 => n594, ZN => n784);
   U383 : OAI221_X1 port map( B1 => n595, B2 => n2139, C1 => n1863, C2 => n2131
                           , A => n786, ZN => n1585);
   U384 : AOI222_X1 port map( A1 => n2127, A2 => n42, B1 => n2121, B2 => n597, 
                           C1 => n2115, C2 => n598, ZN => n786);
   U385 : OAI221_X1 port map( B1 => n599, B2 => n2139, C1 => n1862, C2 => n2131
                           , A => n788, ZN => n1583);
   U386 : AOI222_X1 port map( A1 => n2127, A2 => n41, B1 => n2121, B2 => n601, 
                           C1 => n2115, C2 => n602, ZN => n788);
   U387 : OAI221_X1 port map( B1 => n603, B2 => n2139, C1 => n1861, C2 => n2131
                           , A => n790, ZN => n1581);
   U388 : AOI222_X1 port map( A1 => n2127, A2 => n40, B1 => n2121, B2 => n605, 
                           C1 => n2115, C2 => n606, ZN => n790);
   U389 : OAI221_X1 port map( B1 => n607, B2 => n2139, C1 => n1860, C2 => n2132
                           , A => n792, ZN => n1579);
   U390 : AOI222_X1 port map( A1 => n2127, A2 => n39, B1 => n2121, B2 => n609, 
                           C1 => n2115, C2 => n610, ZN => n792);
   U391 : OAI221_X1 port map( B1 => n611, B2 => n2139, C1 => n1859, C2 => n2132
                           , A => n794, ZN => n1577);
   U392 : AOI222_X1 port map( A1 => n2127, A2 => n38, B1 => n2121, B2 => n613, 
                           C1 => n2115, C2 => n614, ZN => n794);
   U393 : OAI221_X1 port map( B1 => n615, B2 => n2139, C1 => n1858, C2 => n2132
                           , A => n796, ZN => n1575);
   U394 : AOI222_X1 port map( A1 => n2127, A2 => n37, B1 => n2121, B2 => n617, 
                           C1 => n2115, C2 => n618, ZN => n796);
   U395 : OAI221_X1 port map( B1 => n619, B2 => n2138, C1 => n1857, C2 => n2132
                           , A => n798, ZN => n1573);
   U396 : AOI222_X1 port map( A1 => n2126, A2 => n36, B1 => n2120, B2 => n621, 
                           C1 => n2114, C2 => n622, ZN => n798);
   U397 : OAI221_X1 port map( B1 => n2169, B2 => n538, C1 => n1945, C2 => n2159
                           , A => n539, ZN => n1689);
   U398 : AOI222_X1 port map( A1 => n60, A2 => n2153, B1 => n188, B2 => n2148, 
                           C1 => n2146, C2 => n540, ZN => n539);
   U399 : OAI221_X1 port map( B1 => n2169, B2 => n541, C1 => n1944, C2 => n2159
                           , A => n542, ZN => n1688);
   U400 : AOI222_X1 port map( A1 => n59, A2 => n2153, B1 => n187, B2 => n2148, 
                           C1 => n2146, C2 => n543, ZN => n542);
   U401 : OAI221_X1 port map( B1 => n2169, B2 => n544, C1 => n1943, C2 => n2159
                           , A => n545, ZN => n1687);
   U402 : AOI222_X1 port map( A1 => n58, A2 => n2153, B1 => n186, B2 => n2148, 
                           C1 => n2146, C2 => n546, ZN => n545);
   U403 : OAI221_X1 port map( B1 => n2169, B2 => n547, C1 => n1942, C2 => n2159
                           , A => n548, ZN => n1686);
   U404 : AOI222_X1 port map( A1 => n57, A2 => n2153, B1 => n185, B2 => n2148, 
                           C1 => n2146, C2 => n549, ZN => n548);
   U405 : OAI221_X1 port map( B1 => n2169, B2 => n550, C1 => n1941, C2 => n2159
                           , A => n551, ZN => n1685);
   U406 : AOI222_X1 port map( A1 => n56, A2 => n2153, B1 => n184, B2 => n2148, 
                           C1 => n2146, C2 => n552, ZN => n551);
   U407 : OAI221_X1 port map( B1 => n2169, B2 => n553, C1 => n1940, C2 => n2159
                           , A => n554, ZN => n1684);
   U408 : AOI222_X1 port map( A1 => n55, A2 => n2153, B1 => n183, B2 => n2148, 
                           C1 => n2146, C2 => n555, ZN => n554);
   U409 : OAI221_X1 port map( B1 => n2169, B2 => n556, C1 => n1939, C2 => n2159
                           , A => n557, ZN => n1683);
   U410 : AOI222_X1 port map( A1 => n54, A2 => n2153, B1 => n182, B2 => n2148, 
                           C1 => n2146, C2 => n558, ZN => n557);
   U411 : OAI221_X1 port map( B1 => n2169, B2 => n559, C1 => n1938, C2 => n2159
                           , A => n560, ZN => n1682);
   U412 : AOI222_X1 port map( A1 => n53, A2 => n2153, B1 => n181, B2 => n2148, 
                           C1 => n2146, C2 => n561, ZN => n560);
   U413 : OAI221_X1 port map( B1 => n2168, B2 => n583, C1 => n1930, C2 => n2160
                           , A => n584, ZN => n1674);
   U414 : AOI222_X1 port map( A1 => n45, A2 => n2154, B1 => n2149, B2 => n585, 
                           C1 => n2145, C2 => n586, ZN => n584);
   U415 : OAI221_X1 port map( B1 => n2168, B2 => n587, C1 => n1929, C2 => n2160
                           , A => n588, ZN => n1673);
   U416 : AOI222_X1 port map( A1 => n44, A2 => n2154, B1 => n2149, B2 => n589, 
                           C1 => n2145, C2 => n590, ZN => n588);
   U417 : OAI221_X1 port map( B1 => n2168, B2 => n591, C1 => n1928, C2 => n2160
                           , A => n592, ZN => n1672);
   U418 : AOI222_X1 port map( A1 => n43, A2 => n2154, B1 => n2149, B2 => n593, 
                           C1 => n2145, C2 => n594, ZN => n592);
   U419 : OAI221_X1 port map( B1 => n2168, B2 => n595, C1 => n1927, C2 => n2160
                           , A => n596, ZN => n1671);
   U420 : AOI222_X1 port map( A1 => n42, A2 => n2154, B1 => n2149, B2 => n597, 
                           C1 => n2145, C2 => n598, ZN => n596);
   U421 : OAI221_X1 port map( B1 => n2168, B2 => n599, C1 => n1926, C2 => n2160
                           , A => n600, ZN => n1670);
   U422 : AOI222_X1 port map( A1 => n41, A2 => n2154, B1 => n2149, B2 => n601, 
                           C1 => n2145, C2 => n602, ZN => n600);
   U423 : OAI221_X1 port map( B1 => n2168, B2 => n603, C1 => n1925, C2 => n2160
                           , A => n604, ZN => n1669);
   U424 : AOI222_X1 port map( A1 => n40, A2 => n2154, B1 => n2150, B2 => n605, 
                           C1 => n2145, C2 => n606, ZN => n604);
   U425 : OAI221_X1 port map( B1 => n2168, B2 => n607, C1 => n1924, C2 => n2161
                           , A => n608, ZN => n1668);
   U426 : AOI222_X1 port map( A1 => n39, A2 => n2155, B1 => n2150, B2 => n609, 
                           C1 => n2145, C2 => n610, ZN => n608);
   U427 : OAI221_X1 port map( B1 => n2168, B2 => n611, C1 => n1923, C2 => n2161
                           , A => n612, ZN => n1667);
   U428 : AOI222_X1 port map( A1 => n38, A2 => n2155, B1 => n2150, B2 => n613, 
                           C1 => n2145, C2 => n614, ZN => n612);
   U429 : OAI221_X1 port map( B1 => n2168, B2 => n615, C1 => n1922, C2 => n2161
                           , A => n616, ZN => n1666);
   U430 : AOI222_X1 port map( A1 => n37, A2 => n2155, B1 => n2150, B2 => n617, 
                           C1 => n2145, C2 => n618, ZN => n616);
   U431 : OAI22_X1 port map( A1 => n1950, A2 => n2099, B1 => n743, B2 => n2093,
                           ZN => n1501);
   U432 : OAI22_X1 port map( A1 => n1951, A2 => n2099, B1 => n745, B2 => n2093,
                           ZN => n1500);
   U433 : OAI22_X1 port map( A1 => n1952, A2 => n2099, B1 => n747, B2 => n2093,
                           ZN => n1499);
   U434 : OAI22_X1 port map( A1 => n1953, A2 => n2099, B1 => n749, B2 => n2093,
                           ZN => n1498);
   U435 : OAI22_X1 port map( A1 => n1821, A2 => n2087, B1 => n743, B2 => n2081,
                           ZN => n1437);
   U436 : OAI22_X1 port map( A1 => n1820, A2 => n2087, B1 => n745, B2 => n2081,
                           ZN => n1436);
   U437 : OAI22_X1 port map( A1 => n1819, A2 => n2087, B1 => n747, B2 => n2081,
                           ZN => n1435);
   U438 : OAI22_X1 port map( A1 => n1818, A2 => n2087, B1 => n749, B2 => n2081,
                           ZN => n1434);
   U439 : OAI22_X1 port map( A1 => n2010, A2 => n2075, B1 => n743, B2 => n2069,
                           ZN => n1373);
   U440 : OAI22_X1 port map( A1 => n2011, A2 => n2075, B1 => n745, B2 => n2069,
                           ZN => n1372);
   U441 : OAI22_X1 port map( A1 => n2012, A2 => n2075, B1 => n747, B2 => n2069,
                           ZN => n1371);
   U442 : OAI22_X1 port map( A1 => n2013, A2 => n2075, B1 => n749, B2 => n2069,
                           ZN => n1370);
   U443 : OAI22_X1 port map( A1 => n1954, A2 => n2099, B1 => n751, B2 => n2092,
                           ZN => n1497);
   U444 : OAI22_X1 port map( A1 => n1955, A2 => n2098, B1 => n753, B2 => n2092,
                           ZN => n1496);
   U445 : OAI22_X1 port map( A1 => n1956, A2 => n2098, B1 => n755, B2 => n2092,
                           ZN => n1495);
   U446 : OAI22_X1 port map( A1 => n1957, A2 => n2098, B1 => n757, B2 => n2092,
                           ZN => n1494);
   U447 : OAI22_X1 port map( A1 => n1958, A2 => n2098, B1 => n759, B2 => n2092,
                           ZN => n1493);
   U448 : OAI22_X1 port map( A1 => n1959, A2 => n2098, B1 => n761, B2 => n2092,
                           ZN => n1492);
   U449 : OAI22_X1 port map( A1 => n1960, A2 => n2098, B1 => n763, B2 => n2092,
                           ZN => n1491);
   U450 : OAI22_X1 port map( A1 => n1961, A2 => n2098, B1 => n765, B2 => n2092,
                           ZN => n1490);
   U451 : OAI22_X1 port map( A1 => n1962, A2 => n2098, B1 => n767, B2 => n2092,
                           ZN => n1489);
   U452 : OAI22_X1 port map( A1 => n1963, A2 => n2098, B1 => n769, B2 => n2092,
                           ZN => n1488);
   U453 : OAI22_X1 port map( A1 => n1964, A2 => n2098, B1 => n771, B2 => n2092,
                           ZN => n1487);
   U454 : OAI22_X1 port map( A1 => n1965, A2 => n2098, B1 => n773, B2 => n2092,
                           ZN => n1486);
   U455 : OAI22_X1 port map( A1 => n1966, A2 => n2098, B1 => n775, B2 => n2091,
                           ZN => n1485);
   U456 : OAI22_X1 port map( A1 => n1967, A2 => n2097, B1 => n777, B2 => n2091,
                           ZN => n1484);
   U457 : OAI22_X1 port map( A1 => n1968, A2 => n2097, B1 => n779, B2 => n2091,
                           ZN => n1483);
   U458 : OAI22_X1 port map( A1 => n1969, A2 => n2097, B1 => n781, B2 => n2091,
                           ZN => n1482);
   U459 : OAI22_X1 port map( A1 => n1970, A2 => n2097, B1 => n783, B2 => n2091,
                           ZN => n1481);
   U460 : OAI22_X1 port map( A1 => n1971, A2 => n2097, B1 => n785, B2 => n2091,
                           ZN => n1480);
   U461 : OAI22_X1 port map( A1 => n1972, A2 => n2097, B1 => n787, B2 => n2091,
                           ZN => n1479);
   U462 : OAI22_X1 port map( A1 => n1973, A2 => n2097, B1 => n789, B2 => n2091,
                           ZN => n1478);
   U463 : OAI22_X1 port map( A1 => n1974, A2 => n2097, B1 => n791, B2 => n2091,
                           ZN => n1477);
   U464 : OAI22_X1 port map( A1 => n1975, A2 => n2097, B1 => n793, B2 => n2091,
                           ZN => n1476);
   U465 : OAI22_X1 port map( A1 => n1976, A2 => n2097, B1 => n795, B2 => n2091,
                           ZN => n1475);
   U466 : OAI22_X1 port map( A1 => n1977, A2 => n2097, B1 => n797, B2 => n2091,
                           ZN => n1474);
   U467 : OAI22_X1 port map( A1 => n1978, A2 => n2097, B1 => n799, B2 => n2090,
                           ZN => n1473);
   U468 : OAI22_X1 port map( A1 => n1979, A2 => n2096, B1 => n801, B2 => n2090,
                           ZN => n1472);
   U469 : OAI22_X1 port map( A1 => n1980, A2 => n2096, B1 => n803, B2 => n2090,
                           ZN => n1471);
   U470 : OAI22_X1 port map( A1 => n1981, A2 => n2096, B1 => n805, B2 => n2090,
                           ZN => n1470);
   U471 : OAI22_X1 port map( A1 => n1982, A2 => n2096, B1 => n807, B2 => n2090,
                           ZN => n1469);
   U472 : OAI22_X1 port map( A1 => n1983, A2 => n2096, B1 => n809, B2 => n2090,
                           ZN => n1468);
   U473 : OAI22_X1 port map( A1 => n1984, A2 => n2096, B1 => n811, B2 => n2090,
                           ZN => n1467);
   U474 : OAI22_X1 port map( A1 => n1985, A2 => n2096, B1 => n813, B2 => n2090,
                           ZN => n1466);
   U475 : OAI22_X1 port map( A1 => n1986, A2 => n2096, B1 => n815, B2 => n2090,
                           ZN => n1465);
   U476 : OAI22_X1 port map( A1 => n1987, A2 => n2096, B1 => n817, B2 => n2090,
                           ZN => n1464);
   U477 : OAI22_X1 port map( A1 => n1988, A2 => n2096, B1 => n819, B2 => n2090,
                           ZN => n1463);
   U478 : OAI22_X1 port map( A1 => n1989, A2 => n2096, B1 => n821, B2 => n2090,
                           ZN => n1462);
   U479 : OAI22_X1 port map( A1 => n1990, A2 => n2096, B1 => n823, B2 => n2089,
                           ZN => n1461);
   U480 : OAI22_X1 port map( A1 => n1991, A2 => n2095, B1 => n825, B2 => n2089,
                           ZN => n1460);
   U481 : OAI22_X1 port map( A1 => n1992, A2 => n2095, B1 => n827, B2 => n2089,
                           ZN => n1459);
   U482 : OAI22_X1 port map( A1 => n1993, A2 => n2095, B1 => n829, B2 => n2089,
                           ZN => n1458);
   U483 : OAI22_X1 port map( A1 => n1994, A2 => n2095, B1 => n831, B2 => n2089,
                           ZN => n1457);
   U484 : OAI22_X1 port map( A1 => n1995, A2 => n2095, B1 => n833, B2 => n2089,
                           ZN => n1456);
   U485 : OAI22_X1 port map( A1 => n1996, A2 => n2095, B1 => n835, B2 => n2089,
                           ZN => n1455);
   U486 : OAI22_X1 port map( A1 => n1997, A2 => n2095, B1 => n837, B2 => n2089,
                           ZN => n1454);
   U487 : OAI22_X1 port map( A1 => n1998, A2 => n2095, B1 => n839, B2 => n2089,
                           ZN => n1453);
   U488 : OAI22_X1 port map( A1 => n1999, A2 => n2095, B1 => n841, B2 => n2089,
                           ZN => n1452);
   U489 : OAI22_X1 port map( A1 => n2000, A2 => n2095, B1 => n843, B2 => n2089,
                           ZN => n1451);
   U490 : OAI22_X1 port map( A1 => n2001, A2 => n2095, B1 => n845, B2 => n2089,
                           ZN => n1450);
   U491 : OAI22_X1 port map( A1 => n1204, A2 => n2095, B1 => n847, B2 => n2088,
                           ZN => n1449);
   U492 : OAI22_X1 port map( A1 => n1202, A2 => n2094, B1 => n849, B2 => n2088,
                           ZN => n1448);
   U493 : OAI22_X1 port map( A1 => n1200, A2 => n2094, B1 => n851, B2 => n2088,
                           ZN => n1447);
   U494 : OAI22_X1 port map( A1 => n2002, A2 => n2094, B1 => n853, B2 => n2088,
                           ZN => n1446);
   U495 : OAI22_X1 port map( A1 => n2003, A2 => n2094, B1 => n855, B2 => n2088,
                           ZN => n1445);
   U496 : OAI22_X1 port map( A1 => n2004, A2 => n2094, B1 => n857, B2 => n2088,
                           ZN => n1444);
   U497 : OAI22_X1 port map( A1 => n2005, A2 => n2094, B1 => n859, B2 => n2088,
                           ZN => n1443);
   U498 : OAI22_X1 port map( A1 => n2006, A2 => n2094, B1 => n861, B2 => n2088,
                           ZN => n1442);
   U499 : OAI22_X1 port map( A1 => n2007, A2 => n2094, B1 => n863, B2 => n2088,
                           ZN => n1441);
   U500 : OAI22_X1 port map( A1 => n2008, A2 => n2094, B1 => n865, B2 => n2088,
                           ZN => n1440);
   U501 : OAI22_X1 port map( A1 => n2009, A2 => n2094, B1 => n867, B2 => n2088,
                           ZN => n1439);
   U502 : OAI22_X1 port map( A1 => n415, A2 => n2094, B1 => n871, B2 => n2088, 
                           ZN => n1438);
   U503 : OAI22_X1 port map( A1 => n1817, A2 => n2087, B1 => n751, B2 => n2080,
                           ZN => n1433);
   U504 : OAI22_X1 port map( A1 => n1816, A2 => n2086, B1 => n753, B2 => n2080,
                           ZN => n1432);
   U505 : OAI22_X1 port map( A1 => n1815, A2 => n2086, B1 => n755, B2 => n2080,
                           ZN => n1431);
   U506 : OAI22_X1 port map( A1 => n1814, A2 => n2086, B1 => n757, B2 => n2080,
                           ZN => n1430);
   U507 : OAI22_X1 port map( A1 => n1813, A2 => n2086, B1 => n759, B2 => n2080,
                           ZN => n1429);
   U508 : OAI22_X1 port map( A1 => n1812, A2 => n2086, B1 => n761, B2 => n2080,
                           ZN => n1428);
   U509 : OAI22_X1 port map( A1 => n1811, A2 => n2086, B1 => n763, B2 => n2080,
                           ZN => n1427);
   U510 : OAI22_X1 port map( A1 => n1810, A2 => n2086, B1 => n765, B2 => n2080,
                           ZN => n1426);
   U511 : OAI22_X1 port map( A1 => n1809, A2 => n2086, B1 => n767, B2 => n2080,
                           ZN => n1425);
   U512 : OAI22_X1 port map( A1 => n1808, A2 => n2086, B1 => n769, B2 => n2080,
                           ZN => n1424);
   U513 : OAI22_X1 port map( A1 => n1807, A2 => n2086, B1 => n771, B2 => n2080,
                           ZN => n1423);
   U514 : OAI22_X1 port map( A1 => n1806, A2 => n2086, B1 => n773, B2 => n2080,
                           ZN => n1422);
   U515 : OAI22_X1 port map( A1 => n1805, A2 => n2086, B1 => n775, B2 => n2079,
                           ZN => n1421);
   U516 : OAI22_X1 port map( A1 => n1804, A2 => n2085, B1 => n777, B2 => n2079,
                           ZN => n1420);
   U517 : OAI22_X1 port map( A1 => n1803, A2 => n2085, B1 => n779, B2 => n2079,
                           ZN => n1419);
   U518 : OAI22_X1 port map( A1 => n1802, A2 => n2085, B1 => n781, B2 => n2079,
                           ZN => n1418);
   U519 : OAI22_X1 port map( A1 => n1801, A2 => n2085, B1 => n783, B2 => n2079,
                           ZN => n1417);
   U520 : OAI22_X1 port map( A1 => n1800, A2 => n2085, B1 => n785, B2 => n2079,
                           ZN => n1416);
   U521 : OAI22_X1 port map( A1 => n1799, A2 => n2085, B1 => n787, B2 => n2079,
                           ZN => n1415);
   U522 : OAI22_X1 port map( A1 => n1798, A2 => n2085, B1 => n789, B2 => n2079,
                           ZN => n1414);
   U523 : OAI22_X1 port map( A1 => n1797, A2 => n2085, B1 => n791, B2 => n2079,
                           ZN => n1413);
   U524 : OAI22_X1 port map( A1 => n1796, A2 => n2085, B1 => n793, B2 => n2079,
                           ZN => n1412);
   U525 : OAI22_X1 port map( A1 => n1795, A2 => n2085, B1 => n795, B2 => n2079,
                           ZN => n1411);
   U526 : OAI22_X1 port map( A1 => n1794, A2 => n2085, B1 => n797, B2 => n2079,
                           ZN => n1410);
   U527 : OAI22_X1 port map( A1 => n1793, A2 => n2085, B1 => n799, B2 => n2078,
                           ZN => n1409);
   U528 : OAI22_X1 port map( A1 => n2029, A2 => n2084, B1 => n801, B2 => n2078,
                           ZN => n1408);
   U529 : OAI22_X1 port map( A1 => n2030, A2 => n2084, B1 => n803, B2 => n2078,
                           ZN => n1407);
   U530 : OAI22_X1 port map( A1 => n2031, A2 => n2084, B1 => n805, B2 => n2078,
                           ZN => n1406);
   U531 : OAI22_X1 port map( A1 => n2032, A2 => n2084, B1 => n807, B2 => n2078,
                           ZN => n1405);
   U532 : OAI22_X1 port map( A1 => n2033, A2 => n2084, B1 => n809, B2 => n2078,
                           ZN => n1404);
   U533 : OAI22_X1 port map( A1 => n2034, A2 => n2084, B1 => n811, B2 => n2078,
                           ZN => n1403);
   U534 : OAI22_X1 port map( A1 => n2035, A2 => n2084, B1 => n813, B2 => n2078,
                           ZN => n1402);
   U535 : OAI22_X1 port map( A1 => n2036, A2 => n2084, B1 => n815, B2 => n2078,
                           ZN => n1401);
   U536 : OAI22_X1 port map( A1 => n2037, A2 => n2084, B1 => n817, B2 => n2078,
                           ZN => n1400);
   U537 : OAI22_X1 port map( A1 => n2038, A2 => n2084, B1 => n819, B2 => n2078,
                           ZN => n1399);
   U538 : OAI22_X1 port map( A1 => n2039, A2 => n2084, B1 => n821, B2 => n2078,
                           ZN => n1398);
   U539 : OAI22_X1 port map( A1 => n2040, A2 => n2084, B1 => n823, B2 => n2077,
                           ZN => n1397);
   U540 : OAI22_X1 port map( A1 => n2041, A2 => n2083, B1 => n825, B2 => n2077,
                           ZN => n1396);
   U541 : OAI22_X1 port map( A1 => n2042, A2 => n2083, B1 => n827, B2 => n2077,
                           ZN => n1395);
   U542 : OAI22_X1 port map( A1 => n2043, A2 => n2083, B1 => n829, B2 => n2077,
                           ZN => n1394);
   U543 : OAI22_X1 port map( A1 => n2044, A2 => n2083, B1 => n831, B2 => n2077,
                           ZN => n1393);
   U544 : OAI22_X1 port map( A1 => n2045, A2 => n2083, B1 => n833, B2 => n2077,
                           ZN => n1392);
   U545 : OAI22_X1 port map( A1 => n2046, A2 => n2083, B1 => n835, B2 => n2077,
                           ZN => n1391);
   U546 : OAI22_X1 port map( A1 => n2047, A2 => n2083, B1 => n837, B2 => n2077,
                           ZN => n1390);
   U547 : OAI22_X1 port map( A1 => n2048, A2 => n2083, B1 => n839, B2 => n2077,
                           ZN => n1389);
   U548 : OAI22_X1 port map( A1 => n2049, A2 => n2083, B1 => n841, B2 => n2077,
                           ZN => n1388);
   U549 : OAI22_X1 port map( A1 => n2050, A2 => n2083, B1 => n843, B2 => n2077,
                           ZN => n1387);
   U550 : OAI22_X1 port map( A1 => n2051, A2 => n2083, B1 => n845, B2 => n2077,
                           ZN => n1386);
   U551 : OAI22_X1 port map( A1 => n2052, A2 => n2083, B1 => n847, B2 => n2076,
                           ZN => n1385);
   U552 : OAI22_X1 port map( A1 => n2053, A2 => n2082, B1 => n849, B2 => n2076,
                           ZN => n1384);
   U553 : OAI22_X1 port map( A1 => n2054, A2 => n2082, B1 => n851, B2 => n2076,
                           ZN => n1383);
   U554 : OAI22_X1 port map( A1 => n2055, A2 => n2082, B1 => n853, B2 => n2076,
                           ZN => n1382);
   U555 : OAI22_X1 port map( A1 => n2056, A2 => n2082, B1 => n855, B2 => n2076,
                           ZN => n1381);
   U556 : OAI22_X1 port map( A1 => n2057, A2 => n2082, B1 => n857, B2 => n2076,
                           ZN => n1380);
   U557 : OAI22_X1 port map( A1 => n2058, A2 => n2082, B1 => n859, B2 => n2076,
                           ZN => n1379);
   U558 : OAI22_X1 port map( A1 => n2059, A2 => n2082, B1 => n861, B2 => n2076,
                           ZN => n1378);
   U559 : OAI22_X1 port map( A1 => n2060, A2 => n2082, B1 => n863, B2 => n2076,
                           ZN => n1377);
   U560 : OAI22_X1 port map( A1 => n2061, A2 => n2082, B1 => n865, B2 => n2076,
                           ZN => n1376);
   U561 : OAI22_X1 port map( A1 => n2062, A2 => n2082, B1 => n867, B2 => n2076,
                           ZN => n1375);
   U562 : OAI22_X1 port map( A1 => n2063, A2 => n2082, B1 => n871, B2 => n2076,
                           ZN => n1374);
   U563 : OAI22_X1 port map( A1 => n2014, A2 => n2075, B1 => n751, B2 => n2068,
                           ZN => n1369);
   U564 : OAI22_X1 port map( A1 => n2015, A2 => n2074, B1 => n753, B2 => n2068,
                           ZN => n1368);
   U565 : OAI22_X1 port map( A1 => n2016, A2 => n2074, B1 => n755, B2 => n2068,
                           ZN => n1367);
   U566 : OAI22_X1 port map( A1 => n2017, A2 => n2074, B1 => n757, B2 => n2068,
                           ZN => n1366);
   U567 : OAI22_X1 port map( A1 => n2018, A2 => n2074, B1 => n759, B2 => n2068,
                           ZN => n1365);
   U568 : OAI22_X1 port map( A1 => n2019, A2 => n2074, B1 => n761, B2 => n2068,
                           ZN => n1364);
   U569 : OAI22_X1 port map( A1 => n2020, A2 => n2074, B1 => n763, B2 => n2068,
                           ZN => n1363);
   U570 : OAI22_X1 port map( A1 => n2021, A2 => n2074, B1 => n765, B2 => n2068,
                           ZN => n1362);
   U571 : OAI22_X1 port map( A1 => n2022, A2 => n2074, B1 => n767, B2 => n2068,
                           ZN => n1361);
   U572 : OAI22_X1 port map( A1 => n2023, A2 => n2074, B1 => n769, B2 => n2068,
                           ZN => n1360);
   U573 : OAI22_X1 port map( A1 => n2024, A2 => n2074, B1 => n771, B2 => n2068,
                           ZN => n1359);
   U574 : OAI22_X1 port map( A1 => n2025, A2 => n2074, B1 => n773, B2 => n2068,
                           ZN => n1358);
   U575 : OAI22_X1 port map( A1 => n2026, A2 => n2074, B1 => n775, B2 => n2067,
                           ZN => n1357);
   U576 : OAI22_X1 port map( A1 => n2027, A2 => n2073, B1 => n777, B2 => n2067,
                           ZN => n1356);
   U577 : OAI22_X1 port map( A1 => n2028, A2 => n2073, B1 => n779, B2 => n2067,
                           ZN => n1355);
   U578 : OAI22_X1 port map( A1 => n1738, A2 => n2073, B1 => n781, B2 => n2067,
                           ZN => n1354);
   U579 : OAI22_X1 port map( A1 => n1737, A2 => n2073, B1 => n783, B2 => n2067,
                           ZN => n1353);
   U580 : OAI22_X1 port map( A1 => n1736, A2 => n2073, B1 => n785, B2 => n2067,
                           ZN => n1352);
   U581 : OAI22_X1 port map( A1 => n1735, A2 => n2073, B1 => n787, B2 => n2067,
                           ZN => n1351);
   U582 : OAI22_X1 port map( A1 => n1734, A2 => n2073, B1 => n789, B2 => n2067,
                           ZN => n1350);
   U583 : OAI22_X1 port map( A1 => n1733, A2 => n2073, B1 => n791, B2 => n2067,
                           ZN => n1349);
   U584 : OAI22_X1 port map( A1 => n1732, A2 => n2073, B1 => n793, B2 => n2067,
                           ZN => n1348);
   U585 : OAI22_X1 port map( A1 => n1731, A2 => n2073, B1 => n795, B2 => n2067,
                           ZN => n1347);
   U586 : OAI22_X1 port map( A1 => n1730, A2 => n2073, B1 => n797, B2 => n2067,
                           ZN => n1346);
   U587 : OAI22_X1 port map( A1 => n1729, A2 => n2073, B1 => n799, B2 => n2066,
                           ZN => n1345);
   U588 : OAI22_X1 port map( A1 => n1728, A2 => n2072, B1 => n801, B2 => n2066,
                           ZN => n1344);
   U589 : OAI22_X1 port map( A1 => n1727, A2 => n2072, B1 => n803, B2 => n2066,
                           ZN => n1343);
   U590 : OAI22_X1 port map( A1 => n1726, A2 => n2072, B1 => n805, B2 => n2066,
                           ZN => n1342);
   U591 : OAI22_X1 port map( A1 => n1725, A2 => n2072, B1 => n807, B2 => n2066,
                           ZN => n1341);
   U592 : OAI22_X1 port map( A1 => n1724, A2 => n2072, B1 => n809, B2 => n2066,
                           ZN => n1340);
   U593 : OAI22_X1 port map( A1 => n1723, A2 => n2072, B1 => n811, B2 => n2066,
                           ZN => n1339);
   U594 : OAI22_X1 port map( A1 => n1722, A2 => n2072, B1 => n813, B2 => n2066,
                           ZN => n1338);
   U595 : OAI22_X1 port map( A1 => n1721, A2 => n2072, B1 => n815, B2 => n2066,
                           ZN => n1337);
   U596 : OAI22_X1 port map( A1 => n1720, A2 => n2072, B1 => n817, B2 => n2066,
                           ZN => n1336);
   U597 : OAI22_X1 port map( A1 => n1719, A2 => n2072, B1 => n819, B2 => n2066,
                           ZN => n1335);
   U598 : OAI22_X1 port map( A1 => n1718, A2 => n2072, B1 => n821, B2 => n2066,
                           ZN => n1334);
   U599 : OAI22_X1 port map( A1 => n1717, A2 => n2072, B1 => n823, B2 => n2065,
                           ZN => n1333);
   U600 : OAI22_X1 port map( A1 => n1716, A2 => n2071, B1 => n825, B2 => n2065,
                           ZN => n1332);
   U601 : OAI22_X1 port map( A1 => n1715, A2 => n2071, B1 => n827, B2 => n2065,
                           ZN => n1331);
   U602 : OAI22_X1 port map( A1 => n1714, A2 => n2071, B1 => n829, B2 => n2065,
                           ZN => n1330);
   U603 : OAI22_X1 port map( A1 => n1713, A2 => n2071, B1 => n831, B2 => n2065,
                           ZN => n1329);
   U604 : OAI22_X1 port map( A1 => n1712, A2 => n2071, B1 => n833, B2 => n2065,
                           ZN => n1328);
   U605 : OAI22_X1 port map( A1 => n1711, A2 => n2071, B1 => n835, B2 => n2065,
                           ZN => n1327);
   U606 : OAI22_X1 port map( A1 => n1710, A2 => n2071, B1 => n837, B2 => n2065,
                           ZN => n1326);
   U607 : OAI22_X1 port map( A1 => n1709, A2 => n2071, B1 => n839, B2 => n2065,
                           ZN => n1325);
   U608 : OAI22_X1 port map( A1 => n1708, A2 => n2071, B1 => n841, B2 => n2065,
                           ZN => n1324);
   U609 : OAI22_X1 port map( A1 => n1707, A2 => n2071, B1 => n843, B2 => n2065,
                           ZN => n1323);
   U610 : OAI22_X1 port map( A1 => n1706, A2 => n2071, B1 => n845, B2 => n2065,
                           ZN => n1322);
   U611 : OAI22_X1 port map( A1 => n1705, A2 => n2071, B1 => n847, B2 => n2064,
                           ZN => n1321);
   U612 : OAI22_X1 port map( A1 => n1704, A2 => n2070, B1 => n849, B2 => n2064,
                           ZN => n1320);
   U613 : OAI22_X1 port map( A1 => n1703, A2 => n2070, B1 => n851, B2 => n2064,
                           ZN => n1319);
   U614 : OAI22_X1 port map( A1 => n1702, A2 => n2070, B1 => n853, B2 => n2064,
                           ZN => n1318);
   U615 : OAI22_X1 port map( A1 => n1701, A2 => n2070, B1 => n855, B2 => n2064,
                           ZN => n1317);
   U616 : OAI22_X1 port map( A1 => n1700, A2 => n2070, B1 => n857, B2 => n2064,
                           ZN => n1316);
   U617 : OAI22_X1 port map( A1 => n1699, A2 => n2070, B1 => n859, B2 => n2064,
                           ZN => n1315);
   U618 : OAI22_X1 port map( A1 => n1698, A2 => n2070, B1 => n861, B2 => n2064,
                           ZN => n1314);
   U619 : OAI22_X1 port map( A1 => n1697, A2 => n2070, B1 => n863, B2 => n2064,
                           ZN => n1313);
   U620 : OAI22_X1 port map( A1 => n1696, A2 => n2070, B1 => n865, B2 => n2064,
                           ZN => n1312);
   U621 : OAI22_X1 port map( A1 => n1695, A2 => n2070, B1 => n867, B2 => n2064,
                           ZN => n1311);
   U622 : OAI22_X1 port map( A1 => n1694, A2 => n2070, B1 => n871, B2 => n2064,
                           ZN => n1310);
   U623 : INV_X1 port map( A => DATAIN(0), ZN => n743);
   U624 : INV_X1 port map( A => DATAIN(1), ZN => n745);
   U625 : INV_X1 port map( A => DATAIN(2), ZN => n747);
   U626 : INV_X1 port map( A => DATAIN(3), ZN => n749);
   U627 : INV_X1 port map( A => DATAIN(4), ZN => n751);
   U628 : INV_X1 port map( A => DATAIN(5), ZN => n753);
   U629 : INV_X1 port map( A => DATAIN(6), ZN => n755);
   U630 : INV_X1 port map( A => DATAIN(7), ZN => n757);
   U631 : INV_X1 port map( A => DATAIN(8), ZN => n759);
   U632 : INV_X1 port map( A => DATAIN(9), ZN => n761);
   U633 : INV_X1 port map( A => DATAIN(10), ZN => n763);
   U634 : INV_X1 port map( A => DATAIN(11), ZN => n765);
   U635 : INV_X1 port map( A => DATAIN(12), ZN => n767);
   U636 : INV_X1 port map( A => DATAIN(13), ZN => n769);
   U637 : INV_X1 port map( A => DATAIN(14), ZN => n771);
   U638 : INV_X1 port map( A => DATAIN(15), ZN => n773);
   U639 : INV_X1 port map( A => DATAIN(16), ZN => n775);
   U640 : INV_X1 port map( A => DATAIN(17), ZN => n777);
   U641 : INV_X1 port map( A => DATAIN(18), ZN => n779);
   U642 : INV_X1 port map( A => DATAIN(19), ZN => n781);
   U643 : INV_X1 port map( A => DATAIN(20), ZN => n783);
   U644 : INV_X1 port map( A => DATAIN(21), ZN => n785);
   U645 : INV_X1 port map( A => DATAIN(22), ZN => n787);
   U646 : INV_X1 port map( A => DATAIN(23), ZN => n789);
   U647 : INV_X1 port map( A => DATAIN(24), ZN => n791);
   U648 : INV_X1 port map( A => DATAIN(25), ZN => n793);
   U649 : INV_X1 port map( A => DATAIN(26), ZN => n795);
   U650 : INV_X1 port map( A => DATAIN(27), ZN => n797);
   U651 : INV_X1 port map( A => DATAIN(28), ZN => n799);
   U652 : INV_X1 port map( A => DATAIN(29), ZN => n801);
   U653 : INV_X1 port map( A => DATAIN(30), ZN => n803);
   U654 : INV_X1 port map( A => DATAIN(31), ZN => n805);
   U655 : INV_X1 port map( A => DATAIN(32), ZN => n807);
   U656 : INV_X1 port map( A => DATAIN(33), ZN => n809);
   U657 : INV_X1 port map( A => DATAIN(34), ZN => n811);
   U658 : INV_X1 port map( A => DATAIN(35), ZN => n813);
   U659 : INV_X1 port map( A => DATAIN(36), ZN => n815);
   U660 : INV_X1 port map( A => DATAIN(37), ZN => n817);
   U661 : INV_X1 port map( A => DATAIN(38), ZN => n819);
   U662 : INV_X1 port map( A => DATAIN(39), ZN => n821);
   U663 : INV_X1 port map( A => DATAIN(40), ZN => n823);
   U664 : INV_X1 port map( A => DATAIN(41), ZN => n825);
   U665 : INV_X1 port map( A => DATAIN(42), ZN => n827);
   U666 : INV_X1 port map( A => DATAIN(43), ZN => n829);
   U667 : INV_X1 port map( A => DATAIN(44), ZN => n831);
   U668 : INV_X1 port map( A => DATAIN(45), ZN => n833);
   U669 : INV_X1 port map( A => DATAIN(46), ZN => n835);
   U670 : INV_X1 port map( A => DATAIN(47), ZN => n837);
   U671 : INV_X1 port map( A => DATAIN(48), ZN => n839);
   U672 : INV_X1 port map( A => DATAIN(49), ZN => n841);
   U673 : INV_X1 port map( A => DATAIN(50), ZN => n843);
   U674 : INV_X1 port map( A => DATAIN(51), ZN => n845);
   U675 : INV_X1 port map( A => DATAIN(52), ZN => n847);
   U676 : INV_X1 port map( A => DATAIN(53), ZN => n849);
   U677 : INV_X1 port map( A => DATAIN(54), ZN => n851);
   U678 : INV_X1 port map( A => DATAIN(55), ZN => n853);
   U679 : INV_X1 port map( A => DATAIN(56), ZN => n855);
   U680 : INV_X1 port map( A => DATAIN(57), ZN => n857);
   U681 : INV_X1 port map( A => DATAIN(58), ZN => n859);
   U682 : INV_X1 port map( A => DATAIN(59), ZN => n861);
   U683 : INV_X1 port map( A => DATAIN(60), ZN => n863);
   U684 : INV_X1 port map( A => DATAIN(61), ZN => n865);
   U685 : INV_X1 port map( A => DATAIN(62), ZN => n867);
   U686 : INV_X1 port map( A => DATAIN(63), ZN => n871);
   U687 : CLKBUF_X1 port map( A => n979, Z => n2069);
   U688 : CLKBUF_X1 port map( A => n978, Z => n2075);
   U689 : CLKBUF_X1 port map( A => n939, Z => n2081);
   U690 : CLKBUF_X1 port map( A => n938, Z => n2087);
   U691 : CLKBUF_X1 port map( A => n876, Z => n2093);
   U692 : CLKBUF_X1 port map( A => n875, Z => n2099);
   U693 : CLKBUF_X1 port map( A => n742, Z => n2105);
   U694 : CLKBUF_X1 port map( A => n741, Z => n2111);
   U695 : CLKBUF_X1 port map( A => n740, Z => n2117);
   U696 : CLKBUF_X1 port map( A => n739, Z => n2123);
   U697 : CLKBUF_X1 port map( A => n738, Z => n2129);
   U698 : CLKBUF_X1 port map( A => n736, Z => n2135);
   U699 : CLKBUF_X1 port map( A => n735, Z => n2141);
   U700 : CLKBUF_X1 port map( A => n527, Z => n2147);
   U701 : CLKBUF_X1 port map( A => n525, Z => n2158);
   U702 : CLKBUF_X1 port map( A => n523, Z => n2164);
   U703 : CLKBUF_X1 port map( A => n521, Z => n2170);
   U704 : INV_X1 port map( A => ADD_RD2(0), ZN => n2171);
   U705 : INV_X1 port map( A => ADD_RD2(1), ZN => n2172);
   U706 : INV_X1 port map( A => ADD_RD1(0), ZN => n2173);
   U707 : INV_X1 port map( A => ADD_RD1(1), ZN => n2174);
   U708 : INV_X1 port map( A => ADD_WR(0), ZN => n2175);
   U709 : INV_X1 port map( A => ADD_WR(1), ZN => n2176);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4.all;

entity register_file_reg_size64_file_size4_4 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_reg_size64_file_size4_4;

architecture SYN_BEHAVIORAL of register_file_reg_size64_file_size4_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n415, n1200, n1202, n1204, n1310, n1311, n1312, n1313, n1314, n1315
      , n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n871, n872, 
      n873, n875, n876, n936, n938, n939, n975, n978, n979, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176 : std_logic
      ;

begin
   
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => n174,
                           QN => n2028);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => n175,
                           QN => n2027);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => n176,
                           QN => n2026);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => n177,
                           QN => n2025);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => n178,
                           QN => n2024);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => n179,
                           QN => n2023);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => n180,
                           QN => n2022);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => n181,
                           QN => n2021);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => n182,
                           QN => n2020);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => n183, 
                           QN => n2019);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => n184, 
                           QN => n2018);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => n185, 
                           QN => n2017);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => n186, 
                           QN => n2016);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => n187, 
                           QN => n2015);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => n188, 
                           QN => n2014);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => n189, 
                           QN => n2013);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => n190, 
                           QN => n2012);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => n191, 
                           QN => n2011);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => n192, 
                           QN => n2010);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => n65, 
                           QN => n2063);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => n66, 
                           QN => n2062);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n67, 
                           QN => n2061);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => n68, 
                           QN => n2060);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => n69, 
                           QN => n2059);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => n70, 
                           QN => n2058);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => n71, 
                           QN => n2057);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => n72, 
                           QN => n2056);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => n73, 
                           QN => n2055);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => n74, 
                           QN => n2054);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => n75, 
                           QN => n2053);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => n76, 
                           QN => n2052);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => n77, 
                           QN => n2051);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => n78, 
                           QN => n2050);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => n79, 
                           QN => n2049);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => n80, 
                           QN => n2048);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => n81, 
                           QN => n2047);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => n82, 
                           QN => n2046);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => n83, 
                           QN => n2045);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => n84, 
                           QN => n2044);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => n85, 
                           QN => n2043);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => n86, 
                           QN => n2042);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => n87, 
                           QN => n2041);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => n88, 
                           QN => n2040);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => n89, 
                           QN => n2039);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => n90, 
                           QN => n2038);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => n91, 
                           QN => n2037);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => n92, 
                           QN => n2036);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => n93, 
                           QN => n2035);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => n94, 
                           QN => n2034);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => n95, 
                           QN => n2033);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => n96, 
                           QN => n2032);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => n97, 
                           QN => n2031);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => n98, 
                           QN => n2030);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => n99, 
                           QN => n2029);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => n2, 
                           QN => n2009);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => n3, 
                           QN => n2008);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => n4, 
                           QN => n2007);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => n5, 
                           QN => n2006);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => n6, 
                           QN => n2005);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => n7, 
                           QN => n2004);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => n8, 
                           QN => n2003);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => n9, 
                           QN => n2002);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => n13, 
                           QN => n2001);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => n14, 
                           QN => n2000);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => n15, 
                           QN => n1999);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => n16, 
                           QN => n1998);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => n17, 
                           QN => n1997);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => n18, 
                           QN => n1996);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => n19, 
                           QN => n1995);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => n20, 
                           QN => n1994);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => n21, 
                           QN => n1993);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => n22, 
                           QN => n1992);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => n23, 
                           QN => n1991);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => n24, 
                           QN => n1990);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => n25, 
                           QN => n1989);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => n26, 
                           QN => n1988);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n27, 
                           QN => n1987);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => n28, 
                           QN => n1986);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n29, 
                           QN => n1985);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => n30, 
                           QN => n1984);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n31, 
                           QN => n1983);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => n32, 
                           QN => n1982);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n33, 
                           QN => n1981);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => n34, 
                           QN => n1980);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n35, 
                           QN => n1979);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => n36, 
                           QN => n1978);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => n37, 
                           QN => n1977);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => n38, 
                           QN => n1976);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => n39, 
                           QN => n1975);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => n40, 
                           QN => n1974);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => n41, 
                           QN => n1973);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => n42, 
                           QN => n1972);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => n43, 
                           QN => n1971);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => n44, 
                           QN => n1970);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => n45, 
                           QN => n1969);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => n46, 
                           QN => n1968);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => n47, 
                           QN => n1967);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => n48, 
                           QN => n1966);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => n49, 
                           QN => n1965);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => n50, 
                           QN => n1964);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => n51, 
                           QN => n1963);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => n52, 
                           QN => n1962);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => n53, 
                           QN => n1961);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => n54, 
                           QN => n1960);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n55, 
                           QN => n1959);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => n56, 
                           QN => n1958);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n57, 
                           QN => n1957);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => n58, 
                           QN => n1956);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n59, 
                           QN => n1955);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => n60, 
                           QN => n1954);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n61, 
                           QN => n1953);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => n62, 
                           QN => n1952);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n63, 
                           QN => n1951);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => n64, 
                           QN => n1950);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n999,
                           QN => n728);
   OUT2_reg_63_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => OUT2(63), QN
                           => n1822);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n1000
                           , QN => n725);
   OUT2_reg_62_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => OUT2(62), QN
                           => n1823);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n1001
                           , QN => n722);
   OUT2_reg_61_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => OUT2(61), QN
                           => n1824);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n1002
                           , QN => n719);
   OUT2_reg_60_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => OUT2(60), QN
                           => n1825);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n1003
                           , QN => n716);
   OUT2_reg_59_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => OUT2(59), QN
                           => n1826);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n1004
                           , QN => n713);
   OUT2_reg_58_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => OUT2(58), QN
                           => n1827);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n1005
                           , QN => n710);
   OUT2_reg_57_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => OUT2(57), QN
                           => n1828);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n1006
                           , QN => n707);
   OUT2_reg_56_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => OUT2(56), QN
                           => n1829);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n1007
                           , QN => n704);
   OUT2_reg_55_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => OUT2(55), QN
                           => n1830);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n1008
                           , QN => n700);
   OUT2_reg_54_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => OUT2(54), QN
                           => n1831);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n1009
                           , QN => n696);
   OUT2_reg_53_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => OUT2(53), QN
                           => n1832);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n1010
                           , QN => n692);
   OUT2_reg_52_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => OUT2(52), QN
                           => n1833);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n1011
                           , QN => n689);
   OUT2_reg_51_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => OUT2(51), QN
                           => n1834);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n1012
                           , QN => n686);
   OUT2_reg_50_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => OUT2(50), QN
                           => n1835);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n1013
                           , QN => n683);
   OUT2_reg_49_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => OUT2(49), QN
                           => n1836);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n1014
                           , QN => n680);
   OUT2_reg_48_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => OUT2(48), QN
                           => n1837);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n1015
                           , QN => n677);
   OUT2_reg_47_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => OUT2(47), QN
                           => n1838);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n1016
                           , QN => n674);
   OUT2_reg_46_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => OUT2(46), QN
                           => n1839);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n1017
                           , QN => n671);
   OUT2_reg_45_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => OUT2(45), QN
                           => n1840);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n1018
                           , QN => n668);
   OUT2_reg_44_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => OUT2(44), QN
                           => n1841);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n1019
                           , QN => n665);
   OUT2_reg_43_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => OUT2(43), QN
                           => n1842);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n1020
                           , QN => n662);
   OUT2_reg_42_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => OUT2(42), QN
                           => n1843);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n1021
                           , QN => n659);
   OUT2_reg_41_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => OUT2(41), QN
                           => n1844);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n1022
                           , QN => n656);
   OUT2_reg_40_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => OUT2(40), QN
                           => n1845);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n1023
                           , QN => n653);
   OUT2_reg_39_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => OUT2(39), QN
                           => n1846);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n1024
                           , QN => n650);
   OUT2_reg_38_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => OUT2(38), QN
                           => n1847);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n1025
                           , QN => n647);
   OUT2_reg_37_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => OUT2(37), QN
                           => n1848);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n1026
                           , QN => n644);
   OUT2_reg_36_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => OUT2(36), QN
                           => n1849);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n1027
                           , QN => n641);
   OUT2_reg_35_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => OUT2(35), QN
                           => n1850);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n1028
                           , QN => n638);
   OUT2_reg_34_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => OUT2(34), QN
                           => n1851);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n1029
                           , QN => n635);
   OUT2_reg_33_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => OUT2(33), QN
                           => n1852);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n1030
                           , QN => n632);
   OUT2_reg_32_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => OUT2(32), QN
                           => n1853);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n1031
                           , QN => n629);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => OUT2(31), QN
                           => n1854);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n1032
                           , QN => n626);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => OUT2(30), QN
                           => n1855);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n1033
                           , QN => n623);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => OUT2(29), QN
                           => n1856);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n1034
                           , QN => n619);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => OUT2(28), QN
                           => n1857);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n1035
                           , QN => n615);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => OUT2(27), QN
                           => n1858);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n1036
                           , QN => n611);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => OUT2(26), QN
                           => n1859);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n1037
                           , QN => n607);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => OUT2(25), QN
                           => n1860);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n1038
                           , QN => n603);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => OUT2(24), QN
                           => n1861);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n1039
                           , QN => n599);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => OUT2(23), QN
                           => n1862);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n1040
                           , QN => n595);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => OUT2(22), QN
                           => n1863);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n1041
                           , QN => n591);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => OUT2(21), QN
                           => n1864);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n1042
                           , QN => n587);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => OUT2(20), QN
                           => n1865);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n1043
                           , QN => n583);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => OUT2(19), QN
                           => n1866);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n1044
                           , QN => n580);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => OUT2(18), QN
                           => n1867);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n1045
                           , QN => n577);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => OUT2(17), QN
                           => n1868);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n1046
                           , QN => n574);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => OUT2(16), QN
                           => n1869);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n1047
                           , QN => n571);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => OUT2(15), QN
                           => n1870);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n1048
                           , QN => n568);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => OUT2(14), QN
                           => n1871);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n1049
                           , QN => n565);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => OUT2(13), QN
                           => n1872);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n1050
                           , QN => n562);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => OUT2(12), QN
                           => n1873);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n1051
                           , QN => n559);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => OUT2(11), QN
                           => n1874);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n1052
                           , QN => n556);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => OUT2(10), QN
                           => n1875);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n1053,
                           QN => n553);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => OUT2(9), QN 
                           => n1876);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => n1054,
                           QN => n550);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => OUT2(8), QN 
                           => n1877);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => n1055,
                           QN => n547);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => OUT2(7), QN 
                           => n1878);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => n1056,
                           QN => n544);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => OUT2(6), QN 
                           => n1879);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => n1057,
                           QN => n541);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => OUT2(5), QN 
                           => n1880);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => n1058,
                           QN => n538);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => OUT2(4), QN 
                           => n1881);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => n1059,
                           QN => n535);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => OUT2(3), QN 
                           => n1882);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n1060,
                           QN => n532);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => OUT2(2), QN 
                           => n1883);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n1061,
                           QN => n529);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => OUT2(1), QN 
                           => n1884);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n1062,
                           QN => n522);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => OUT2(0), QN 
                           => n1885);
   OUT1_reg_63_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => OUT1(63), QN
                           => n1886);
   OUT1_reg_62_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => OUT1(62), QN
                           => n1887);
   OUT1_reg_61_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => OUT1(61), QN
                           => n1888);
   OUT1_reg_60_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => OUT1(60), QN
                           => n1889);
   OUT1_reg_59_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => OUT1(59), QN
                           => n1890);
   OUT1_reg_58_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => OUT1(58), QN
                           => n1891);
   OUT1_reg_57_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => OUT1(57), QN
                           => n1892);
   OUT1_reg_56_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => OUT1(56), QN
                           => n1893);
   OUT1_reg_55_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => OUT1(55), QN
                           => n1894);
   OUT1_reg_54_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => OUT1(54), QN
                           => n1895);
   OUT1_reg_53_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => OUT1(53), QN
                           => n1896);
   OUT1_reg_52_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => OUT1(52), QN
                           => n1897);
   OUT1_reg_51_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => OUT1(51), QN
                           => n1898);
   OUT1_reg_50_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => OUT1(50), QN
                           => n1899);
   OUT1_reg_49_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => OUT1(49), QN
                           => n1900);
   OUT1_reg_48_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => OUT1(48), QN
                           => n1901);
   OUT1_reg_47_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => OUT1(47), QN
                           => n1902);
   OUT1_reg_46_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => OUT1(46), QN
                           => n1903);
   OUT1_reg_45_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => OUT1(45), QN
                           => n1904);
   OUT1_reg_44_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => OUT1(44), QN
                           => n1905);
   OUT1_reg_43_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => OUT1(43), QN
                           => n1906);
   OUT1_reg_42_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => OUT1(42), QN
                           => n1907);
   OUT1_reg_41_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => OUT1(41), QN
                           => n1908);
   OUT1_reg_40_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => OUT1(40), QN
                           => n1909);
   OUT1_reg_39_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => OUT1(39), QN
                           => n1910);
   OUT1_reg_38_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => OUT1(38), QN
                           => n1911);
   OUT1_reg_37_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => OUT1(37), QN
                           => n1912);
   OUT1_reg_36_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => OUT1(36), QN
                           => n1913);
   OUT1_reg_35_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => OUT1(35), QN
                           => n1914);
   OUT1_reg_34_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => OUT1(34), QN
                           => n1915);
   OUT1_reg_33_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => OUT1(33), QN
                           => n1916);
   OUT1_reg_32_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => OUT1(32), QN
                           => n1917);
   OUT1_reg_31_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => OUT1(31), QN
                           => n1918);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => OUT1(30), QN
                           => n1919);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => OUT1(29), QN
                           => n1920);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => OUT1(28), QN
                           => n1921);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => OUT1(27), QN
                           => n1922);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => OUT1(26), QN
                           => n1923);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => OUT1(25), QN
                           => n1924);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => OUT1(24), QN
                           => n1925);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => OUT1(23), QN
                           => n1926);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => OUT1(22), QN
                           => n1927);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => OUT1(21), QN
                           => n1928);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => OUT1(20), QN
                           => n1929);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => OUT1(19), QN
                           => n1930);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => OUT1(18), QN
                           => n1931);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => OUT1(17), QN
                           => n1932);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => OUT1(16), QN
                           => n1933);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => OUT1(15), QN
                           => n1934);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => OUT1(14), QN
                           => n1935);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => OUT1(13), QN
                           => n1936);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => OUT1(12), QN
                           => n1937);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => OUT1(11), QN
                           => n1938);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => OUT1(10), QN
                           => n1939);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => OUT1(9), QN 
                           => n1940);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => OUT1(8), QN 
                           => n1941);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => OUT1(7), QN 
                           => n1942);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => OUT1(6), QN 
                           => n1943);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => OUT1(5), QN 
                           => n1944);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => OUT1(4), QN 
                           => n1945);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => OUT1(3), QN 
                           => n1946);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => OUT1(2), QN 
                           => n1947);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => OUT1(1), QN 
                           => n1948);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => OUT1(0), QN 
                           => n1949);
   U859 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n2164, A3 => ADD_RD1(1), 
                           ZN => n521);
   U860 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n2135, A3 => ADD_RD2(1), 
                           ZN => n735);
   U861 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n873, A3 => ADD_WR(1), ZN 
                           => n872);
   U862 : NAND3_X1 port map( A1 => n873, A2 => n2175, A3 => ADD_WR(1), ZN => 
                           n936);
   U863 : NAND3_X1 port map( A1 => n873, A2 => n2176, A3 => ADD_WR(0), ZN => 
                           n975);
   U864 : NAND3_X1 port map( A1 => n2175, A2 => n2176, A3 => n873, ZN => n998);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => n537, 
                           QN => n1818);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => n534, 
                           QN => n1819);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => n531, 
                           QN => n1820);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => n528, 
                           QN => n1821);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => n730,
                           QN => n415);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => n702,
                           QN => n1200);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => n698,
                           QN => n1202);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => n694,
                           QN => n1204);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => n622,
                           QN => n1793);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => n618,
                           QN => n1794);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => n614,
                           QN => n1795);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => n610,
                           QN => n1796);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => n606,
                           QN => n1797);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => n602,
                           QN => n1798);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => n598,
                           QN => n1799);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => n594,
                           QN => n1800);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => n590,
                           QN => n1801);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => n586,
                           QN => n1802);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => n582,
                           QN => n1803);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => n579,
                           QN => n1804);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => n576,
                           QN => n1805);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => n573,
                           QN => n1806);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => n570,
                           QN => n1807);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => n567,
                           QN => n1808);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => n564,
                           QN => n1809);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => n561,
                           QN => n1810);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => n558,
                           QN => n1811);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => n555, 
                           QN => n1812);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => n552, 
                           QN => n1813);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => n549, 
                           QN => n1814);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => n546, 
                           QN => n1815);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => n543, 
                           QN => n1816);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => n540, 
                           QN => n1817);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => n731,
                           QN => n1694);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => n727,
                           QN => n1695);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => n724,
                           QN => n1696);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => n721,
                           QN => n1697);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => n718,
                           QN => n1698);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => n715,
                           QN => n1699);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => n712,
                           QN => n1700);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => n709,
                           QN => n1701);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => n706,
                           QN => n1702);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => n703,
                           QN => n1703);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => n699,
                           QN => n1704);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => n695,
                           QN => n1705);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => n691,
                           QN => n1706);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => n688,
                           QN => n1707);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => n685,
                           QN => n1708);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => n682,
                           QN => n1709);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => n679,
                           QN => n1710);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => n676,
                           QN => n1711);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => n673,
                           QN => n1712);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => n670,
                           QN => n1713);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => n667,
                           QN => n1714);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => n664,
                           QN => n1715);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => n661,
                           QN => n1716);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => n658,
                           QN => n1717);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => n655,
                           QN => n1718);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => n652,
                           QN => n1719);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => n649,
                           QN => n1720);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => n646,
                           QN => n1721);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => n643,
                           QN => n1722);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => n640,
                           QN => n1723);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => n637,
                           QN => n1724);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => n634,
                           QN => n1725);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => n631,
                           QN => n1726);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => n628,
                           QN => n1727);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n625,
                           QN => n1728);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => n621,
                           QN => n1729);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => n617,
                           QN => n1730);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => n613,
                           QN => n1731);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => n609,
                           QN => n1732);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => n605,
                           QN => n1733);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => n601,
                           QN => n1734);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => n597,
                           QN => n1735);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => n593,
                           QN => n1736);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => n589,
                           QN => n1737);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => n585,
                           QN => n1738);
   U3 : BUF_X1 port map( A => n521, Z => n2167);
   U4 : BUF_X1 port map( A => n521, Z => n2166);
   U5 : BUF_X1 port map( A => n521, Z => n2165);
   U6 : BUF_X1 port map( A => n735, Z => n2139);
   U7 : BUF_X1 port map( A => n735, Z => n2138);
   U8 : BUF_X1 port map( A => n735, Z => n2137);
   U9 : BUF_X1 port map( A => n735, Z => n2136);
   U10 : BUF_X1 port map( A => n521, Z => n2169);
   U11 : BUF_X1 port map( A => n521, Z => n2168);
   U12 : BUF_X1 port map( A => n735, Z => n2140);
   U13 : BUF_X1 port map( A => n526, Z => n2151);
   U14 : BUF_X1 port map( A => n526, Z => n2152);
   U15 : BUF_X1 port map( A => n527, Z => n2144);
   U16 : BUF_X1 port map( A => n527, Z => n2146);
   U17 : BUF_X1 port map( A => n527, Z => n2145);
   U18 : BUF_X1 port map( A => n523, Z => n2159);
   U19 : BUF_X1 port map( A => n523, Z => n2160);
   U20 : BUF_X1 port map( A => n523, Z => n2161);
   U21 : BUF_X1 port map( A => n523, Z => n2162);
   U22 : BUF_X1 port map( A => n523, Z => n2163);
   U23 : BUF_X1 port map( A => n736, Z => n2130);
   U24 : BUF_X1 port map( A => n736, Z => n2131);
   U25 : BUF_X1 port map( A => n736, Z => n2132);
   U26 : BUF_X1 port map( A => n736, Z => n2133);
   U27 : BUF_X1 port map( A => n736, Z => n2134);
   U28 : BUF_X1 port map( A => n525, Z => n2154);
   U29 : BUF_X1 port map( A => n525, Z => n2155);
   U30 : BUF_X1 port map( A => n525, Z => n2156);
   U31 : BUF_X1 port map( A => n525, Z => n2157);
   U32 : BUF_X1 port map( A => n738, Z => n2128);
   U33 : BUF_X1 port map( A => n738, Z => n2127);
   U34 : BUF_X1 port map( A => n738, Z => n2126);
   U35 : BUF_X1 port map( A => n738, Z => n2125);
   U36 : BUF_X1 port map( A => n738, Z => n2124);
   U37 : BUF_X1 port map( A => n742, Z => n2104);
   U38 : BUF_X1 port map( A => n742, Z => n2103);
   U39 : BUF_X1 port map( A => n742, Z => n2102);
   U40 : BUF_X1 port map( A => n742, Z => n2101);
   U41 : BUF_X1 port map( A => n739, Z => n2122);
   U42 : BUF_X1 port map( A => n739, Z => n2121);
   U43 : BUF_X1 port map( A => n739, Z => n2120);
   U44 : BUF_X1 port map( A => n739, Z => n2119);
   U45 : BUF_X1 port map( A => n739, Z => n2118);
   U46 : BUF_X1 port map( A => n740, Z => n2116);
   U47 : BUF_X1 port map( A => n740, Z => n2115);
   U48 : BUF_X1 port map( A => n740, Z => n2114);
   U49 : BUF_X1 port map( A => n740, Z => n2113);
   U50 : BUF_X1 port map( A => n740, Z => n2112);
   U51 : BUF_X1 port map( A => n741, Z => n2106);
   U52 : BUF_X1 port map( A => n875, Z => n2094);
   U53 : BUF_X1 port map( A => n938, Z => n2082);
   U54 : BUF_X1 port map( A => n978, Z => n2070);
   U55 : BUF_X1 port map( A => n741, Z => n2110);
   U56 : BUF_X1 port map( A => n741, Z => n2109);
   U57 : BUF_X1 port map( A => n741, Z => n2108);
   U58 : BUF_X1 port map( A => n741, Z => n2107);
   U59 : BUF_X1 port map( A => n875, Z => n2098);
   U60 : BUF_X1 port map( A => n875, Z => n2097);
   U61 : BUF_X1 port map( A => n875, Z => n2096);
   U62 : BUF_X1 port map( A => n875, Z => n2095);
   U63 : BUF_X1 port map( A => n938, Z => n2086);
   U64 : BUF_X1 port map( A => n938, Z => n2085);
   U65 : BUF_X1 port map( A => n938, Z => n2084);
   U66 : BUF_X1 port map( A => n938, Z => n2083);
   U67 : BUF_X1 port map( A => n978, Z => n2074);
   U68 : BUF_X1 port map( A => n978, Z => n2073);
   U69 : BUF_X1 port map( A => n978, Z => n2072);
   U70 : BUF_X1 port map( A => n978, Z => n2071);
   U71 : BUF_X1 port map( A => n526, Z => n2148);
   U72 : BUF_X1 port map( A => n526, Z => n2150);
   U73 : BUF_X1 port map( A => n876, Z => n2092);
   U74 : BUF_X1 port map( A => n876, Z => n2091);
   U75 : BUF_X1 port map( A => n876, Z => n2090);
   U76 : BUF_X1 port map( A => n876, Z => n2089);
   U77 : BUF_X1 port map( A => n876, Z => n2088);
   U78 : BUF_X1 port map( A => n939, Z => n2080);
   U79 : BUF_X1 port map( A => n939, Z => n2079);
   U80 : BUF_X1 port map( A => n939, Z => n2078);
   U81 : BUF_X1 port map( A => n939, Z => n2077);
   U82 : BUF_X1 port map( A => n939, Z => n2076);
   U83 : BUF_X1 port map( A => n979, Z => n2068);
   U84 : BUF_X1 port map( A => n979, Z => n2067);
   U85 : BUF_X1 port map( A => n979, Z => n2066);
   U86 : BUF_X1 port map( A => n979, Z => n2065);
   U87 : BUF_X1 port map( A => n979, Z => n2064);
   U88 : BUF_X1 port map( A => n527, Z => n2143);
   U89 : BUF_X1 port map( A => n527, Z => n2142);
   U90 : BUF_X1 port map( A => n526, Z => n2149);
   U91 : BUF_X1 port map( A => n525, Z => n2153);
   U92 : BUF_X1 port map( A => n742, Z => n2100);
   U93 : NAND2_X1 port map( A1 => n734, A2 => n872, ZN => n741);
   U94 : NAND2_X1 port map( A1 => n734, A2 => n936, ZN => n875);
   U95 : NAND2_X1 port map( A1 => n734, A2 => n2094, ZN => n876);
   U96 : NAND2_X1 port map( A1 => n734, A2 => n975, ZN => n938);
   U97 : NAND2_X1 port map( A1 => n734, A2 => n2082, ZN => n939);
   U98 : NAND2_X1 port map( A1 => n734, A2 => n998, ZN => n978);
   U99 : NAND2_X1 port map( A1 => n734, A2 => n2070, ZN => n979);
   U100 : OAI22_X1 port map( A1 => n538, A2 => n2111, B1 => n2104, B2 => n751, 
                           ZN => n1620);
   U101 : OAI22_X1 port map( A1 => n541, A2 => n2110, B1 => n2104, B2 => n753, 
                           ZN => n1618);
   U102 : OAI22_X1 port map( A1 => n544, A2 => n2110, B1 => n2104, B2 => n755, 
                           ZN => n1616);
   U103 : OAI22_X1 port map( A1 => n547, A2 => n2110, B1 => n2104, B2 => n757, 
                           ZN => n1614);
   U104 : OAI22_X1 port map( A1 => n550, A2 => n2110, B1 => n2104, B2 => n759, 
                           ZN => n1612);
   U105 : OAI22_X1 port map( A1 => n553, A2 => n2110, B1 => n2104, B2 => n761, 
                           ZN => n1610);
   U106 : OAI22_X1 port map( A1 => n556, A2 => n2110, B1 => n2104, B2 => n763, 
                           ZN => n1608);
   U107 : OAI22_X1 port map( A1 => n559, A2 => n2110, B1 => n2104, B2 => n765, 
                           ZN => n1606);
   U108 : OAI22_X1 port map( A1 => n562, A2 => n2110, B1 => n2104, B2 => n767, 
                           ZN => n1604);
   U109 : OAI22_X1 port map( A1 => n565, A2 => n2110, B1 => n2104, B2 => n769, 
                           ZN => n1602);
   U110 : OAI22_X1 port map( A1 => n568, A2 => n2110, B1 => n2104, B2 => n771, 
                           ZN => n1600);
   U111 : OAI22_X1 port map( A1 => n571, A2 => n2110, B1 => n2104, B2 => n773, 
                           ZN => n1598);
   U112 : OAI22_X1 port map( A1 => n574, A2 => n2110, B1 => n2103, B2 => n775, 
                           ZN => n1596);
   U113 : OAI22_X1 port map( A1 => n577, A2 => n2109, B1 => n2103, B2 => n777, 
                           ZN => n1594);
   U114 : OAI22_X1 port map( A1 => n580, A2 => n2109, B1 => n2103, B2 => n779, 
                           ZN => n1592);
   U115 : OAI22_X1 port map( A1 => n583, A2 => n2109, B1 => n2103, B2 => n781, 
                           ZN => n1590);
   U116 : OAI22_X1 port map( A1 => n587, A2 => n2109, B1 => n2103, B2 => n783, 
                           ZN => n1588);
   U117 : OAI22_X1 port map( A1 => n591, A2 => n2109, B1 => n2103, B2 => n785, 
                           ZN => n1586);
   U118 : OAI22_X1 port map( A1 => n595, A2 => n2109, B1 => n2103, B2 => n787, 
                           ZN => n1584);
   U119 : OAI22_X1 port map( A1 => n599, A2 => n2109, B1 => n2103, B2 => n789, 
                           ZN => n1582);
   U120 : OAI22_X1 port map( A1 => n603, A2 => n2109, B1 => n2103, B2 => n791, 
                           ZN => n1580);
   U121 : OAI22_X1 port map( A1 => n607, A2 => n2109, B1 => n2103, B2 => n793, 
                           ZN => n1578);
   U122 : OAI22_X1 port map( A1 => n611, A2 => n2109, B1 => n2103, B2 => n795, 
                           ZN => n1576);
   U123 : OAI22_X1 port map( A1 => n615, A2 => n2109, B1 => n2103, B2 => n797, 
                           ZN => n1574);
   U124 : OAI22_X1 port map( A1 => n619, A2 => n2109, B1 => n2102, B2 => n799, 
                           ZN => n1572);
   U125 : OAI22_X1 port map( A1 => n623, A2 => n2108, B1 => n2102, B2 => n801, 
                           ZN => n1570);
   U126 : OAI22_X1 port map( A1 => n626, A2 => n2108, B1 => n2102, B2 => n803, 
                           ZN => n1568);
   U127 : OAI22_X1 port map( A1 => n629, A2 => n2108, B1 => n2102, B2 => n805, 
                           ZN => n1566);
   U128 : OAI22_X1 port map( A1 => n632, A2 => n2108, B1 => n2102, B2 => n807, 
                           ZN => n1564);
   U129 : OAI22_X1 port map( A1 => n635, A2 => n2108, B1 => n2102, B2 => n809, 
                           ZN => n1562);
   U130 : OAI22_X1 port map( A1 => n638, A2 => n2108, B1 => n2102, B2 => n811, 
                           ZN => n1560);
   U131 : OAI22_X1 port map( A1 => n641, A2 => n2108, B1 => n2102, B2 => n813, 
                           ZN => n1558);
   U132 : OAI22_X1 port map( A1 => n644, A2 => n2108, B1 => n2102, B2 => n815, 
                           ZN => n1556);
   U133 : OAI22_X1 port map( A1 => n647, A2 => n2108, B1 => n2102, B2 => n817, 
                           ZN => n1554);
   U134 : OAI22_X1 port map( A1 => n650, A2 => n2108, B1 => n2102, B2 => n819, 
                           ZN => n1552);
   U135 : OAI22_X1 port map( A1 => n653, A2 => n2108, B1 => n2102, B2 => n821, 
                           ZN => n1550);
   U136 : OAI22_X1 port map( A1 => n656, A2 => n2108, B1 => n2101, B2 => n823, 
                           ZN => n1548);
   U137 : OAI22_X1 port map( A1 => n659, A2 => n2107, B1 => n2101, B2 => n825, 
                           ZN => n1546);
   U138 : OAI22_X1 port map( A1 => n662, A2 => n2107, B1 => n2101, B2 => n827, 
                           ZN => n1544);
   U139 : OAI22_X1 port map( A1 => n665, A2 => n2107, B1 => n2101, B2 => n829, 
                           ZN => n1542);
   U140 : OAI22_X1 port map( A1 => n668, A2 => n2107, B1 => n2101, B2 => n831, 
                           ZN => n1540);
   U141 : OAI22_X1 port map( A1 => n671, A2 => n2107, B1 => n2101, B2 => n833, 
                           ZN => n1538);
   U142 : OAI22_X1 port map( A1 => n674, A2 => n2107, B1 => n2101, B2 => n835, 
                           ZN => n1536);
   U143 : OAI22_X1 port map( A1 => n677, A2 => n2107, B1 => n2101, B2 => n837, 
                           ZN => n1534);
   U144 : OAI22_X1 port map( A1 => n680, A2 => n2107, B1 => n2101, B2 => n839, 
                           ZN => n1532);
   U145 : OAI22_X1 port map( A1 => n683, A2 => n2107, B1 => n2101, B2 => n841, 
                           ZN => n1530);
   U146 : OAI22_X1 port map( A1 => n686, A2 => n2107, B1 => n2101, B2 => n843, 
                           ZN => n1528);
   U147 : OAI22_X1 port map( A1 => n689, A2 => n2107, B1 => n2101, B2 => n845, 
                           ZN => n1526);
   U148 : OAI22_X1 port map( A1 => n522, A2 => n2111, B1 => n2105, B2 => n743, 
                           ZN => n1628);
   U149 : OAI22_X1 port map( A1 => n529, A2 => n2111, B1 => n2105, B2 => n745, 
                           ZN => n1626);
   U150 : OAI22_X1 port map( A1 => n532, A2 => n2111, B1 => n2105, B2 => n747, 
                           ZN => n1624);
   U151 : OAI22_X1 port map( A1 => n535, A2 => n2111, B1 => n2105, B2 => n749, 
                           ZN => n1622);
   U152 : OAI22_X1 port map( A1 => n692, A2 => n2107, B1 => n2100, B2 => n847, 
                           ZN => n1524);
   U153 : OAI22_X1 port map( A1 => n696, A2 => n2106, B1 => n2100, B2 => n849, 
                           ZN => n1522);
   U154 : OAI22_X1 port map( A1 => n700, A2 => n2106, B1 => n2100, B2 => n851, 
                           ZN => n1520);
   U155 : OAI22_X1 port map( A1 => n704, A2 => n2106, B1 => n2100, B2 => n853, 
                           ZN => n1518);
   U156 : OAI22_X1 port map( A1 => n707, A2 => n2106, B1 => n2100, B2 => n855, 
                           ZN => n1516);
   U157 : OAI22_X1 port map( A1 => n710, A2 => n2106, B1 => n2100, B2 => n857, 
                           ZN => n1514);
   U158 : OAI22_X1 port map( A1 => n713, A2 => n2106, B1 => n2100, B2 => n859, 
                           ZN => n1512);
   U159 : OAI22_X1 port map( A1 => n716, A2 => n2106, B1 => n2100, B2 => n861, 
                           ZN => n1510);
   U160 : OAI22_X1 port map( A1 => n719, A2 => n2106, B1 => n2100, B2 => n863, 
                           ZN => n1508);
   U161 : OAI22_X1 port map( A1 => n722, A2 => n2106, B1 => n2100, B2 => n865, 
                           ZN => n1506);
   U162 : OAI22_X1 port map( A1 => n725, A2 => n2106, B1 => n2100, B2 => n867, 
                           ZN => n1504);
   U163 : OAI22_X1 port map( A1 => n728, A2 => n2106, B1 => n2100, B2 => n871, 
                           ZN => n1502);
   U164 : AND3_X1 port map( A1 => n2173, A2 => n2174, A3 => n2164, ZN => n526);
   U165 : AND3_X1 port map( A1 => n2164, A2 => n2174, A3 => ADD_RD1(0), ZN => 
                           n527);
   U166 : AND3_X1 port map( A1 => n2164, A2 => n2173, A3 => ADD_RD1(1), ZN => 
                           n525);
   U167 : NAND2_X1 port map( A1 => n734, A2 => n2106, ZN => n742);
   U168 : AND3_X1 port map( A1 => n2135, A2 => n2172, A3 => ADD_RD2(0), ZN => 
                           n740);
   U169 : AND3_X1 port map( A1 => n2135, A2 => n2171, A3 => ADD_RD2(1), ZN => 
                           n738);
   U170 : AND3_X1 port map( A1 => n2171, A2 => n2172, A3 => n2135, ZN => n739);
   U171 : AND2_X1 port map( A1 => RD2, A2 => n734, ZN => n736);
   U172 : AND2_X1 port map( A1 => RD1, A2 => n734, ZN => n523);
   U173 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n873);
   U174 : OAI221_X1 port map( B1 => n2169, B2 => n562, C1 => n1937, C2 => n2160
                           , A => n563, ZN => n1681);
   U175 : AOI222_X1 port map( A1 => n52, A2 => n2153, B1 => n180, B2 => n2149, 
                           C1 => n2146, C2 => n564, ZN => n563);
   U176 : OAI221_X1 port map( B1 => n2169, B2 => n565, C1 => n1936, C2 => n2160
                           , A => n566, ZN => n1680);
   U177 : AOI222_X1 port map( A1 => n51, A2 => n2154, B1 => n179, B2 => n2149, 
                           C1 => n2146, C2 => n567, ZN => n566);
   U178 : OAI221_X1 port map( B1 => n2169, B2 => n568, C1 => n1935, C2 => n2160
                           , A => n569, ZN => n1679);
   U179 : AOI222_X1 port map( A1 => n50, A2 => n2154, B1 => n178, B2 => n2149, 
                           C1 => n2146, C2 => n570, ZN => n569);
   U180 : OAI221_X1 port map( B1 => n2169, B2 => n571, C1 => n1934, C2 => n2161
                           , A => n572, ZN => n1678);
   U181 : AOI222_X1 port map( A1 => n49, A2 => n2154, B1 => n177, B2 => n2149, 
                           C1 => n2145, C2 => n573, ZN => n572);
   U182 : OAI221_X1 port map( B1 => n2168, B2 => n574, C1 => n1933, C2 => n2160
                           , A => n575, ZN => n1677);
   U183 : AOI222_X1 port map( A1 => n48, A2 => n2154, B1 => n176, B2 => n2149, 
                           C1 => n2145, C2 => n576, ZN => n575);
   U184 : OAI221_X1 port map( B1 => n2168, B2 => n577, C1 => n1932, C2 => n2160
                           , A => n578, ZN => n1676);
   U185 : AOI222_X1 port map( A1 => n47, A2 => n2154, B1 => n175, B2 => n2149, 
                           C1 => n2145, C2 => n579, ZN => n578);
   U186 : OAI221_X1 port map( B1 => n2168, B2 => n580, C1 => n1931, C2 => n2160
                           , A => n581, ZN => n1675);
   U187 : AOI222_X1 port map( A1 => n46, A2 => n2154, B1 => n174, B2 => n2149, 
                           C1 => n2145, C2 => n582, ZN => n581);
   U188 : OAI221_X1 port map( B1 => n538, B2 => n2140, C1 => n1881, C2 => n2130
                           , A => n750, ZN => n1621);
   U189 : AOI222_X1 port map( A1 => n2128, A2 => n60, B1 => n2122, B2 => n188, 
                           C1 => n2116, C2 => n540, ZN => n750);
   U190 : OAI221_X1 port map( B1 => n541, B2 => n2140, C1 => n1880, C2 => n2130
                           , A => n752, ZN => n1619);
   U191 : AOI222_X1 port map( A1 => n2128, A2 => n59, B1 => n2122, B2 => n187, 
                           C1 => n2116, C2 => n543, ZN => n752);
   U192 : OAI221_X1 port map( B1 => n544, B2 => n2140, C1 => n1879, C2 => n2130
                           , A => n754, ZN => n1617);
   U193 : AOI222_X1 port map( A1 => n2128, A2 => n58, B1 => n2122, B2 => n186, 
                           C1 => n2116, C2 => n546, ZN => n754);
   U194 : OAI221_X1 port map( B1 => n547, B2 => n2140, C1 => n1878, C2 => n2130
                           , A => n756, ZN => n1615);
   U195 : AOI222_X1 port map( A1 => n2128, A2 => n57, B1 => n2122, B2 => n185, 
                           C1 => n2116, C2 => n549, ZN => n756);
   U196 : OAI221_X1 port map( B1 => n550, B2 => n2140, C1 => n1877, C2 => n2130
                           , A => n758, ZN => n1613);
   U197 : AOI222_X1 port map( A1 => n2128, A2 => n56, B1 => n2122, B2 => n184, 
                           C1 => n2116, C2 => n552, ZN => n758);
   U198 : OAI221_X1 port map( B1 => n553, B2 => n2140, C1 => n1876, C2 => n2130
                           , A => n760, ZN => n1611);
   U199 : AOI222_X1 port map( A1 => n2128, A2 => n55, B1 => n2122, B2 => n183, 
                           C1 => n2116, C2 => n555, ZN => n760);
   U200 : OAI221_X1 port map( B1 => n556, B2 => n2140, C1 => n1875, C2 => n2130
                           , A => n762, ZN => n1609);
   U201 : AOI222_X1 port map( A1 => n2128, A2 => n54, B1 => n2122, B2 => n182, 
                           C1 => n2116, C2 => n558, ZN => n762);
   U202 : OAI221_X1 port map( B1 => n559, B2 => n2140, C1 => n1874, C2 => n2130
                           , A => n764, ZN => n1607);
   U203 : AOI222_X1 port map( A1 => n2128, A2 => n53, B1 => n2122, B2 => n181, 
                           C1 => n2116, C2 => n561, ZN => n764);
   U204 : OAI221_X1 port map( B1 => n562, B2 => n2140, C1 => n1873, C2 => n2131
                           , A => n766, ZN => n1605);
   U205 : AOI222_X1 port map( A1 => n2128, A2 => n52, B1 => n2122, B2 => n180, 
                           C1 => n2116, C2 => n564, ZN => n766);
   U206 : OAI221_X1 port map( B1 => n565, B2 => n2140, C1 => n1872, C2 => n2131
                           , A => n768, ZN => n1603);
   U207 : AOI222_X1 port map( A1 => n2128, A2 => n51, B1 => n2122, B2 => n179, 
                           C1 => n2116, C2 => n567, ZN => n768);
   U208 : OAI221_X1 port map( B1 => n568, B2 => n2140, C1 => n1871, C2 => n2131
                           , A => n770, ZN => n1601);
   U209 : AOI222_X1 port map( A1 => n2128, A2 => n50, B1 => n2122, B2 => n178, 
                           C1 => n2116, C2 => n570, ZN => n770);
   U210 : OAI221_X1 port map( B1 => n571, B2 => n2140, C1 => n1870, C2 => n2132
                           , A => n772, ZN => n1599);
   U211 : AOI222_X1 port map( A1 => n2128, A2 => n49, B1 => n2122, B2 => n177, 
                           C1 => n2116, C2 => n573, ZN => n772);
   U212 : OAI221_X1 port map( B1 => n574, B2 => n2139, C1 => n1869, C2 => n2131
                           , A => n774, ZN => n1597);
   U213 : AOI222_X1 port map( A1 => n2127, A2 => n48, B1 => n2121, B2 => n176, 
                           C1 => n2115, C2 => n576, ZN => n774);
   U214 : OAI221_X1 port map( B1 => n577, B2 => n2139, C1 => n1868, C2 => n2131
                           , A => n776, ZN => n1595);
   U215 : AOI222_X1 port map( A1 => n2127, A2 => n47, B1 => n2121, B2 => n175, 
                           C1 => n2115, C2 => n579, ZN => n776);
   U216 : OAI221_X1 port map( B1 => n580, B2 => n2139, C1 => n1867, C2 => n2131
                           , A => n778, ZN => n1593);
   U217 : AOI222_X1 port map( A1 => n2127, A2 => n46, B1 => n2121, B2 => n174, 
                           C1 => n2115, C2 => n582, ZN => n778);
   U218 : OAI221_X1 port map( B1 => n2165, B2 => n716, C1 => n1890, C2 => n2164
                           , A => n717, ZN => n1634);
   U219 : AOI222_X1 port map( A1 => n5, A2 => n2157, B1 => n2152, B2 => n718, 
                           C1 => n69, C2 => n2142, ZN => n717);
   U220 : OAI221_X1 port map( B1 => n2165, B2 => n722, C1 => n1888, C2 => n2164
                           , A => n723, ZN => n1632);
   U221 : AOI222_X1 port map( A1 => n3, A2 => n2157, B1 => n2152, B2 => n724, 
                           C1 => n67, C2 => n2142, ZN => n723);
   U222 : OAI221_X1 port map( B1 => n2165, B2 => n725, C1 => n1887, C2 => n2164
                           , A => n726, ZN => n1631);
   U223 : AOI222_X1 port map( A1 => n2, A2 => n2157, B1 => n2152, B2 => n727, 
                           C1 => n66, C2 => n2142, ZN => n726);
   U224 : OAI221_X1 port map( B1 => n2165, B2 => n728, C1 => n1886, C2 => n2164
                           , A => n729, ZN => n1630);
   U225 : AOI222_X1 port map( A1 => n2158, A2 => n730, B1 => n2150, B2 => n731,
                           C1 => n65, C2 => n2142, ZN => n729);
   U226 : OAI221_X1 port map( B1 => n623, B2 => n2138, C1 => n1856, C2 => n2132
                           , A => n800, ZN => n1571);
   U227 : AOI222_X1 port map( A1 => n2126, A2 => n35, B1 => n2120, B2 => n625, 
                           C1 => n2114, C2 => n99, ZN => n800);
   U228 : OAI221_X1 port map( B1 => n626, B2 => n2138, C1 => n1855, C2 => n2132
                           , A => n802, ZN => n1569);
   U229 : AOI222_X1 port map( A1 => n2126, A2 => n34, B1 => n2120, B2 => n628, 
                           C1 => n2114, C2 => n98, ZN => n802);
   U230 : OAI221_X1 port map( B1 => n629, B2 => n2138, C1 => n1854, C2 => n2132
                           , A => n804, ZN => n1567);
   U231 : AOI222_X1 port map( A1 => n2126, A2 => n33, B1 => n2120, B2 => n631, 
                           C1 => n2114, C2 => n97, ZN => n804);
   U232 : OAI221_X1 port map( B1 => n632, B2 => n2138, C1 => n1853, C2 => n2132
                           , A => n806, ZN => n1565);
   U233 : AOI222_X1 port map( A1 => n2126, A2 => n32, B1 => n2120, B2 => n634, 
                           C1 => n2114, C2 => n96, ZN => n806);
   U234 : OAI221_X1 port map( B1 => n635, B2 => n2138, C1 => n1852, C2 => n2132
                           , A => n808, ZN => n1563);
   U235 : AOI222_X1 port map( A1 => n2126, A2 => n31, B1 => n2120, B2 => n637, 
                           C1 => n2114, C2 => n95, ZN => n808);
   U236 : OAI221_X1 port map( B1 => n638, B2 => n2138, C1 => n1851, C2 => n2132
                           , A => n810, ZN => n1561);
   U237 : AOI222_X1 port map( A1 => n2126, A2 => n30, B1 => n2120, B2 => n640, 
                           C1 => n2114, C2 => n94, ZN => n810);
   U238 : OAI221_X1 port map( B1 => n641, B2 => n2138, C1 => n1850, C2 => n2132
                           , A => n812, ZN => n1559);
   U239 : AOI222_X1 port map( A1 => n2126, A2 => n29, B1 => n2120, B2 => n643, 
                           C1 => n2114, C2 => n93, ZN => n812);
   U240 : OAI221_X1 port map( B1 => n644, B2 => n2138, C1 => n1849, C2 => n2133
                           , A => n814, ZN => n1557);
   U241 : AOI222_X1 port map( A1 => n2126, A2 => n28, B1 => n2120, B2 => n646, 
                           C1 => n2114, C2 => n92, ZN => n814);
   U242 : OAI221_X1 port map( B1 => n647, B2 => n2138, C1 => n1848, C2 => n2133
                           , A => n816, ZN => n1555);
   U243 : AOI222_X1 port map( A1 => n2126, A2 => n27, B1 => n2120, B2 => n649, 
                           C1 => n2114, C2 => n91, ZN => n816);
   U244 : OAI221_X1 port map( B1 => n650, B2 => n2138, C1 => n1847, C2 => n2133
                           , A => n818, ZN => n1553);
   U245 : AOI222_X1 port map( A1 => n2126, A2 => n26, B1 => n2120, B2 => n652, 
                           C1 => n2114, C2 => n90, ZN => n818);
   U246 : OAI221_X1 port map( B1 => n653, B2 => n2138, C1 => n1846, C2 => n2133
                           , A => n820, ZN => n1551);
   U247 : AOI222_X1 port map( A1 => n2126, A2 => n25, B1 => n2120, B2 => n655, 
                           C1 => n2114, C2 => n89, ZN => n820);
   U248 : OAI221_X1 port map( B1 => n656, B2 => n2137, C1 => n1845, C2 => n2133
                           , A => n822, ZN => n1549);
   U249 : AOI222_X1 port map( A1 => n2125, A2 => n24, B1 => n2119, B2 => n658, 
                           C1 => n2113, C2 => n88, ZN => n822);
   U250 : OAI221_X1 port map( B1 => n659, B2 => n2137, C1 => n1844, C2 => n2133
                           , A => n824, ZN => n1547);
   U251 : AOI222_X1 port map( A1 => n2125, A2 => n23, B1 => n2119, B2 => n661, 
                           C1 => n2113, C2 => n87, ZN => n824);
   U252 : OAI221_X1 port map( B1 => n662, B2 => n2137, C1 => n1843, C2 => n2133
                           , A => n826, ZN => n1545);
   U253 : AOI222_X1 port map( A1 => n2125, A2 => n22, B1 => n2119, B2 => n664, 
                           C1 => n2113, C2 => n86, ZN => n826);
   U254 : OAI221_X1 port map( B1 => n665, B2 => n2137, C1 => n1842, C2 => n2133
                           , A => n828, ZN => n1543);
   U255 : AOI222_X1 port map( A1 => n2125, A2 => n21, B1 => n2119, B2 => n667, 
                           C1 => n2113, C2 => n85, ZN => n828);
   U256 : OAI221_X1 port map( B1 => n668, B2 => n2137, C1 => n1841, C2 => n2133
                           , A => n830, ZN => n1541);
   U257 : AOI222_X1 port map( A1 => n2125, A2 => n20, B1 => n2119, B2 => n670, 
                           C1 => n2113, C2 => n84, ZN => n830);
   U258 : OAI221_X1 port map( B1 => n671, B2 => n2137, C1 => n1840, C2 => n2133
                           , A => n832, ZN => n1539);
   U259 : AOI222_X1 port map( A1 => n2125, A2 => n19, B1 => n2119, B2 => n673, 
                           C1 => n2113, C2 => n83, ZN => n832);
   U260 : OAI221_X1 port map( B1 => n674, B2 => n2137, C1 => n1839, C2 => n2133
                           , A => n834, ZN => n1537);
   U261 : AOI222_X1 port map( A1 => n2125, A2 => n18, B1 => n2119, B2 => n676, 
                           C1 => n2113, C2 => n82, ZN => n834);
   U262 : OAI221_X1 port map( B1 => n677, B2 => n2137, C1 => n1838, C2 => n2133
                           , A => n836, ZN => n1535);
   U263 : AOI222_X1 port map( A1 => n2125, A2 => n17, B1 => n2119, B2 => n679, 
                           C1 => n2113, C2 => n81, ZN => n836);
   U264 : OAI221_X1 port map( B1 => n680, B2 => n2137, C1 => n1837, C2 => n2134
                           , A => n838, ZN => n1533);
   U265 : AOI222_X1 port map( A1 => n2125, A2 => n16, B1 => n2119, B2 => n682, 
                           C1 => n2113, C2 => n80, ZN => n838);
   U266 : OAI221_X1 port map( B1 => n683, B2 => n2137, C1 => n1836, C2 => n2134
                           , A => n840, ZN => n1531);
   U267 : AOI222_X1 port map( A1 => n2125, A2 => n15, B1 => n2119, B2 => n685, 
                           C1 => n2113, C2 => n79, ZN => n840);
   U268 : OAI221_X1 port map( B1 => n686, B2 => n2137, C1 => n1835, C2 => n2134
                           , A => n842, ZN => n1529);
   U269 : AOI222_X1 port map( A1 => n2125, A2 => n14, B1 => n2119, B2 => n688, 
                           C1 => n2113, C2 => n78, ZN => n842);
   U270 : OAI221_X1 port map( B1 => n689, B2 => n2137, C1 => n1834, C2 => n2134
                           , A => n844, ZN => n1527);
   U271 : AOI222_X1 port map( A1 => n2125, A2 => n13, B1 => n2119, B2 => n691, 
                           C1 => n2113, C2 => n77, ZN => n844);
   U272 : OAI221_X1 port map( B1 => n692, B2 => n2136, C1 => n1833, C2 => n2134
                           , A => n846, ZN => n1525);
   U273 : AOI222_X1 port map( A1 => n2124, A2 => n694, B1 => n2118, B2 => n695,
                           C1 => n2112, C2 => n76, ZN => n846);
   U274 : OAI221_X1 port map( B1 => n696, B2 => n2136, C1 => n1832, C2 => n2134
                           , A => n848, ZN => n1523);
   U275 : AOI222_X1 port map( A1 => n2124, A2 => n698, B1 => n2118, B2 => n699,
                           C1 => n2112, C2 => n75, ZN => n848);
   U276 : OAI221_X1 port map( B1 => n700, B2 => n2136, C1 => n1831, C2 => n2134
                           , A => n850, ZN => n1521);
   U277 : AOI222_X1 port map( A1 => n2124, A2 => n702, B1 => n2118, B2 => n703,
                           C1 => n2112, C2 => n74, ZN => n850);
   U278 : OAI221_X1 port map( B1 => n704, B2 => n2136, C1 => n1830, C2 => n2134
                           , A => n852, ZN => n1519);
   U279 : AOI222_X1 port map( A1 => n2124, A2 => n9, B1 => n2118, B2 => n706, 
                           C1 => n2112, C2 => n73, ZN => n852);
   U280 : OAI221_X1 port map( B1 => n707, B2 => n2136, C1 => n1829, C2 => n2134
                           , A => n854, ZN => n1517);
   U281 : AOI222_X1 port map( A1 => n2124, A2 => n8, B1 => n2118, B2 => n709, 
                           C1 => n2112, C2 => n72, ZN => n854);
   U282 : OAI221_X1 port map( B1 => n710, B2 => n2136, C1 => n1828, C2 => n2134
                           , A => n856, ZN => n1515);
   U283 : AOI222_X1 port map( A1 => n2124, A2 => n7, B1 => n2118, B2 => n712, 
                           C1 => n2112, C2 => n71, ZN => n856);
   U284 : OAI221_X1 port map( B1 => n713, B2 => n2136, C1 => n1827, C2 => n2134
                           , A => n858, ZN => n1513);
   U285 : AOI222_X1 port map( A1 => n2124, A2 => n6, B1 => n2118, B2 => n715, 
                           C1 => n2112, C2 => n70, ZN => n858);
   U286 : OAI221_X1 port map( B1 => n716, B2 => n2136, C1 => n1826, C2 => n2135
                           , A => n860, ZN => n1511);
   U287 : AOI222_X1 port map( A1 => n2124, A2 => n5, B1 => n2118, B2 => n718, 
                           C1 => n2112, C2 => n69, ZN => n860);
   U288 : OAI221_X1 port map( B1 => n719, B2 => n2136, C1 => n1825, C2 => n2134
                           , A => n862, ZN => n1509);
   U289 : AOI222_X1 port map( A1 => n2124, A2 => n4, B1 => n2118, B2 => n721, 
                           C1 => n2112, C2 => n68, ZN => n862);
   U290 : OAI221_X1 port map( B1 => n722, B2 => n2136, C1 => n1824, C2 => n2135
                           , A => n864, ZN => n1507);
   U291 : AOI222_X1 port map( A1 => n2124, A2 => n3, B1 => n2118, B2 => n724, 
                           C1 => n2112, C2 => n67, ZN => n864);
   U292 : OAI221_X1 port map( B1 => n725, B2 => n2136, C1 => n1823, C2 => n2135
                           , A => n866, ZN => n1505);
   U293 : AOI222_X1 port map( A1 => n2124, A2 => n2, B1 => n2118, B2 => n727, 
                           C1 => n2112, C2 => n66, ZN => n866);
   U294 : OAI221_X1 port map( B1 => n728, B2 => n2136, C1 => n1822, C2 => n2135
                           , A => n868, ZN => n1503);
   U295 : AOI222_X1 port map( A1 => n2124, A2 => n730, B1 => n2118, B2 => n731,
                           C1 => n2112, C2 => n65, ZN => n868);
   U296 : INV_X1 port map( A => RESET, ZN => n734);
   U297 : OAI221_X1 port map( B1 => n2170, B2 => n522, C1 => n1949, C2 => n2159
                           , A => n524, ZN => n1693);
   U298 : AOI222_X1 port map( A1 => n64, A2 => n2155, B1 => n192, B2 => n2148, 
                           C1 => n2147, C2 => n528, ZN => n524);
   U299 : OAI221_X1 port map( B1 => n2170, B2 => n529, C1 => n1948, C2 => n2159
                           , A => n530, ZN => n1692);
   U300 : AOI222_X1 port map( A1 => n63, A2 => n2153, B1 => n191, B2 => n2148, 
                           C1 => n2147, C2 => n531, ZN => n530);
   U301 : OAI221_X1 port map( B1 => n2170, B2 => n532, C1 => n1947, C2 => n2159
                           , A => n533, ZN => n1691);
   U302 : AOI222_X1 port map( A1 => n62, A2 => n2153, B1 => n190, B2 => n2148, 
                           C1 => n2146, C2 => n534, ZN => n533);
   U303 : OAI221_X1 port map( B1 => n2170, B2 => n535, C1 => n1946, C2 => n2159
                           , A => n536, ZN => n1690);
   U304 : AOI222_X1 port map( A1 => n61, A2 => n2153, B1 => n189, B2 => n2148, 
                           C1 => n2146, C2 => n537, ZN => n536);
   U305 : OAI221_X1 port map( B1 => n2167, B2 => n619, C1 => n1921, C2 => n2161
                           , A => n620, ZN => n1665);
   U306 : AOI222_X1 port map( A1 => n36, A2 => n2155, B1 => n2150, B2 => n621, 
                           C1 => n2144, C2 => n622, ZN => n620);
   U307 : OAI221_X1 port map( B1 => n2167, B2 => n623, C1 => n1920, C2 => n2161
                           , A => n624, ZN => n1664);
   U308 : AOI222_X1 port map( A1 => n35, A2 => n2155, B1 => n2150, B2 => n625, 
                           C1 => n99, C2 => n2144, ZN => n624);
   U309 : OAI221_X1 port map( B1 => n2167, B2 => n626, C1 => n1919, C2 => n2161
                           , A => n627, ZN => n1663);
   U310 : AOI222_X1 port map( A1 => n34, A2 => n2155, B1 => n2150, B2 => n628, 
                           C1 => n98, C2 => n2144, ZN => n627);
   U311 : OAI221_X1 port map( B1 => n2167, B2 => n629, C1 => n1918, C2 => n2161
                           , A => n630, ZN => n1662);
   U312 : AOI222_X1 port map( A1 => n33, A2 => n2155, B1 => n2150, B2 => n631, 
                           C1 => n97, C2 => n2144, ZN => n630);
   U313 : OAI221_X1 port map( B1 => n2167, B2 => n632, C1 => n1917, C2 => n2161
                           , A => n633, ZN => n1661);
   U314 : AOI222_X1 port map( A1 => n32, A2 => n2155, B1 => n2150, B2 => n634, 
                           C1 => n96, C2 => n2144, ZN => n633);
   U315 : OAI221_X1 port map( B1 => n2167, B2 => n635, C1 => n1916, C2 => n2161
                           , A => n636, ZN => n1660);
   U316 : AOI222_X1 port map( A1 => n31, A2 => n2155, B1 => n2150, B2 => n637, 
                           C1 => n95, C2 => n2144, ZN => n636);
   U317 : OAI221_X1 port map( B1 => n2167, B2 => n638, C1 => n1915, C2 => n2161
                           , A => n639, ZN => n1659);
   U318 : AOI222_X1 port map( A1 => n30, A2 => n2155, B1 => n2150, B2 => n640, 
                           C1 => n94, C2 => n2144, ZN => n639);
   U319 : OAI221_X1 port map( B1 => n2167, B2 => n641, C1 => n1914, C2 => n2161
                           , A => n642, ZN => n1658);
   U320 : AOI222_X1 port map( A1 => n29, A2 => n2155, B1 => n2150, B2 => n643, 
                           C1 => n93, C2 => n2144, ZN => n642);
   U321 : OAI221_X1 port map( B1 => n2167, B2 => n644, C1 => n1913, C2 => n2162
                           , A => n645, ZN => n1657);
   U322 : AOI222_X1 port map( A1 => n28, A2 => n2156, B1 => n2150, B2 => n646, 
                           C1 => n92, C2 => n2144, ZN => n645);
   U323 : OAI221_X1 port map( B1 => n2167, B2 => n647, C1 => n1912, C2 => n2162
                           , A => n648, ZN => n1656);
   U324 : AOI222_X1 port map( A1 => n27, A2 => n2156, B1 => n2151, B2 => n649, 
                           C1 => n91, C2 => n2144, ZN => n648);
   U325 : OAI221_X1 port map( B1 => n2167, B2 => n650, C1 => n1911, C2 => n2162
                           , A => n651, ZN => n1655);
   U326 : AOI222_X1 port map( A1 => n26, A2 => n2156, B1 => n2151, B2 => n652, 
                           C1 => n90, C2 => n2144, ZN => n651);
   U327 : OAI221_X1 port map( B1 => n2167, B2 => n653, C1 => n1910, C2 => n2162
                           , A => n654, ZN => n1654);
   U328 : AOI222_X1 port map( A1 => n25, A2 => n2156, B1 => n2151, B2 => n655, 
                           C1 => n89, C2 => n2144, ZN => n654);
   U329 : OAI221_X1 port map( B1 => n2166, B2 => n656, C1 => n1909, C2 => n2162
                           , A => n657, ZN => n1653);
   U330 : AOI222_X1 port map( A1 => n24, A2 => n2156, B1 => n2151, B2 => n658, 
                           C1 => n88, C2 => n2143, ZN => n657);
   U331 : OAI221_X1 port map( B1 => n2166, B2 => n659, C1 => n1908, C2 => n2162
                           , A => n660, ZN => n1652);
   U332 : AOI222_X1 port map( A1 => n23, A2 => n2156, B1 => n2151, B2 => n661, 
                           C1 => n87, C2 => n2143, ZN => n660);
   U333 : OAI221_X1 port map( B1 => n2166, B2 => n662, C1 => n1907, C2 => n2162
                           , A => n663, ZN => n1651);
   U334 : AOI222_X1 port map( A1 => n22, A2 => n2156, B1 => n2151, B2 => n664, 
                           C1 => n86, C2 => n2143, ZN => n663);
   U335 : OAI221_X1 port map( B1 => n2166, B2 => n665, C1 => n1906, C2 => n2162
                           , A => n666, ZN => n1650);
   U336 : AOI222_X1 port map( A1 => n21, A2 => n2156, B1 => n2151, B2 => n667, 
                           C1 => n85, C2 => n2143, ZN => n666);
   U337 : OAI221_X1 port map( B1 => n2166, B2 => n668, C1 => n1905, C2 => n2162
                           , A => n669, ZN => n1649);
   U338 : AOI222_X1 port map( A1 => n20, A2 => n2156, B1 => n2151, B2 => n670, 
                           C1 => n84, C2 => n2143, ZN => n669);
   U339 : OAI221_X1 port map( B1 => n2166, B2 => n671, C1 => n1904, C2 => n2162
                           , A => n672, ZN => n1648);
   U340 : AOI222_X1 port map( A1 => n19, A2 => n2156, B1 => n2151, B2 => n673, 
                           C1 => n83, C2 => n2143, ZN => n672);
   U341 : OAI221_X1 port map( B1 => n2166, B2 => n674, C1 => n1903, C2 => n2162
                           , A => n675, ZN => n1647);
   U342 : AOI222_X1 port map( A1 => n18, A2 => n2156, B1 => n2151, B2 => n676, 
                           C1 => n82, C2 => n2143, ZN => n675);
   U343 : OAI221_X1 port map( B1 => n2166, B2 => n677, C1 => n1902, C2 => n2162
                           , A => n678, ZN => n1646);
   U344 : AOI222_X1 port map( A1 => n17, A2 => n2156, B1 => n2151, B2 => n679, 
                           C1 => n81, C2 => n2143, ZN => n678);
   U345 : OAI221_X1 port map( B1 => n2166, B2 => n680, C1 => n1901, C2 => n2163
                           , A => n681, ZN => n1645);
   U346 : AOI222_X1 port map( A1 => n16, A2 => n2157, B1 => n2151, B2 => n682, 
                           C1 => n80, C2 => n2143, ZN => n681);
   U347 : OAI221_X1 port map( B1 => n2166, B2 => n683, C1 => n1900, C2 => n2163
                           , A => n684, ZN => n1644);
   U348 : AOI222_X1 port map( A1 => n15, A2 => n2157, B1 => n2151, B2 => n685, 
                           C1 => n79, C2 => n2143, ZN => n684);
   U349 : OAI221_X1 port map( B1 => n2166, B2 => n686, C1 => n1899, C2 => n2163
                           , A => n687, ZN => n1643);
   U350 : AOI222_X1 port map( A1 => n14, A2 => n2157, B1 => n2152, B2 => n688, 
                           C1 => n78, C2 => n2143, ZN => n687);
   U351 : OAI221_X1 port map( B1 => n2166, B2 => n689, C1 => n1898, C2 => n2163
                           , A => n690, ZN => n1642);
   U352 : AOI222_X1 port map( A1 => n13, A2 => n2157, B1 => n2152, B2 => n691, 
                           C1 => n77, C2 => n2143, ZN => n690);
   U353 : OAI221_X1 port map( B1 => n2165, B2 => n692, C1 => n1897, C2 => n2163
                           , A => n693, ZN => n1641);
   U354 : AOI222_X1 port map( A1 => n2158, A2 => n694, B1 => n2152, B2 => n695,
                           C1 => n76, C2 => n2142, ZN => n693);
   U355 : OAI221_X1 port map( B1 => n2165, B2 => n696, C1 => n1896, C2 => n2163
                           , A => n697, ZN => n1640);
   U356 : AOI222_X1 port map( A1 => n2158, A2 => n698, B1 => n2152, B2 => n699,
                           C1 => n75, C2 => n2142, ZN => n697);
   U357 : OAI221_X1 port map( B1 => n2165, B2 => n700, C1 => n1895, C2 => n2163
                           , A => n701, ZN => n1639);
   U358 : AOI222_X1 port map( A1 => n2158, A2 => n702, B1 => n2152, B2 => n703,
                           C1 => n74, C2 => n2142, ZN => n701);
   U359 : OAI221_X1 port map( B1 => n2165, B2 => n704, C1 => n1894, C2 => n2163
                           , A => n705, ZN => n1638);
   U360 : AOI222_X1 port map( A1 => n9, A2 => n2157, B1 => n2152, B2 => n706, 
                           C1 => n73, C2 => n2142, ZN => n705);
   U361 : OAI221_X1 port map( B1 => n2165, B2 => n707, C1 => n1893, C2 => n2163
                           , A => n708, ZN => n1637);
   U362 : AOI222_X1 port map( A1 => n8, A2 => n2157, B1 => n2152, B2 => n709, 
                           C1 => n72, C2 => n2142, ZN => n708);
   U363 : OAI221_X1 port map( B1 => n2165, B2 => n710, C1 => n1892, C2 => n2163
                           , A => n711, ZN => n1636);
   U364 : AOI222_X1 port map( A1 => n7, A2 => n2157, B1 => n2152, B2 => n712, 
                           C1 => n71, C2 => n2142, ZN => n711);
   U365 : OAI221_X1 port map( B1 => n2165, B2 => n713, C1 => n1891, C2 => n2163
                           , A => n714, ZN => n1635);
   U366 : AOI222_X1 port map( A1 => n6, A2 => n2157, B1 => n2152, B2 => n715, 
                           C1 => n70, C2 => n2142, ZN => n714);
   U367 : OAI221_X1 port map( B1 => n2165, B2 => n719, C1 => n1889, C2 => n2163
                           , A => n720, ZN => n1633);
   U368 : AOI222_X1 port map( A1 => n4, A2 => n2157, B1 => n2152, B2 => n721, 
                           C1 => n68, C2 => n2142, ZN => n720);
   U369 : OAI221_X1 port map( B1 => n522, B2 => n2141, C1 => n1885, C2 => n2130
                           , A => n737, ZN => n1629);
   U370 : AOI222_X1 port map( A1 => n2129, A2 => n64, B1 => n2123, B2 => n192, 
                           C1 => n2117, C2 => n528, ZN => n737);
   U371 : OAI221_X1 port map( B1 => n529, B2 => n2141, C1 => n1884, C2 => n2130
                           , A => n744, ZN => n1627);
   U372 : AOI222_X1 port map( A1 => n2129, A2 => n63, B1 => n2123, B2 => n191, 
                           C1 => n2117, C2 => n531, ZN => n744);
   U373 : OAI221_X1 port map( B1 => n532, B2 => n2141, C1 => n1883, C2 => n2130
                           , A => n746, ZN => n1625);
   U374 : AOI222_X1 port map( A1 => n2129, A2 => n62, B1 => n2123, B2 => n190, 
                           C1 => n2117, C2 => n534, ZN => n746);
   U375 : OAI221_X1 port map( B1 => n535, B2 => n2141, C1 => n1882, C2 => n2130
                           , A => n748, ZN => n1623);
   U376 : AOI222_X1 port map( A1 => n2129, A2 => n61, B1 => n2123, B2 => n189, 
                           C1 => n2117, C2 => n537, ZN => n748);
   U377 : OAI221_X1 port map( B1 => n583, B2 => n2139, C1 => n1866, C2 => n2131
                           , A => n780, ZN => n1591);
   U378 : AOI222_X1 port map( A1 => n2127, A2 => n45, B1 => n2121, B2 => n585, 
                           C1 => n2115, C2 => n586, ZN => n780);
   U379 : OAI221_X1 port map( B1 => n587, B2 => n2139, C1 => n1865, C2 => n2131
                           , A => n782, ZN => n1589);
   U380 : AOI222_X1 port map( A1 => n2127, A2 => n44, B1 => n2121, B2 => n589, 
                           C1 => n2115, C2 => n590, ZN => n782);
   U381 : OAI221_X1 port map( B1 => n591, B2 => n2139, C1 => n1864, C2 => n2131
                           , A => n784, ZN => n1587);
   U382 : AOI222_X1 port map( A1 => n2127, A2 => n43, B1 => n2121, B2 => n593, 
                           C1 => n2115, C2 => n594, ZN => n784);
   U383 : OAI221_X1 port map( B1 => n595, B2 => n2139, C1 => n1863, C2 => n2131
                           , A => n786, ZN => n1585);
   U384 : AOI222_X1 port map( A1 => n2127, A2 => n42, B1 => n2121, B2 => n597, 
                           C1 => n2115, C2 => n598, ZN => n786);
   U385 : OAI221_X1 port map( B1 => n599, B2 => n2139, C1 => n1862, C2 => n2131
                           , A => n788, ZN => n1583);
   U386 : AOI222_X1 port map( A1 => n2127, A2 => n41, B1 => n2121, B2 => n601, 
                           C1 => n2115, C2 => n602, ZN => n788);
   U387 : OAI221_X1 port map( B1 => n603, B2 => n2139, C1 => n1861, C2 => n2131
                           , A => n790, ZN => n1581);
   U388 : AOI222_X1 port map( A1 => n2127, A2 => n40, B1 => n2121, B2 => n605, 
                           C1 => n2115, C2 => n606, ZN => n790);
   U389 : OAI221_X1 port map( B1 => n607, B2 => n2139, C1 => n1860, C2 => n2132
                           , A => n792, ZN => n1579);
   U390 : AOI222_X1 port map( A1 => n2127, A2 => n39, B1 => n2121, B2 => n609, 
                           C1 => n2115, C2 => n610, ZN => n792);
   U391 : OAI221_X1 port map( B1 => n611, B2 => n2139, C1 => n1859, C2 => n2132
                           , A => n794, ZN => n1577);
   U392 : AOI222_X1 port map( A1 => n2127, A2 => n38, B1 => n2121, B2 => n613, 
                           C1 => n2115, C2 => n614, ZN => n794);
   U393 : OAI221_X1 port map( B1 => n615, B2 => n2139, C1 => n1858, C2 => n2132
                           , A => n796, ZN => n1575);
   U394 : AOI222_X1 port map( A1 => n2127, A2 => n37, B1 => n2121, B2 => n617, 
                           C1 => n2115, C2 => n618, ZN => n796);
   U395 : OAI221_X1 port map( B1 => n619, B2 => n2138, C1 => n1857, C2 => n2132
                           , A => n798, ZN => n1573);
   U396 : AOI222_X1 port map( A1 => n2126, A2 => n36, B1 => n2120, B2 => n621, 
                           C1 => n2114, C2 => n622, ZN => n798);
   U397 : OAI221_X1 port map( B1 => n2169, B2 => n538, C1 => n1945, C2 => n2159
                           , A => n539, ZN => n1689);
   U398 : AOI222_X1 port map( A1 => n60, A2 => n2153, B1 => n188, B2 => n2148, 
                           C1 => n2146, C2 => n540, ZN => n539);
   U399 : OAI221_X1 port map( B1 => n2169, B2 => n541, C1 => n1944, C2 => n2159
                           , A => n542, ZN => n1688);
   U400 : AOI222_X1 port map( A1 => n59, A2 => n2153, B1 => n187, B2 => n2148, 
                           C1 => n2146, C2 => n543, ZN => n542);
   U401 : OAI221_X1 port map( B1 => n2169, B2 => n544, C1 => n1943, C2 => n2159
                           , A => n545, ZN => n1687);
   U402 : AOI222_X1 port map( A1 => n58, A2 => n2153, B1 => n186, B2 => n2148, 
                           C1 => n2146, C2 => n546, ZN => n545);
   U403 : OAI221_X1 port map( B1 => n2169, B2 => n547, C1 => n1942, C2 => n2159
                           , A => n548, ZN => n1686);
   U404 : AOI222_X1 port map( A1 => n57, A2 => n2153, B1 => n185, B2 => n2148, 
                           C1 => n2146, C2 => n549, ZN => n548);
   U405 : OAI221_X1 port map( B1 => n2169, B2 => n550, C1 => n1941, C2 => n2159
                           , A => n551, ZN => n1685);
   U406 : AOI222_X1 port map( A1 => n56, A2 => n2153, B1 => n184, B2 => n2148, 
                           C1 => n2146, C2 => n552, ZN => n551);
   U407 : OAI221_X1 port map( B1 => n2169, B2 => n553, C1 => n1940, C2 => n2159
                           , A => n554, ZN => n1684);
   U408 : AOI222_X1 port map( A1 => n55, A2 => n2153, B1 => n183, B2 => n2148, 
                           C1 => n2146, C2 => n555, ZN => n554);
   U409 : OAI221_X1 port map( B1 => n2169, B2 => n556, C1 => n1939, C2 => n2159
                           , A => n557, ZN => n1683);
   U410 : AOI222_X1 port map( A1 => n54, A2 => n2153, B1 => n182, B2 => n2148, 
                           C1 => n2146, C2 => n558, ZN => n557);
   U411 : OAI221_X1 port map( B1 => n2169, B2 => n559, C1 => n1938, C2 => n2159
                           , A => n560, ZN => n1682);
   U412 : AOI222_X1 port map( A1 => n53, A2 => n2153, B1 => n181, B2 => n2148, 
                           C1 => n2146, C2 => n561, ZN => n560);
   U413 : OAI221_X1 port map( B1 => n2168, B2 => n583, C1 => n1930, C2 => n2160
                           , A => n584, ZN => n1674);
   U414 : AOI222_X1 port map( A1 => n45, A2 => n2154, B1 => n2149, B2 => n585, 
                           C1 => n2145, C2 => n586, ZN => n584);
   U415 : OAI221_X1 port map( B1 => n2168, B2 => n587, C1 => n1929, C2 => n2160
                           , A => n588, ZN => n1673);
   U416 : AOI222_X1 port map( A1 => n44, A2 => n2154, B1 => n2149, B2 => n589, 
                           C1 => n2145, C2 => n590, ZN => n588);
   U417 : OAI221_X1 port map( B1 => n2168, B2 => n591, C1 => n1928, C2 => n2160
                           , A => n592, ZN => n1672);
   U418 : AOI222_X1 port map( A1 => n43, A2 => n2154, B1 => n2149, B2 => n593, 
                           C1 => n2145, C2 => n594, ZN => n592);
   U419 : OAI221_X1 port map( B1 => n2168, B2 => n595, C1 => n1927, C2 => n2160
                           , A => n596, ZN => n1671);
   U420 : AOI222_X1 port map( A1 => n42, A2 => n2154, B1 => n2149, B2 => n597, 
                           C1 => n2145, C2 => n598, ZN => n596);
   U421 : OAI221_X1 port map( B1 => n2168, B2 => n599, C1 => n1926, C2 => n2160
                           , A => n600, ZN => n1670);
   U422 : AOI222_X1 port map( A1 => n41, A2 => n2154, B1 => n2149, B2 => n601, 
                           C1 => n2145, C2 => n602, ZN => n600);
   U423 : OAI221_X1 port map( B1 => n2168, B2 => n603, C1 => n1925, C2 => n2160
                           , A => n604, ZN => n1669);
   U424 : AOI222_X1 port map( A1 => n40, A2 => n2154, B1 => n2150, B2 => n605, 
                           C1 => n2145, C2 => n606, ZN => n604);
   U425 : OAI221_X1 port map( B1 => n2168, B2 => n607, C1 => n1924, C2 => n2161
                           , A => n608, ZN => n1668);
   U426 : AOI222_X1 port map( A1 => n39, A2 => n2155, B1 => n2150, B2 => n609, 
                           C1 => n2145, C2 => n610, ZN => n608);
   U427 : OAI221_X1 port map( B1 => n2168, B2 => n611, C1 => n1923, C2 => n2161
                           , A => n612, ZN => n1667);
   U428 : AOI222_X1 port map( A1 => n38, A2 => n2155, B1 => n2150, B2 => n613, 
                           C1 => n2145, C2 => n614, ZN => n612);
   U429 : OAI221_X1 port map( B1 => n2168, B2 => n615, C1 => n1922, C2 => n2161
                           , A => n616, ZN => n1666);
   U430 : AOI222_X1 port map( A1 => n37, A2 => n2155, B1 => n2150, B2 => n617, 
                           C1 => n2145, C2 => n618, ZN => n616);
   U431 : OAI22_X1 port map( A1 => n1950, A2 => n2099, B1 => n743, B2 => n2093,
                           ZN => n1501);
   U432 : OAI22_X1 port map( A1 => n1951, A2 => n2099, B1 => n745, B2 => n2093,
                           ZN => n1500);
   U433 : OAI22_X1 port map( A1 => n1952, A2 => n2099, B1 => n747, B2 => n2093,
                           ZN => n1499);
   U434 : OAI22_X1 port map( A1 => n1953, A2 => n2099, B1 => n749, B2 => n2093,
                           ZN => n1498);
   U435 : OAI22_X1 port map( A1 => n1821, A2 => n2087, B1 => n743, B2 => n2081,
                           ZN => n1437);
   U436 : OAI22_X1 port map( A1 => n1820, A2 => n2087, B1 => n745, B2 => n2081,
                           ZN => n1436);
   U437 : OAI22_X1 port map( A1 => n1819, A2 => n2087, B1 => n747, B2 => n2081,
                           ZN => n1435);
   U438 : OAI22_X1 port map( A1 => n1818, A2 => n2087, B1 => n749, B2 => n2081,
                           ZN => n1434);
   U439 : OAI22_X1 port map( A1 => n2010, A2 => n2075, B1 => n743, B2 => n2069,
                           ZN => n1373);
   U440 : OAI22_X1 port map( A1 => n2011, A2 => n2075, B1 => n745, B2 => n2069,
                           ZN => n1372);
   U441 : OAI22_X1 port map( A1 => n2012, A2 => n2075, B1 => n747, B2 => n2069,
                           ZN => n1371);
   U442 : OAI22_X1 port map( A1 => n2013, A2 => n2075, B1 => n749, B2 => n2069,
                           ZN => n1370);
   U443 : OAI22_X1 port map( A1 => n1954, A2 => n2099, B1 => n751, B2 => n2092,
                           ZN => n1497);
   U444 : OAI22_X1 port map( A1 => n1955, A2 => n2098, B1 => n753, B2 => n2092,
                           ZN => n1496);
   U445 : OAI22_X1 port map( A1 => n1956, A2 => n2098, B1 => n755, B2 => n2092,
                           ZN => n1495);
   U446 : OAI22_X1 port map( A1 => n1957, A2 => n2098, B1 => n757, B2 => n2092,
                           ZN => n1494);
   U447 : OAI22_X1 port map( A1 => n1958, A2 => n2098, B1 => n759, B2 => n2092,
                           ZN => n1493);
   U448 : OAI22_X1 port map( A1 => n1959, A2 => n2098, B1 => n761, B2 => n2092,
                           ZN => n1492);
   U449 : OAI22_X1 port map( A1 => n1960, A2 => n2098, B1 => n763, B2 => n2092,
                           ZN => n1491);
   U450 : OAI22_X1 port map( A1 => n1961, A2 => n2098, B1 => n765, B2 => n2092,
                           ZN => n1490);
   U451 : OAI22_X1 port map( A1 => n1962, A2 => n2098, B1 => n767, B2 => n2092,
                           ZN => n1489);
   U452 : OAI22_X1 port map( A1 => n1963, A2 => n2098, B1 => n769, B2 => n2092,
                           ZN => n1488);
   U453 : OAI22_X1 port map( A1 => n1964, A2 => n2098, B1 => n771, B2 => n2092,
                           ZN => n1487);
   U454 : OAI22_X1 port map( A1 => n1965, A2 => n2098, B1 => n773, B2 => n2092,
                           ZN => n1486);
   U455 : OAI22_X1 port map( A1 => n1966, A2 => n2098, B1 => n775, B2 => n2091,
                           ZN => n1485);
   U456 : OAI22_X1 port map( A1 => n1967, A2 => n2097, B1 => n777, B2 => n2091,
                           ZN => n1484);
   U457 : OAI22_X1 port map( A1 => n1968, A2 => n2097, B1 => n779, B2 => n2091,
                           ZN => n1483);
   U458 : OAI22_X1 port map( A1 => n1969, A2 => n2097, B1 => n781, B2 => n2091,
                           ZN => n1482);
   U459 : OAI22_X1 port map( A1 => n1970, A2 => n2097, B1 => n783, B2 => n2091,
                           ZN => n1481);
   U460 : OAI22_X1 port map( A1 => n1971, A2 => n2097, B1 => n785, B2 => n2091,
                           ZN => n1480);
   U461 : OAI22_X1 port map( A1 => n1972, A2 => n2097, B1 => n787, B2 => n2091,
                           ZN => n1479);
   U462 : OAI22_X1 port map( A1 => n1973, A2 => n2097, B1 => n789, B2 => n2091,
                           ZN => n1478);
   U463 : OAI22_X1 port map( A1 => n1974, A2 => n2097, B1 => n791, B2 => n2091,
                           ZN => n1477);
   U464 : OAI22_X1 port map( A1 => n1975, A2 => n2097, B1 => n793, B2 => n2091,
                           ZN => n1476);
   U465 : OAI22_X1 port map( A1 => n1976, A2 => n2097, B1 => n795, B2 => n2091,
                           ZN => n1475);
   U466 : OAI22_X1 port map( A1 => n1977, A2 => n2097, B1 => n797, B2 => n2091,
                           ZN => n1474);
   U467 : OAI22_X1 port map( A1 => n1978, A2 => n2097, B1 => n799, B2 => n2090,
                           ZN => n1473);
   U468 : OAI22_X1 port map( A1 => n1979, A2 => n2096, B1 => n801, B2 => n2090,
                           ZN => n1472);
   U469 : OAI22_X1 port map( A1 => n1980, A2 => n2096, B1 => n803, B2 => n2090,
                           ZN => n1471);
   U470 : OAI22_X1 port map( A1 => n1981, A2 => n2096, B1 => n805, B2 => n2090,
                           ZN => n1470);
   U471 : OAI22_X1 port map( A1 => n1982, A2 => n2096, B1 => n807, B2 => n2090,
                           ZN => n1469);
   U472 : OAI22_X1 port map( A1 => n1983, A2 => n2096, B1 => n809, B2 => n2090,
                           ZN => n1468);
   U473 : OAI22_X1 port map( A1 => n1984, A2 => n2096, B1 => n811, B2 => n2090,
                           ZN => n1467);
   U474 : OAI22_X1 port map( A1 => n1985, A2 => n2096, B1 => n813, B2 => n2090,
                           ZN => n1466);
   U475 : OAI22_X1 port map( A1 => n1986, A2 => n2096, B1 => n815, B2 => n2090,
                           ZN => n1465);
   U476 : OAI22_X1 port map( A1 => n1987, A2 => n2096, B1 => n817, B2 => n2090,
                           ZN => n1464);
   U477 : OAI22_X1 port map( A1 => n1988, A2 => n2096, B1 => n819, B2 => n2090,
                           ZN => n1463);
   U478 : OAI22_X1 port map( A1 => n1989, A2 => n2096, B1 => n821, B2 => n2090,
                           ZN => n1462);
   U479 : OAI22_X1 port map( A1 => n1990, A2 => n2096, B1 => n823, B2 => n2089,
                           ZN => n1461);
   U480 : OAI22_X1 port map( A1 => n1991, A2 => n2095, B1 => n825, B2 => n2089,
                           ZN => n1460);
   U481 : OAI22_X1 port map( A1 => n1992, A2 => n2095, B1 => n827, B2 => n2089,
                           ZN => n1459);
   U482 : OAI22_X1 port map( A1 => n1993, A2 => n2095, B1 => n829, B2 => n2089,
                           ZN => n1458);
   U483 : OAI22_X1 port map( A1 => n1994, A2 => n2095, B1 => n831, B2 => n2089,
                           ZN => n1457);
   U484 : OAI22_X1 port map( A1 => n1995, A2 => n2095, B1 => n833, B2 => n2089,
                           ZN => n1456);
   U485 : OAI22_X1 port map( A1 => n1996, A2 => n2095, B1 => n835, B2 => n2089,
                           ZN => n1455);
   U486 : OAI22_X1 port map( A1 => n1997, A2 => n2095, B1 => n837, B2 => n2089,
                           ZN => n1454);
   U487 : OAI22_X1 port map( A1 => n1998, A2 => n2095, B1 => n839, B2 => n2089,
                           ZN => n1453);
   U488 : OAI22_X1 port map( A1 => n1999, A2 => n2095, B1 => n841, B2 => n2089,
                           ZN => n1452);
   U489 : OAI22_X1 port map( A1 => n2000, A2 => n2095, B1 => n843, B2 => n2089,
                           ZN => n1451);
   U490 : OAI22_X1 port map( A1 => n2001, A2 => n2095, B1 => n845, B2 => n2089,
                           ZN => n1450);
   U491 : OAI22_X1 port map( A1 => n1204, A2 => n2095, B1 => n847, B2 => n2088,
                           ZN => n1449);
   U492 : OAI22_X1 port map( A1 => n1202, A2 => n2094, B1 => n849, B2 => n2088,
                           ZN => n1448);
   U493 : OAI22_X1 port map( A1 => n1200, A2 => n2094, B1 => n851, B2 => n2088,
                           ZN => n1447);
   U494 : OAI22_X1 port map( A1 => n2002, A2 => n2094, B1 => n853, B2 => n2088,
                           ZN => n1446);
   U495 : OAI22_X1 port map( A1 => n2003, A2 => n2094, B1 => n855, B2 => n2088,
                           ZN => n1445);
   U496 : OAI22_X1 port map( A1 => n2004, A2 => n2094, B1 => n857, B2 => n2088,
                           ZN => n1444);
   U497 : OAI22_X1 port map( A1 => n2005, A2 => n2094, B1 => n859, B2 => n2088,
                           ZN => n1443);
   U498 : OAI22_X1 port map( A1 => n2006, A2 => n2094, B1 => n861, B2 => n2088,
                           ZN => n1442);
   U499 : OAI22_X1 port map( A1 => n2007, A2 => n2094, B1 => n863, B2 => n2088,
                           ZN => n1441);
   U500 : OAI22_X1 port map( A1 => n2008, A2 => n2094, B1 => n865, B2 => n2088,
                           ZN => n1440);
   U501 : OAI22_X1 port map( A1 => n2009, A2 => n2094, B1 => n867, B2 => n2088,
                           ZN => n1439);
   U502 : OAI22_X1 port map( A1 => n415, A2 => n2094, B1 => n871, B2 => n2088, 
                           ZN => n1438);
   U503 : OAI22_X1 port map( A1 => n1817, A2 => n2087, B1 => n751, B2 => n2080,
                           ZN => n1433);
   U504 : OAI22_X1 port map( A1 => n1816, A2 => n2086, B1 => n753, B2 => n2080,
                           ZN => n1432);
   U505 : OAI22_X1 port map( A1 => n1815, A2 => n2086, B1 => n755, B2 => n2080,
                           ZN => n1431);
   U506 : OAI22_X1 port map( A1 => n1814, A2 => n2086, B1 => n757, B2 => n2080,
                           ZN => n1430);
   U507 : OAI22_X1 port map( A1 => n1813, A2 => n2086, B1 => n759, B2 => n2080,
                           ZN => n1429);
   U508 : OAI22_X1 port map( A1 => n1812, A2 => n2086, B1 => n761, B2 => n2080,
                           ZN => n1428);
   U509 : OAI22_X1 port map( A1 => n1811, A2 => n2086, B1 => n763, B2 => n2080,
                           ZN => n1427);
   U510 : OAI22_X1 port map( A1 => n1810, A2 => n2086, B1 => n765, B2 => n2080,
                           ZN => n1426);
   U511 : OAI22_X1 port map( A1 => n1809, A2 => n2086, B1 => n767, B2 => n2080,
                           ZN => n1425);
   U512 : OAI22_X1 port map( A1 => n1808, A2 => n2086, B1 => n769, B2 => n2080,
                           ZN => n1424);
   U513 : OAI22_X1 port map( A1 => n1807, A2 => n2086, B1 => n771, B2 => n2080,
                           ZN => n1423);
   U514 : OAI22_X1 port map( A1 => n1806, A2 => n2086, B1 => n773, B2 => n2080,
                           ZN => n1422);
   U515 : OAI22_X1 port map( A1 => n1805, A2 => n2086, B1 => n775, B2 => n2079,
                           ZN => n1421);
   U516 : OAI22_X1 port map( A1 => n1804, A2 => n2085, B1 => n777, B2 => n2079,
                           ZN => n1420);
   U517 : OAI22_X1 port map( A1 => n1803, A2 => n2085, B1 => n779, B2 => n2079,
                           ZN => n1419);
   U518 : OAI22_X1 port map( A1 => n1802, A2 => n2085, B1 => n781, B2 => n2079,
                           ZN => n1418);
   U519 : OAI22_X1 port map( A1 => n1801, A2 => n2085, B1 => n783, B2 => n2079,
                           ZN => n1417);
   U520 : OAI22_X1 port map( A1 => n1800, A2 => n2085, B1 => n785, B2 => n2079,
                           ZN => n1416);
   U521 : OAI22_X1 port map( A1 => n1799, A2 => n2085, B1 => n787, B2 => n2079,
                           ZN => n1415);
   U522 : OAI22_X1 port map( A1 => n1798, A2 => n2085, B1 => n789, B2 => n2079,
                           ZN => n1414);
   U523 : OAI22_X1 port map( A1 => n1797, A2 => n2085, B1 => n791, B2 => n2079,
                           ZN => n1413);
   U524 : OAI22_X1 port map( A1 => n1796, A2 => n2085, B1 => n793, B2 => n2079,
                           ZN => n1412);
   U525 : OAI22_X1 port map( A1 => n1795, A2 => n2085, B1 => n795, B2 => n2079,
                           ZN => n1411);
   U526 : OAI22_X1 port map( A1 => n1794, A2 => n2085, B1 => n797, B2 => n2079,
                           ZN => n1410);
   U527 : OAI22_X1 port map( A1 => n1793, A2 => n2085, B1 => n799, B2 => n2078,
                           ZN => n1409);
   U528 : OAI22_X1 port map( A1 => n2029, A2 => n2084, B1 => n801, B2 => n2078,
                           ZN => n1408);
   U529 : OAI22_X1 port map( A1 => n2030, A2 => n2084, B1 => n803, B2 => n2078,
                           ZN => n1407);
   U530 : OAI22_X1 port map( A1 => n2031, A2 => n2084, B1 => n805, B2 => n2078,
                           ZN => n1406);
   U531 : OAI22_X1 port map( A1 => n2032, A2 => n2084, B1 => n807, B2 => n2078,
                           ZN => n1405);
   U532 : OAI22_X1 port map( A1 => n2033, A2 => n2084, B1 => n809, B2 => n2078,
                           ZN => n1404);
   U533 : OAI22_X1 port map( A1 => n2034, A2 => n2084, B1 => n811, B2 => n2078,
                           ZN => n1403);
   U534 : OAI22_X1 port map( A1 => n2035, A2 => n2084, B1 => n813, B2 => n2078,
                           ZN => n1402);
   U535 : OAI22_X1 port map( A1 => n2036, A2 => n2084, B1 => n815, B2 => n2078,
                           ZN => n1401);
   U536 : OAI22_X1 port map( A1 => n2037, A2 => n2084, B1 => n817, B2 => n2078,
                           ZN => n1400);
   U537 : OAI22_X1 port map( A1 => n2038, A2 => n2084, B1 => n819, B2 => n2078,
                           ZN => n1399);
   U538 : OAI22_X1 port map( A1 => n2039, A2 => n2084, B1 => n821, B2 => n2078,
                           ZN => n1398);
   U539 : OAI22_X1 port map( A1 => n2040, A2 => n2084, B1 => n823, B2 => n2077,
                           ZN => n1397);
   U540 : OAI22_X1 port map( A1 => n2041, A2 => n2083, B1 => n825, B2 => n2077,
                           ZN => n1396);
   U541 : OAI22_X1 port map( A1 => n2042, A2 => n2083, B1 => n827, B2 => n2077,
                           ZN => n1395);
   U542 : OAI22_X1 port map( A1 => n2043, A2 => n2083, B1 => n829, B2 => n2077,
                           ZN => n1394);
   U543 : OAI22_X1 port map( A1 => n2044, A2 => n2083, B1 => n831, B2 => n2077,
                           ZN => n1393);
   U544 : OAI22_X1 port map( A1 => n2045, A2 => n2083, B1 => n833, B2 => n2077,
                           ZN => n1392);
   U545 : OAI22_X1 port map( A1 => n2046, A2 => n2083, B1 => n835, B2 => n2077,
                           ZN => n1391);
   U546 : OAI22_X1 port map( A1 => n2047, A2 => n2083, B1 => n837, B2 => n2077,
                           ZN => n1390);
   U547 : OAI22_X1 port map( A1 => n2048, A2 => n2083, B1 => n839, B2 => n2077,
                           ZN => n1389);
   U548 : OAI22_X1 port map( A1 => n2049, A2 => n2083, B1 => n841, B2 => n2077,
                           ZN => n1388);
   U549 : OAI22_X1 port map( A1 => n2050, A2 => n2083, B1 => n843, B2 => n2077,
                           ZN => n1387);
   U550 : OAI22_X1 port map( A1 => n2051, A2 => n2083, B1 => n845, B2 => n2077,
                           ZN => n1386);
   U551 : OAI22_X1 port map( A1 => n2052, A2 => n2083, B1 => n847, B2 => n2076,
                           ZN => n1385);
   U552 : OAI22_X1 port map( A1 => n2053, A2 => n2082, B1 => n849, B2 => n2076,
                           ZN => n1384);
   U553 : OAI22_X1 port map( A1 => n2054, A2 => n2082, B1 => n851, B2 => n2076,
                           ZN => n1383);
   U554 : OAI22_X1 port map( A1 => n2055, A2 => n2082, B1 => n853, B2 => n2076,
                           ZN => n1382);
   U555 : OAI22_X1 port map( A1 => n2056, A2 => n2082, B1 => n855, B2 => n2076,
                           ZN => n1381);
   U556 : OAI22_X1 port map( A1 => n2057, A2 => n2082, B1 => n857, B2 => n2076,
                           ZN => n1380);
   U557 : OAI22_X1 port map( A1 => n2058, A2 => n2082, B1 => n859, B2 => n2076,
                           ZN => n1379);
   U558 : OAI22_X1 port map( A1 => n2059, A2 => n2082, B1 => n861, B2 => n2076,
                           ZN => n1378);
   U559 : OAI22_X1 port map( A1 => n2060, A2 => n2082, B1 => n863, B2 => n2076,
                           ZN => n1377);
   U560 : OAI22_X1 port map( A1 => n2061, A2 => n2082, B1 => n865, B2 => n2076,
                           ZN => n1376);
   U561 : OAI22_X1 port map( A1 => n2062, A2 => n2082, B1 => n867, B2 => n2076,
                           ZN => n1375);
   U562 : OAI22_X1 port map( A1 => n2063, A2 => n2082, B1 => n871, B2 => n2076,
                           ZN => n1374);
   U563 : OAI22_X1 port map( A1 => n2014, A2 => n2075, B1 => n751, B2 => n2068,
                           ZN => n1369);
   U564 : OAI22_X1 port map( A1 => n2015, A2 => n2074, B1 => n753, B2 => n2068,
                           ZN => n1368);
   U565 : OAI22_X1 port map( A1 => n2016, A2 => n2074, B1 => n755, B2 => n2068,
                           ZN => n1367);
   U566 : OAI22_X1 port map( A1 => n2017, A2 => n2074, B1 => n757, B2 => n2068,
                           ZN => n1366);
   U567 : OAI22_X1 port map( A1 => n2018, A2 => n2074, B1 => n759, B2 => n2068,
                           ZN => n1365);
   U568 : OAI22_X1 port map( A1 => n2019, A2 => n2074, B1 => n761, B2 => n2068,
                           ZN => n1364);
   U569 : OAI22_X1 port map( A1 => n2020, A2 => n2074, B1 => n763, B2 => n2068,
                           ZN => n1363);
   U570 : OAI22_X1 port map( A1 => n2021, A2 => n2074, B1 => n765, B2 => n2068,
                           ZN => n1362);
   U571 : OAI22_X1 port map( A1 => n2022, A2 => n2074, B1 => n767, B2 => n2068,
                           ZN => n1361);
   U572 : OAI22_X1 port map( A1 => n2023, A2 => n2074, B1 => n769, B2 => n2068,
                           ZN => n1360);
   U573 : OAI22_X1 port map( A1 => n2024, A2 => n2074, B1 => n771, B2 => n2068,
                           ZN => n1359);
   U574 : OAI22_X1 port map( A1 => n2025, A2 => n2074, B1 => n773, B2 => n2068,
                           ZN => n1358);
   U575 : OAI22_X1 port map( A1 => n2026, A2 => n2074, B1 => n775, B2 => n2067,
                           ZN => n1357);
   U576 : OAI22_X1 port map( A1 => n2027, A2 => n2073, B1 => n777, B2 => n2067,
                           ZN => n1356);
   U577 : OAI22_X1 port map( A1 => n2028, A2 => n2073, B1 => n779, B2 => n2067,
                           ZN => n1355);
   U578 : OAI22_X1 port map( A1 => n1738, A2 => n2073, B1 => n781, B2 => n2067,
                           ZN => n1354);
   U579 : OAI22_X1 port map( A1 => n1737, A2 => n2073, B1 => n783, B2 => n2067,
                           ZN => n1353);
   U580 : OAI22_X1 port map( A1 => n1736, A2 => n2073, B1 => n785, B2 => n2067,
                           ZN => n1352);
   U581 : OAI22_X1 port map( A1 => n1735, A2 => n2073, B1 => n787, B2 => n2067,
                           ZN => n1351);
   U582 : OAI22_X1 port map( A1 => n1734, A2 => n2073, B1 => n789, B2 => n2067,
                           ZN => n1350);
   U583 : OAI22_X1 port map( A1 => n1733, A2 => n2073, B1 => n791, B2 => n2067,
                           ZN => n1349);
   U584 : OAI22_X1 port map( A1 => n1732, A2 => n2073, B1 => n793, B2 => n2067,
                           ZN => n1348);
   U585 : OAI22_X1 port map( A1 => n1731, A2 => n2073, B1 => n795, B2 => n2067,
                           ZN => n1347);
   U586 : OAI22_X1 port map( A1 => n1730, A2 => n2073, B1 => n797, B2 => n2067,
                           ZN => n1346);
   U587 : OAI22_X1 port map( A1 => n1729, A2 => n2073, B1 => n799, B2 => n2066,
                           ZN => n1345);
   U588 : OAI22_X1 port map( A1 => n1728, A2 => n2072, B1 => n801, B2 => n2066,
                           ZN => n1344);
   U589 : OAI22_X1 port map( A1 => n1727, A2 => n2072, B1 => n803, B2 => n2066,
                           ZN => n1343);
   U590 : OAI22_X1 port map( A1 => n1726, A2 => n2072, B1 => n805, B2 => n2066,
                           ZN => n1342);
   U591 : OAI22_X1 port map( A1 => n1725, A2 => n2072, B1 => n807, B2 => n2066,
                           ZN => n1341);
   U592 : OAI22_X1 port map( A1 => n1724, A2 => n2072, B1 => n809, B2 => n2066,
                           ZN => n1340);
   U593 : OAI22_X1 port map( A1 => n1723, A2 => n2072, B1 => n811, B2 => n2066,
                           ZN => n1339);
   U594 : OAI22_X1 port map( A1 => n1722, A2 => n2072, B1 => n813, B2 => n2066,
                           ZN => n1338);
   U595 : OAI22_X1 port map( A1 => n1721, A2 => n2072, B1 => n815, B2 => n2066,
                           ZN => n1337);
   U596 : OAI22_X1 port map( A1 => n1720, A2 => n2072, B1 => n817, B2 => n2066,
                           ZN => n1336);
   U597 : OAI22_X1 port map( A1 => n1719, A2 => n2072, B1 => n819, B2 => n2066,
                           ZN => n1335);
   U598 : OAI22_X1 port map( A1 => n1718, A2 => n2072, B1 => n821, B2 => n2066,
                           ZN => n1334);
   U599 : OAI22_X1 port map( A1 => n1717, A2 => n2072, B1 => n823, B2 => n2065,
                           ZN => n1333);
   U600 : OAI22_X1 port map( A1 => n1716, A2 => n2071, B1 => n825, B2 => n2065,
                           ZN => n1332);
   U601 : OAI22_X1 port map( A1 => n1715, A2 => n2071, B1 => n827, B2 => n2065,
                           ZN => n1331);
   U602 : OAI22_X1 port map( A1 => n1714, A2 => n2071, B1 => n829, B2 => n2065,
                           ZN => n1330);
   U603 : OAI22_X1 port map( A1 => n1713, A2 => n2071, B1 => n831, B2 => n2065,
                           ZN => n1329);
   U604 : OAI22_X1 port map( A1 => n1712, A2 => n2071, B1 => n833, B2 => n2065,
                           ZN => n1328);
   U605 : OAI22_X1 port map( A1 => n1711, A2 => n2071, B1 => n835, B2 => n2065,
                           ZN => n1327);
   U606 : OAI22_X1 port map( A1 => n1710, A2 => n2071, B1 => n837, B2 => n2065,
                           ZN => n1326);
   U607 : OAI22_X1 port map( A1 => n1709, A2 => n2071, B1 => n839, B2 => n2065,
                           ZN => n1325);
   U608 : OAI22_X1 port map( A1 => n1708, A2 => n2071, B1 => n841, B2 => n2065,
                           ZN => n1324);
   U609 : OAI22_X1 port map( A1 => n1707, A2 => n2071, B1 => n843, B2 => n2065,
                           ZN => n1323);
   U610 : OAI22_X1 port map( A1 => n1706, A2 => n2071, B1 => n845, B2 => n2065,
                           ZN => n1322);
   U611 : OAI22_X1 port map( A1 => n1705, A2 => n2071, B1 => n847, B2 => n2064,
                           ZN => n1321);
   U612 : OAI22_X1 port map( A1 => n1704, A2 => n2070, B1 => n849, B2 => n2064,
                           ZN => n1320);
   U613 : OAI22_X1 port map( A1 => n1703, A2 => n2070, B1 => n851, B2 => n2064,
                           ZN => n1319);
   U614 : OAI22_X1 port map( A1 => n1702, A2 => n2070, B1 => n853, B2 => n2064,
                           ZN => n1318);
   U615 : OAI22_X1 port map( A1 => n1701, A2 => n2070, B1 => n855, B2 => n2064,
                           ZN => n1317);
   U616 : OAI22_X1 port map( A1 => n1700, A2 => n2070, B1 => n857, B2 => n2064,
                           ZN => n1316);
   U617 : OAI22_X1 port map( A1 => n1699, A2 => n2070, B1 => n859, B2 => n2064,
                           ZN => n1315);
   U618 : OAI22_X1 port map( A1 => n1698, A2 => n2070, B1 => n861, B2 => n2064,
                           ZN => n1314);
   U619 : OAI22_X1 port map( A1 => n1697, A2 => n2070, B1 => n863, B2 => n2064,
                           ZN => n1313);
   U620 : OAI22_X1 port map( A1 => n1696, A2 => n2070, B1 => n865, B2 => n2064,
                           ZN => n1312);
   U621 : OAI22_X1 port map( A1 => n1695, A2 => n2070, B1 => n867, B2 => n2064,
                           ZN => n1311);
   U622 : OAI22_X1 port map( A1 => n1694, A2 => n2070, B1 => n871, B2 => n2064,
                           ZN => n1310);
   U623 : INV_X1 port map( A => DATAIN(0), ZN => n743);
   U624 : INV_X1 port map( A => DATAIN(1), ZN => n745);
   U625 : INV_X1 port map( A => DATAIN(2), ZN => n747);
   U626 : INV_X1 port map( A => DATAIN(3), ZN => n749);
   U627 : INV_X1 port map( A => DATAIN(4), ZN => n751);
   U628 : INV_X1 port map( A => DATAIN(5), ZN => n753);
   U629 : INV_X1 port map( A => DATAIN(6), ZN => n755);
   U630 : INV_X1 port map( A => DATAIN(7), ZN => n757);
   U631 : INV_X1 port map( A => DATAIN(8), ZN => n759);
   U632 : INV_X1 port map( A => DATAIN(9), ZN => n761);
   U633 : INV_X1 port map( A => DATAIN(10), ZN => n763);
   U634 : INV_X1 port map( A => DATAIN(11), ZN => n765);
   U635 : INV_X1 port map( A => DATAIN(12), ZN => n767);
   U636 : INV_X1 port map( A => DATAIN(13), ZN => n769);
   U637 : INV_X1 port map( A => DATAIN(14), ZN => n771);
   U638 : INV_X1 port map( A => DATAIN(15), ZN => n773);
   U639 : INV_X1 port map( A => DATAIN(16), ZN => n775);
   U640 : INV_X1 port map( A => DATAIN(17), ZN => n777);
   U641 : INV_X1 port map( A => DATAIN(18), ZN => n779);
   U642 : INV_X1 port map( A => DATAIN(19), ZN => n781);
   U643 : INV_X1 port map( A => DATAIN(20), ZN => n783);
   U644 : INV_X1 port map( A => DATAIN(21), ZN => n785);
   U645 : INV_X1 port map( A => DATAIN(22), ZN => n787);
   U646 : INV_X1 port map( A => DATAIN(23), ZN => n789);
   U647 : INV_X1 port map( A => DATAIN(24), ZN => n791);
   U648 : INV_X1 port map( A => DATAIN(25), ZN => n793);
   U649 : INV_X1 port map( A => DATAIN(26), ZN => n795);
   U650 : INV_X1 port map( A => DATAIN(27), ZN => n797);
   U651 : INV_X1 port map( A => DATAIN(28), ZN => n799);
   U652 : INV_X1 port map( A => DATAIN(29), ZN => n801);
   U653 : INV_X1 port map( A => DATAIN(30), ZN => n803);
   U654 : INV_X1 port map( A => DATAIN(31), ZN => n805);
   U655 : INV_X1 port map( A => DATAIN(32), ZN => n807);
   U656 : INV_X1 port map( A => DATAIN(33), ZN => n809);
   U657 : INV_X1 port map( A => DATAIN(34), ZN => n811);
   U658 : INV_X1 port map( A => DATAIN(35), ZN => n813);
   U659 : INV_X1 port map( A => DATAIN(36), ZN => n815);
   U660 : INV_X1 port map( A => DATAIN(37), ZN => n817);
   U661 : INV_X1 port map( A => DATAIN(38), ZN => n819);
   U662 : INV_X1 port map( A => DATAIN(39), ZN => n821);
   U663 : INV_X1 port map( A => DATAIN(40), ZN => n823);
   U664 : INV_X1 port map( A => DATAIN(41), ZN => n825);
   U665 : INV_X1 port map( A => DATAIN(42), ZN => n827);
   U666 : INV_X1 port map( A => DATAIN(43), ZN => n829);
   U667 : INV_X1 port map( A => DATAIN(44), ZN => n831);
   U668 : INV_X1 port map( A => DATAIN(45), ZN => n833);
   U669 : INV_X1 port map( A => DATAIN(46), ZN => n835);
   U670 : INV_X1 port map( A => DATAIN(47), ZN => n837);
   U671 : INV_X1 port map( A => DATAIN(48), ZN => n839);
   U672 : INV_X1 port map( A => DATAIN(49), ZN => n841);
   U673 : INV_X1 port map( A => DATAIN(50), ZN => n843);
   U674 : INV_X1 port map( A => DATAIN(51), ZN => n845);
   U675 : INV_X1 port map( A => DATAIN(52), ZN => n847);
   U676 : INV_X1 port map( A => DATAIN(53), ZN => n849);
   U677 : INV_X1 port map( A => DATAIN(54), ZN => n851);
   U678 : INV_X1 port map( A => DATAIN(55), ZN => n853);
   U679 : INV_X1 port map( A => DATAIN(56), ZN => n855);
   U680 : INV_X1 port map( A => DATAIN(57), ZN => n857);
   U681 : INV_X1 port map( A => DATAIN(58), ZN => n859);
   U682 : INV_X1 port map( A => DATAIN(59), ZN => n861);
   U683 : INV_X1 port map( A => DATAIN(60), ZN => n863);
   U684 : INV_X1 port map( A => DATAIN(61), ZN => n865);
   U685 : INV_X1 port map( A => DATAIN(62), ZN => n867);
   U686 : INV_X1 port map( A => DATAIN(63), ZN => n871);
   U687 : CLKBUF_X1 port map( A => n979, Z => n2069);
   U688 : CLKBUF_X1 port map( A => n978, Z => n2075);
   U689 : CLKBUF_X1 port map( A => n939, Z => n2081);
   U690 : CLKBUF_X1 port map( A => n938, Z => n2087);
   U691 : CLKBUF_X1 port map( A => n876, Z => n2093);
   U692 : CLKBUF_X1 port map( A => n875, Z => n2099);
   U693 : CLKBUF_X1 port map( A => n742, Z => n2105);
   U694 : CLKBUF_X1 port map( A => n741, Z => n2111);
   U695 : CLKBUF_X1 port map( A => n740, Z => n2117);
   U696 : CLKBUF_X1 port map( A => n739, Z => n2123);
   U697 : CLKBUF_X1 port map( A => n738, Z => n2129);
   U698 : CLKBUF_X1 port map( A => n736, Z => n2135);
   U699 : CLKBUF_X1 port map( A => n735, Z => n2141);
   U700 : CLKBUF_X1 port map( A => n527, Z => n2147);
   U701 : CLKBUF_X1 port map( A => n525, Z => n2158);
   U702 : CLKBUF_X1 port map( A => n523, Z => n2164);
   U703 : CLKBUF_X1 port map( A => n521, Z => n2170);
   U704 : INV_X1 port map( A => ADD_RD2(0), ZN => n2171);
   U705 : INV_X1 port map( A => ADD_RD2(1), ZN => n2172);
   U706 : INV_X1 port map( A => ADD_RD1(0), ZN => n2173);
   U707 : INV_X1 port map( A => ADD_RD1(1), ZN => n2174);
   U708 : INV_X1 port map( A => ADD_WR(0), ZN => n2175);
   U709 : INV_X1 port map( A => ADD_WR(1), ZN => n2176);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4.all;

entity register_file_reg_size64_file_size4_5 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_reg_size64_file_size4_5;

architecture SYN_BEHAVIORAL of register_file_reg_size64_file_size4_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n415, n1200, n1202, n1204, n1310, n1311, n1312, n1313, n1314, n1315
      , n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n871, n872, 
      n873, n875, n876, n936, n938, n939, n975, n978, n979, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176 : std_logic
      ;

begin
   
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => n174,
                           QN => n2028);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => n175,
                           QN => n2027);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => n176,
                           QN => n2026);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => n177,
                           QN => n2025);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => n178,
                           QN => n2024);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => n179,
                           QN => n2023);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => n180,
                           QN => n2022);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => n181,
                           QN => n2021);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => n182,
                           QN => n2020);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => n183, 
                           QN => n2019);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => n184, 
                           QN => n2018);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => n185, 
                           QN => n2017);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => n186, 
                           QN => n2016);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => n187, 
                           QN => n2015);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => n188, 
                           QN => n2014);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => n189, 
                           QN => n2013);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => n190, 
                           QN => n2012);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => n191, 
                           QN => n2011);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => n192, 
                           QN => n2010);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => n65, 
                           QN => n2063);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => n66, 
                           QN => n2062);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n67, 
                           QN => n2061);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => n68, 
                           QN => n2060);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => n69, 
                           QN => n2059);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => n70, 
                           QN => n2058);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => n71, 
                           QN => n2057);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => n72, 
                           QN => n2056);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => n73, 
                           QN => n2055);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => n74, 
                           QN => n2054);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => n75, 
                           QN => n2053);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => n76, 
                           QN => n2052);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => n77, 
                           QN => n2051);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => n78, 
                           QN => n2050);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => n79, 
                           QN => n2049);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => n80, 
                           QN => n2048);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => n81, 
                           QN => n2047);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => n82, 
                           QN => n2046);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => n83, 
                           QN => n2045);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => n84, 
                           QN => n2044);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => n85, 
                           QN => n2043);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => n86, 
                           QN => n2042);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => n87, 
                           QN => n2041);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => n88, 
                           QN => n2040);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => n89, 
                           QN => n2039);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => n90, 
                           QN => n2038);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => n91, 
                           QN => n2037);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => n92, 
                           QN => n2036);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => n93, 
                           QN => n2035);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => n94, 
                           QN => n2034);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => n95, 
                           QN => n2033);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => n96, 
                           QN => n2032);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => n97, 
                           QN => n2031);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => n98, 
                           QN => n2030);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => n99, 
                           QN => n2029);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => n2, 
                           QN => n2009);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => n3, 
                           QN => n2008);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => n4, 
                           QN => n2007);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => n5, 
                           QN => n2006);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => n6, 
                           QN => n2005);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => n7, 
                           QN => n2004);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => n8, 
                           QN => n2003);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => n9, 
                           QN => n2002);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => n13, 
                           QN => n2001);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => n14, 
                           QN => n2000);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => n15, 
                           QN => n1999);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => n16, 
                           QN => n1998);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => n17, 
                           QN => n1997);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => n18, 
                           QN => n1996);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => n19, 
                           QN => n1995);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => n20, 
                           QN => n1994);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => n21, 
                           QN => n1993);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => n22, 
                           QN => n1992);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => n23, 
                           QN => n1991);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => n24, 
                           QN => n1990);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => n25, 
                           QN => n1989);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => n26, 
                           QN => n1988);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n27, 
                           QN => n1987);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => n28, 
                           QN => n1986);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n29, 
                           QN => n1985);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => n30, 
                           QN => n1984);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n31, 
                           QN => n1983);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => n32, 
                           QN => n1982);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n33, 
                           QN => n1981);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => n34, 
                           QN => n1980);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n35, 
                           QN => n1979);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => n36, 
                           QN => n1978);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => n37, 
                           QN => n1977);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => n38, 
                           QN => n1976);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => n39, 
                           QN => n1975);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => n40, 
                           QN => n1974);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => n41, 
                           QN => n1973);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => n42, 
                           QN => n1972);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => n43, 
                           QN => n1971);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => n44, 
                           QN => n1970);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => n45, 
                           QN => n1969);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => n46, 
                           QN => n1968);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => n47, 
                           QN => n1967);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => n48, 
                           QN => n1966);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => n49, 
                           QN => n1965);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => n50, 
                           QN => n1964);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => n51, 
                           QN => n1963);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => n52, 
                           QN => n1962);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => n53, 
                           QN => n1961);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => n54, 
                           QN => n1960);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n55, 
                           QN => n1959);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => n56, 
                           QN => n1958);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n57, 
                           QN => n1957);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => n58, 
                           QN => n1956);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n59, 
                           QN => n1955);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => n60, 
                           QN => n1954);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n61, 
                           QN => n1953);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => n62, 
                           QN => n1952);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n63, 
                           QN => n1951);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => n64, 
                           QN => n1950);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n999,
                           QN => n728);
   OUT2_reg_63_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => OUT2(63), QN
                           => n1822);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n1000
                           , QN => n725);
   OUT2_reg_62_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => OUT2(62), QN
                           => n1823);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n1001
                           , QN => n722);
   OUT2_reg_61_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => OUT2(61), QN
                           => n1824);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n1002
                           , QN => n719);
   OUT2_reg_60_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => OUT2(60), QN
                           => n1825);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n1003
                           , QN => n716);
   OUT2_reg_59_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => OUT2(59), QN
                           => n1826);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n1004
                           , QN => n713);
   OUT2_reg_58_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => OUT2(58), QN
                           => n1827);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n1005
                           , QN => n710);
   OUT2_reg_57_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => OUT2(57), QN
                           => n1828);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n1006
                           , QN => n707);
   OUT2_reg_56_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => OUT2(56), QN
                           => n1829);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n1007
                           , QN => n704);
   OUT2_reg_55_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => OUT2(55), QN
                           => n1830);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n1008
                           , QN => n700);
   OUT2_reg_54_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => OUT2(54), QN
                           => n1831);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n1009
                           , QN => n696);
   OUT2_reg_53_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => OUT2(53), QN
                           => n1832);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n1010
                           , QN => n692);
   OUT2_reg_52_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => OUT2(52), QN
                           => n1833);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n1011
                           , QN => n689);
   OUT2_reg_51_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => OUT2(51), QN
                           => n1834);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n1012
                           , QN => n686);
   OUT2_reg_50_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => OUT2(50), QN
                           => n1835);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n1013
                           , QN => n683);
   OUT2_reg_49_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => OUT2(49), QN
                           => n1836);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n1014
                           , QN => n680);
   OUT2_reg_48_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => OUT2(48), QN
                           => n1837);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n1015
                           , QN => n677);
   OUT2_reg_47_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => OUT2(47), QN
                           => n1838);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n1016
                           , QN => n674);
   OUT2_reg_46_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => OUT2(46), QN
                           => n1839);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n1017
                           , QN => n671);
   OUT2_reg_45_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => OUT2(45), QN
                           => n1840);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n1018
                           , QN => n668);
   OUT2_reg_44_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => OUT2(44), QN
                           => n1841);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n1019
                           , QN => n665);
   OUT2_reg_43_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => OUT2(43), QN
                           => n1842);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n1020
                           , QN => n662);
   OUT2_reg_42_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => OUT2(42), QN
                           => n1843);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n1021
                           , QN => n659);
   OUT2_reg_41_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => OUT2(41), QN
                           => n1844);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n1022
                           , QN => n656);
   OUT2_reg_40_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => OUT2(40), QN
                           => n1845);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n1023
                           , QN => n653);
   OUT2_reg_39_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => OUT2(39), QN
                           => n1846);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n1024
                           , QN => n650);
   OUT2_reg_38_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => OUT2(38), QN
                           => n1847);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n1025
                           , QN => n647);
   OUT2_reg_37_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => OUT2(37), QN
                           => n1848);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n1026
                           , QN => n644);
   OUT2_reg_36_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => OUT2(36), QN
                           => n1849);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n1027
                           , QN => n641);
   OUT2_reg_35_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => OUT2(35), QN
                           => n1850);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n1028
                           , QN => n638);
   OUT2_reg_34_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => OUT2(34), QN
                           => n1851);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n1029
                           , QN => n635);
   OUT2_reg_33_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => OUT2(33), QN
                           => n1852);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n1030
                           , QN => n632);
   OUT2_reg_32_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => OUT2(32), QN
                           => n1853);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n1031
                           , QN => n629);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => OUT2(31), QN
                           => n1854);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n1032
                           , QN => n626);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => OUT2(30), QN
                           => n1855);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n1033
                           , QN => n623);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => OUT2(29), QN
                           => n1856);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n1034
                           , QN => n619);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => OUT2(28), QN
                           => n1857);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n1035
                           , QN => n615);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => OUT2(27), QN
                           => n1858);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n1036
                           , QN => n611);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => OUT2(26), QN
                           => n1859);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n1037
                           , QN => n607);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => OUT2(25), QN
                           => n1860);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n1038
                           , QN => n603);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => OUT2(24), QN
                           => n1861);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n1039
                           , QN => n599);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => OUT2(23), QN
                           => n1862);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n1040
                           , QN => n595);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => OUT2(22), QN
                           => n1863);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n1041
                           , QN => n591);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => OUT2(21), QN
                           => n1864);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n1042
                           , QN => n587);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => OUT2(20), QN
                           => n1865);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n1043
                           , QN => n583);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => OUT2(19), QN
                           => n1866);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n1044
                           , QN => n580);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => OUT2(18), QN
                           => n1867);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n1045
                           , QN => n577);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => OUT2(17), QN
                           => n1868);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n1046
                           , QN => n574);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => OUT2(16), QN
                           => n1869);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n1047
                           , QN => n571);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => OUT2(15), QN
                           => n1870);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n1048
                           , QN => n568);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => OUT2(14), QN
                           => n1871);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n1049
                           , QN => n565);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => OUT2(13), QN
                           => n1872);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n1050
                           , QN => n562);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => OUT2(12), QN
                           => n1873);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n1051
                           , QN => n559);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => OUT2(11), QN
                           => n1874);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n1052
                           , QN => n556);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => OUT2(10), QN
                           => n1875);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n1053,
                           QN => n553);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => OUT2(9), QN 
                           => n1876);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => n1054,
                           QN => n550);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => OUT2(8), QN 
                           => n1877);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => n1055,
                           QN => n547);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => OUT2(7), QN 
                           => n1878);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => n1056,
                           QN => n544);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => OUT2(6), QN 
                           => n1879);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => n1057,
                           QN => n541);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => OUT2(5), QN 
                           => n1880);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => n1058,
                           QN => n538);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => OUT2(4), QN 
                           => n1881);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => n1059,
                           QN => n535);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => OUT2(3), QN 
                           => n1882);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n1060,
                           QN => n532);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => OUT2(2), QN 
                           => n1883);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n1061,
                           QN => n529);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => OUT2(1), QN 
                           => n1884);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n1062,
                           QN => n522);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => OUT2(0), QN 
                           => n1885);
   OUT1_reg_63_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => OUT1(63), QN
                           => n1886);
   OUT1_reg_62_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => OUT1(62), QN
                           => n1887);
   OUT1_reg_61_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => OUT1(61), QN
                           => n1888);
   OUT1_reg_60_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => OUT1(60), QN
                           => n1889);
   OUT1_reg_59_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => OUT1(59), QN
                           => n1890);
   OUT1_reg_58_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => OUT1(58), QN
                           => n1891);
   OUT1_reg_57_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => OUT1(57), QN
                           => n1892);
   OUT1_reg_56_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => OUT1(56), QN
                           => n1893);
   OUT1_reg_55_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => OUT1(55), QN
                           => n1894);
   OUT1_reg_54_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => OUT1(54), QN
                           => n1895);
   OUT1_reg_53_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => OUT1(53), QN
                           => n1896);
   OUT1_reg_52_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => OUT1(52), QN
                           => n1897);
   OUT1_reg_51_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => OUT1(51), QN
                           => n1898);
   OUT1_reg_50_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => OUT1(50), QN
                           => n1899);
   OUT1_reg_49_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => OUT1(49), QN
                           => n1900);
   OUT1_reg_48_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => OUT1(48), QN
                           => n1901);
   OUT1_reg_47_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => OUT1(47), QN
                           => n1902);
   OUT1_reg_46_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => OUT1(46), QN
                           => n1903);
   OUT1_reg_45_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => OUT1(45), QN
                           => n1904);
   OUT1_reg_44_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => OUT1(44), QN
                           => n1905);
   OUT1_reg_43_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => OUT1(43), QN
                           => n1906);
   OUT1_reg_42_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => OUT1(42), QN
                           => n1907);
   OUT1_reg_41_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => OUT1(41), QN
                           => n1908);
   OUT1_reg_40_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => OUT1(40), QN
                           => n1909);
   OUT1_reg_39_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => OUT1(39), QN
                           => n1910);
   OUT1_reg_38_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => OUT1(38), QN
                           => n1911);
   OUT1_reg_37_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => OUT1(37), QN
                           => n1912);
   OUT1_reg_36_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => OUT1(36), QN
                           => n1913);
   OUT1_reg_35_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => OUT1(35), QN
                           => n1914);
   OUT1_reg_34_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => OUT1(34), QN
                           => n1915);
   OUT1_reg_33_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => OUT1(33), QN
                           => n1916);
   OUT1_reg_32_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => OUT1(32), QN
                           => n1917);
   OUT1_reg_31_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => OUT1(31), QN
                           => n1918);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => OUT1(30), QN
                           => n1919);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => OUT1(29), QN
                           => n1920);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => OUT1(28), QN
                           => n1921);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => OUT1(27), QN
                           => n1922);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => OUT1(26), QN
                           => n1923);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => OUT1(25), QN
                           => n1924);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => OUT1(24), QN
                           => n1925);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => OUT1(23), QN
                           => n1926);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => OUT1(22), QN
                           => n1927);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => OUT1(21), QN
                           => n1928);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => OUT1(20), QN
                           => n1929);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => OUT1(19), QN
                           => n1930);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => OUT1(18), QN
                           => n1931);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => OUT1(17), QN
                           => n1932);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => OUT1(16), QN
                           => n1933);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => OUT1(15), QN
                           => n1934);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => OUT1(14), QN
                           => n1935);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => OUT1(13), QN
                           => n1936);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => OUT1(12), QN
                           => n1937);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => OUT1(11), QN
                           => n1938);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => OUT1(10), QN
                           => n1939);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => OUT1(9), QN 
                           => n1940);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => OUT1(8), QN 
                           => n1941);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => OUT1(7), QN 
                           => n1942);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => OUT1(6), QN 
                           => n1943);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => OUT1(5), QN 
                           => n1944);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => OUT1(4), QN 
                           => n1945);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => OUT1(3), QN 
                           => n1946);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => OUT1(2), QN 
                           => n1947);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => OUT1(1), QN 
                           => n1948);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => OUT1(0), QN 
                           => n1949);
   U859 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n2164, A3 => ADD_RD1(1), 
                           ZN => n521);
   U860 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n2135, A3 => ADD_RD2(1), 
                           ZN => n735);
   U861 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n873, A3 => ADD_WR(1), ZN 
                           => n872);
   U862 : NAND3_X1 port map( A1 => n873, A2 => n2175, A3 => ADD_WR(1), ZN => 
                           n936);
   U863 : NAND3_X1 port map( A1 => n873, A2 => n2176, A3 => ADD_WR(0), ZN => 
                           n975);
   U864 : NAND3_X1 port map( A1 => n2175, A2 => n2176, A3 => n873, ZN => n998);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => n537, 
                           QN => n1818);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => n534, 
                           QN => n1819);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => n531, 
                           QN => n1820);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => n528, 
                           QN => n1821);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => n730,
                           QN => n415);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => n702,
                           QN => n1200);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => n698,
                           QN => n1202);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => n694,
                           QN => n1204);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => n622,
                           QN => n1793);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => n618,
                           QN => n1794);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => n614,
                           QN => n1795);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => n610,
                           QN => n1796);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => n606,
                           QN => n1797);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => n602,
                           QN => n1798);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => n598,
                           QN => n1799);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => n594,
                           QN => n1800);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => n590,
                           QN => n1801);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => n586,
                           QN => n1802);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => n582,
                           QN => n1803);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => n579,
                           QN => n1804);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => n576,
                           QN => n1805);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => n573,
                           QN => n1806);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => n570,
                           QN => n1807);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => n567,
                           QN => n1808);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => n564,
                           QN => n1809);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => n561,
                           QN => n1810);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => n558,
                           QN => n1811);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => n555, 
                           QN => n1812);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => n552, 
                           QN => n1813);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => n549, 
                           QN => n1814);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => n546, 
                           QN => n1815);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => n543, 
                           QN => n1816);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => n540, 
                           QN => n1817);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => n731,
                           QN => n1694);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => n727,
                           QN => n1695);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => n724,
                           QN => n1696);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => n721,
                           QN => n1697);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => n718,
                           QN => n1698);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => n715,
                           QN => n1699);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => n712,
                           QN => n1700);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => n709,
                           QN => n1701);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => n706,
                           QN => n1702);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => n703,
                           QN => n1703);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => n699,
                           QN => n1704);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => n695,
                           QN => n1705);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => n691,
                           QN => n1706);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => n688,
                           QN => n1707);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => n685,
                           QN => n1708);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => n682,
                           QN => n1709);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => n679,
                           QN => n1710);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => n676,
                           QN => n1711);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => n673,
                           QN => n1712);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => n670,
                           QN => n1713);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => n667,
                           QN => n1714);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => n664,
                           QN => n1715);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => n661,
                           QN => n1716);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => n658,
                           QN => n1717);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => n655,
                           QN => n1718);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => n652,
                           QN => n1719);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => n649,
                           QN => n1720);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => n646,
                           QN => n1721);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => n643,
                           QN => n1722);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => n640,
                           QN => n1723);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => n637,
                           QN => n1724);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => n634,
                           QN => n1725);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => n631,
                           QN => n1726);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => n628,
                           QN => n1727);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n625,
                           QN => n1728);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => n621,
                           QN => n1729);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => n617,
                           QN => n1730);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => n613,
                           QN => n1731);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => n609,
                           QN => n1732);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => n605,
                           QN => n1733);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => n601,
                           QN => n1734);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => n597,
                           QN => n1735);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => n593,
                           QN => n1736);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => n589,
                           QN => n1737);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => n585,
                           QN => n1738);
   U3 : BUF_X1 port map( A => n521, Z => n2167);
   U4 : BUF_X1 port map( A => n521, Z => n2166);
   U5 : BUF_X1 port map( A => n521, Z => n2165);
   U6 : BUF_X1 port map( A => n735, Z => n2139);
   U7 : BUF_X1 port map( A => n735, Z => n2138);
   U8 : BUF_X1 port map( A => n735, Z => n2137);
   U9 : BUF_X1 port map( A => n735, Z => n2136);
   U10 : BUF_X1 port map( A => n521, Z => n2169);
   U11 : BUF_X1 port map( A => n521, Z => n2168);
   U12 : BUF_X1 port map( A => n735, Z => n2140);
   U13 : BUF_X1 port map( A => n526, Z => n2151);
   U14 : BUF_X1 port map( A => n526, Z => n2152);
   U15 : BUF_X1 port map( A => n527, Z => n2144);
   U16 : BUF_X1 port map( A => n527, Z => n2146);
   U17 : BUF_X1 port map( A => n527, Z => n2145);
   U18 : BUF_X1 port map( A => n523, Z => n2159);
   U19 : BUF_X1 port map( A => n523, Z => n2160);
   U20 : BUF_X1 port map( A => n523, Z => n2161);
   U21 : BUF_X1 port map( A => n523, Z => n2162);
   U22 : BUF_X1 port map( A => n523, Z => n2163);
   U23 : BUF_X1 port map( A => n736, Z => n2130);
   U24 : BUF_X1 port map( A => n736, Z => n2131);
   U25 : BUF_X1 port map( A => n736, Z => n2132);
   U26 : BUF_X1 port map( A => n736, Z => n2133);
   U27 : BUF_X1 port map( A => n736, Z => n2134);
   U28 : BUF_X1 port map( A => n525, Z => n2154);
   U29 : BUF_X1 port map( A => n525, Z => n2155);
   U30 : BUF_X1 port map( A => n525, Z => n2156);
   U31 : BUF_X1 port map( A => n525, Z => n2157);
   U32 : BUF_X1 port map( A => n738, Z => n2128);
   U33 : BUF_X1 port map( A => n738, Z => n2127);
   U34 : BUF_X1 port map( A => n738, Z => n2126);
   U35 : BUF_X1 port map( A => n738, Z => n2125);
   U36 : BUF_X1 port map( A => n738, Z => n2124);
   U37 : BUF_X1 port map( A => n742, Z => n2104);
   U38 : BUF_X1 port map( A => n742, Z => n2103);
   U39 : BUF_X1 port map( A => n742, Z => n2102);
   U40 : BUF_X1 port map( A => n742, Z => n2101);
   U41 : BUF_X1 port map( A => n739, Z => n2122);
   U42 : BUF_X1 port map( A => n739, Z => n2121);
   U43 : BUF_X1 port map( A => n739, Z => n2120);
   U44 : BUF_X1 port map( A => n739, Z => n2119);
   U45 : BUF_X1 port map( A => n739, Z => n2118);
   U46 : BUF_X1 port map( A => n740, Z => n2116);
   U47 : BUF_X1 port map( A => n740, Z => n2115);
   U48 : BUF_X1 port map( A => n740, Z => n2114);
   U49 : BUF_X1 port map( A => n740, Z => n2113);
   U50 : BUF_X1 port map( A => n740, Z => n2112);
   U51 : BUF_X1 port map( A => n741, Z => n2106);
   U52 : BUF_X1 port map( A => n875, Z => n2094);
   U53 : BUF_X1 port map( A => n938, Z => n2082);
   U54 : BUF_X1 port map( A => n978, Z => n2070);
   U55 : BUF_X1 port map( A => n741, Z => n2110);
   U56 : BUF_X1 port map( A => n741, Z => n2109);
   U57 : BUF_X1 port map( A => n741, Z => n2108);
   U58 : BUF_X1 port map( A => n741, Z => n2107);
   U59 : BUF_X1 port map( A => n875, Z => n2098);
   U60 : BUF_X1 port map( A => n875, Z => n2097);
   U61 : BUF_X1 port map( A => n875, Z => n2096);
   U62 : BUF_X1 port map( A => n875, Z => n2095);
   U63 : BUF_X1 port map( A => n938, Z => n2086);
   U64 : BUF_X1 port map( A => n938, Z => n2085);
   U65 : BUF_X1 port map( A => n938, Z => n2084);
   U66 : BUF_X1 port map( A => n938, Z => n2083);
   U67 : BUF_X1 port map( A => n978, Z => n2074);
   U68 : BUF_X1 port map( A => n978, Z => n2073);
   U69 : BUF_X1 port map( A => n978, Z => n2072);
   U70 : BUF_X1 port map( A => n978, Z => n2071);
   U71 : BUF_X1 port map( A => n526, Z => n2148);
   U72 : BUF_X1 port map( A => n526, Z => n2150);
   U73 : BUF_X1 port map( A => n876, Z => n2092);
   U74 : BUF_X1 port map( A => n876, Z => n2091);
   U75 : BUF_X1 port map( A => n876, Z => n2090);
   U76 : BUF_X1 port map( A => n876, Z => n2089);
   U77 : BUF_X1 port map( A => n876, Z => n2088);
   U78 : BUF_X1 port map( A => n939, Z => n2080);
   U79 : BUF_X1 port map( A => n939, Z => n2079);
   U80 : BUF_X1 port map( A => n939, Z => n2078);
   U81 : BUF_X1 port map( A => n939, Z => n2077);
   U82 : BUF_X1 port map( A => n939, Z => n2076);
   U83 : BUF_X1 port map( A => n979, Z => n2068);
   U84 : BUF_X1 port map( A => n979, Z => n2067);
   U85 : BUF_X1 port map( A => n979, Z => n2066);
   U86 : BUF_X1 port map( A => n979, Z => n2065);
   U87 : BUF_X1 port map( A => n979, Z => n2064);
   U88 : BUF_X1 port map( A => n527, Z => n2143);
   U89 : BUF_X1 port map( A => n527, Z => n2142);
   U90 : BUF_X1 port map( A => n526, Z => n2149);
   U91 : BUF_X1 port map( A => n525, Z => n2153);
   U92 : BUF_X1 port map( A => n742, Z => n2100);
   U93 : NAND2_X1 port map( A1 => n734, A2 => n872, ZN => n741);
   U94 : NAND2_X1 port map( A1 => n734, A2 => n936, ZN => n875);
   U95 : NAND2_X1 port map( A1 => n734, A2 => n2094, ZN => n876);
   U96 : NAND2_X1 port map( A1 => n734, A2 => n975, ZN => n938);
   U97 : NAND2_X1 port map( A1 => n734, A2 => n2082, ZN => n939);
   U98 : NAND2_X1 port map( A1 => n734, A2 => n998, ZN => n978);
   U99 : NAND2_X1 port map( A1 => n734, A2 => n2070, ZN => n979);
   U100 : OAI22_X1 port map( A1 => n538, A2 => n2111, B1 => n2104, B2 => n751, 
                           ZN => n1620);
   U101 : OAI22_X1 port map( A1 => n541, A2 => n2110, B1 => n2104, B2 => n753, 
                           ZN => n1618);
   U102 : OAI22_X1 port map( A1 => n544, A2 => n2110, B1 => n2104, B2 => n755, 
                           ZN => n1616);
   U103 : OAI22_X1 port map( A1 => n547, A2 => n2110, B1 => n2104, B2 => n757, 
                           ZN => n1614);
   U104 : OAI22_X1 port map( A1 => n550, A2 => n2110, B1 => n2104, B2 => n759, 
                           ZN => n1612);
   U105 : OAI22_X1 port map( A1 => n553, A2 => n2110, B1 => n2104, B2 => n761, 
                           ZN => n1610);
   U106 : OAI22_X1 port map( A1 => n556, A2 => n2110, B1 => n2104, B2 => n763, 
                           ZN => n1608);
   U107 : OAI22_X1 port map( A1 => n559, A2 => n2110, B1 => n2104, B2 => n765, 
                           ZN => n1606);
   U108 : OAI22_X1 port map( A1 => n562, A2 => n2110, B1 => n2104, B2 => n767, 
                           ZN => n1604);
   U109 : OAI22_X1 port map( A1 => n565, A2 => n2110, B1 => n2104, B2 => n769, 
                           ZN => n1602);
   U110 : OAI22_X1 port map( A1 => n568, A2 => n2110, B1 => n2104, B2 => n771, 
                           ZN => n1600);
   U111 : OAI22_X1 port map( A1 => n571, A2 => n2110, B1 => n2104, B2 => n773, 
                           ZN => n1598);
   U112 : OAI22_X1 port map( A1 => n574, A2 => n2110, B1 => n2103, B2 => n775, 
                           ZN => n1596);
   U113 : OAI22_X1 port map( A1 => n577, A2 => n2109, B1 => n2103, B2 => n777, 
                           ZN => n1594);
   U114 : OAI22_X1 port map( A1 => n580, A2 => n2109, B1 => n2103, B2 => n779, 
                           ZN => n1592);
   U115 : OAI22_X1 port map( A1 => n583, A2 => n2109, B1 => n2103, B2 => n781, 
                           ZN => n1590);
   U116 : OAI22_X1 port map( A1 => n587, A2 => n2109, B1 => n2103, B2 => n783, 
                           ZN => n1588);
   U117 : OAI22_X1 port map( A1 => n591, A2 => n2109, B1 => n2103, B2 => n785, 
                           ZN => n1586);
   U118 : OAI22_X1 port map( A1 => n595, A2 => n2109, B1 => n2103, B2 => n787, 
                           ZN => n1584);
   U119 : OAI22_X1 port map( A1 => n599, A2 => n2109, B1 => n2103, B2 => n789, 
                           ZN => n1582);
   U120 : OAI22_X1 port map( A1 => n603, A2 => n2109, B1 => n2103, B2 => n791, 
                           ZN => n1580);
   U121 : OAI22_X1 port map( A1 => n607, A2 => n2109, B1 => n2103, B2 => n793, 
                           ZN => n1578);
   U122 : OAI22_X1 port map( A1 => n611, A2 => n2109, B1 => n2103, B2 => n795, 
                           ZN => n1576);
   U123 : OAI22_X1 port map( A1 => n615, A2 => n2109, B1 => n2103, B2 => n797, 
                           ZN => n1574);
   U124 : OAI22_X1 port map( A1 => n619, A2 => n2109, B1 => n2102, B2 => n799, 
                           ZN => n1572);
   U125 : OAI22_X1 port map( A1 => n623, A2 => n2108, B1 => n2102, B2 => n801, 
                           ZN => n1570);
   U126 : OAI22_X1 port map( A1 => n626, A2 => n2108, B1 => n2102, B2 => n803, 
                           ZN => n1568);
   U127 : OAI22_X1 port map( A1 => n629, A2 => n2108, B1 => n2102, B2 => n805, 
                           ZN => n1566);
   U128 : OAI22_X1 port map( A1 => n632, A2 => n2108, B1 => n2102, B2 => n807, 
                           ZN => n1564);
   U129 : OAI22_X1 port map( A1 => n635, A2 => n2108, B1 => n2102, B2 => n809, 
                           ZN => n1562);
   U130 : OAI22_X1 port map( A1 => n638, A2 => n2108, B1 => n2102, B2 => n811, 
                           ZN => n1560);
   U131 : OAI22_X1 port map( A1 => n641, A2 => n2108, B1 => n2102, B2 => n813, 
                           ZN => n1558);
   U132 : OAI22_X1 port map( A1 => n644, A2 => n2108, B1 => n2102, B2 => n815, 
                           ZN => n1556);
   U133 : OAI22_X1 port map( A1 => n647, A2 => n2108, B1 => n2102, B2 => n817, 
                           ZN => n1554);
   U134 : OAI22_X1 port map( A1 => n650, A2 => n2108, B1 => n2102, B2 => n819, 
                           ZN => n1552);
   U135 : OAI22_X1 port map( A1 => n653, A2 => n2108, B1 => n2102, B2 => n821, 
                           ZN => n1550);
   U136 : OAI22_X1 port map( A1 => n656, A2 => n2108, B1 => n2101, B2 => n823, 
                           ZN => n1548);
   U137 : OAI22_X1 port map( A1 => n659, A2 => n2107, B1 => n2101, B2 => n825, 
                           ZN => n1546);
   U138 : OAI22_X1 port map( A1 => n662, A2 => n2107, B1 => n2101, B2 => n827, 
                           ZN => n1544);
   U139 : OAI22_X1 port map( A1 => n665, A2 => n2107, B1 => n2101, B2 => n829, 
                           ZN => n1542);
   U140 : OAI22_X1 port map( A1 => n668, A2 => n2107, B1 => n2101, B2 => n831, 
                           ZN => n1540);
   U141 : OAI22_X1 port map( A1 => n671, A2 => n2107, B1 => n2101, B2 => n833, 
                           ZN => n1538);
   U142 : OAI22_X1 port map( A1 => n674, A2 => n2107, B1 => n2101, B2 => n835, 
                           ZN => n1536);
   U143 : OAI22_X1 port map( A1 => n677, A2 => n2107, B1 => n2101, B2 => n837, 
                           ZN => n1534);
   U144 : OAI22_X1 port map( A1 => n680, A2 => n2107, B1 => n2101, B2 => n839, 
                           ZN => n1532);
   U145 : OAI22_X1 port map( A1 => n683, A2 => n2107, B1 => n2101, B2 => n841, 
                           ZN => n1530);
   U146 : OAI22_X1 port map( A1 => n686, A2 => n2107, B1 => n2101, B2 => n843, 
                           ZN => n1528);
   U147 : OAI22_X1 port map( A1 => n689, A2 => n2107, B1 => n2101, B2 => n845, 
                           ZN => n1526);
   U148 : OAI22_X1 port map( A1 => n522, A2 => n2111, B1 => n2105, B2 => n743, 
                           ZN => n1628);
   U149 : OAI22_X1 port map( A1 => n529, A2 => n2111, B1 => n2105, B2 => n745, 
                           ZN => n1626);
   U150 : OAI22_X1 port map( A1 => n532, A2 => n2111, B1 => n2105, B2 => n747, 
                           ZN => n1624);
   U151 : OAI22_X1 port map( A1 => n535, A2 => n2111, B1 => n2105, B2 => n749, 
                           ZN => n1622);
   U152 : OAI22_X1 port map( A1 => n692, A2 => n2107, B1 => n2100, B2 => n847, 
                           ZN => n1524);
   U153 : OAI22_X1 port map( A1 => n696, A2 => n2106, B1 => n2100, B2 => n849, 
                           ZN => n1522);
   U154 : OAI22_X1 port map( A1 => n700, A2 => n2106, B1 => n2100, B2 => n851, 
                           ZN => n1520);
   U155 : OAI22_X1 port map( A1 => n704, A2 => n2106, B1 => n2100, B2 => n853, 
                           ZN => n1518);
   U156 : OAI22_X1 port map( A1 => n707, A2 => n2106, B1 => n2100, B2 => n855, 
                           ZN => n1516);
   U157 : OAI22_X1 port map( A1 => n710, A2 => n2106, B1 => n2100, B2 => n857, 
                           ZN => n1514);
   U158 : OAI22_X1 port map( A1 => n713, A2 => n2106, B1 => n2100, B2 => n859, 
                           ZN => n1512);
   U159 : OAI22_X1 port map( A1 => n716, A2 => n2106, B1 => n2100, B2 => n861, 
                           ZN => n1510);
   U160 : OAI22_X1 port map( A1 => n719, A2 => n2106, B1 => n2100, B2 => n863, 
                           ZN => n1508);
   U161 : OAI22_X1 port map( A1 => n722, A2 => n2106, B1 => n2100, B2 => n865, 
                           ZN => n1506);
   U162 : OAI22_X1 port map( A1 => n725, A2 => n2106, B1 => n2100, B2 => n867, 
                           ZN => n1504);
   U163 : OAI22_X1 port map( A1 => n728, A2 => n2106, B1 => n2100, B2 => n871, 
                           ZN => n1502);
   U164 : AND3_X1 port map( A1 => n2173, A2 => n2174, A3 => n2164, ZN => n526);
   U165 : AND3_X1 port map( A1 => n2164, A2 => n2174, A3 => ADD_RD1(0), ZN => 
                           n527);
   U166 : AND3_X1 port map( A1 => n2164, A2 => n2173, A3 => ADD_RD1(1), ZN => 
                           n525);
   U167 : NAND2_X1 port map( A1 => n734, A2 => n2106, ZN => n742);
   U168 : AND3_X1 port map( A1 => n2135, A2 => n2172, A3 => ADD_RD2(0), ZN => 
                           n740);
   U169 : AND3_X1 port map( A1 => n2135, A2 => n2171, A3 => ADD_RD2(1), ZN => 
                           n738);
   U170 : AND3_X1 port map( A1 => n2171, A2 => n2172, A3 => n2135, ZN => n739);
   U171 : AND2_X1 port map( A1 => RD1, A2 => n734, ZN => n523);
   U172 : AND2_X1 port map( A1 => RD2, A2 => n734, ZN => n736);
   U173 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n873);
   U174 : OAI221_X1 port map( B1 => n2169, B2 => n562, C1 => n1937, C2 => n2160
                           , A => n563, ZN => n1681);
   U175 : AOI222_X1 port map( A1 => n52, A2 => n2153, B1 => n180, B2 => n2149, 
                           C1 => n2146, C2 => n564, ZN => n563);
   U176 : OAI221_X1 port map( B1 => n2169, B2 => n565, C1 => n1936, C2 => n2160
                           , A => n566, ZN => n1680);
   U177 : AOI222_X1 port map( A1 => n51, A2 => n2154, B1 => n179, B2 => n2149, 
                           C1 => n2146, C2 => n567, ZN => n566);
   U178 : OAI221_X1 port map( B1 => n2169, B2 => n568, C1 => n1935, C2 => n2160
                           , A => n569, ZN => n1679);
   U179 : AOI222_X1 port map( A1 => n50, A2 => n2154, B1 => n178, B2 => n2149, 
                           C1 => n2146, C2 => n570, ZN => n569);
   U180 : OAI221_X1 port map( B1 => n2169, B2 => n571, C1 => n1934, C2 => n2161
                           , A => n572, ZN => n1678);
   U181 : AOI222_X1 port map( A1 => n49, A2 => n2154, B1 => n177, B2 => n2149, 
                           C1 => n2145, C2 => n573, ZN => n572);
   U182 : OAI221_X1 port map( B1 => n2168, B2 => n574, C1 => n1933, C2 => n2160
                           , A => n575, ZN => n1677);
   U183 : AOI222_X1 port map( A1 => n48, A2 => n2154, B1 => n176, B2 => n2149, 
                           C1 => n2145, C2 => n576, ZN => n575);
   U184 : OAI221_X1 port map( B1 => n2168, B2 => n577, C1 => n1932, C2 => n2160
                           , A => n578, ZN => n1676);
   U185 : AOI222_X1 port map( A1 => n47, A2 => n2154, B1 => n175, B2 => n2149, 
                           C1 => n2145, C2 => n579, ZN => n578);
   U186 : OAI221_X1 port map( B1 => n2168, B2 => n580, C1 => n1931, C2 => n2160
                           , A => n581, ZN => n1675);
   U187 : AOI222_X1 port map( A1 => n46, A2 => n2154, B1 => n174, B2 => n2149, 
                           C1 => n2145, C2 => n582, ZN => n581);
   U188 : OAI221_X1 port map( B1 => n538, B2 => n2140, C1 => n1881, C2 => n2130
                           , A => n750, ZN => n1621);
   U189 : AOI222_X1 port map( A1 => n2128, A2 => n60, B1 => n2122, B2 => n188, 
                           C1 => n2116, C2 => n540, ZN => n750);
   U190 : OAI221_X1 port map( B1 => n541, B2 => n2140, C1 => n1880, C2 => n2130
                           , A => n752, ZN => n1619);
   U191 : AOI222_X1 port map( A1 => n2128, A2 => n59, B1 => n2122, B2 => n187, 
                           C1 => n2116, C2 => n543, ZN => n752);
   U192 : OAI221_X1 port map( B1 => n544, B2 => n2140, C1 => n1879, C2 => n2130
                           , A => n754, ZN => n1617);
   U193 : AOI222_X1 port map( A1 => n2128, A2 => n58, B1 => n2122, B2 => n186, 
                           C1 => n2116, C2 => n546, ZN => n754);
   U194 : OAI221_X1 port map( B1 => n547, B2 => n2140, C1 => n1878, C2 => n2130
                           , A => n756, ZN => n1615);
   U195 : AOI222_X1 port map( A1 => n2128, A2 => n57, B1 => n2122, B2 => n185, 
                           C1 => n2116, C2 => n549, ZN => n756);
   U196 : OAI221_X1 port map( B1 => n550, B2 => n2140, C1 => n1877, C2 => n2130
                           , A => n758, ZN => n1613);
   U197 : AOI222_X1 port map( A1 => n2128, A2 => n56, B1 => n2122, B2 => n184, 
                           C1 => n2116, C2 => n552, ZN => n758);
   U198 : OAI221_X1 port map( B1 => n553, B2 => n2140, C1 => n1876, C2 => n2130
                           , A => n760, ZN => n1611);
   U199 : AOI222_X1 port map( A1 => n2128, A2 => n55, B1 => n2122, B2 => n183, 
                           C1 => n2116, C2 => n555, ZN => n760);
   U200 : OAI221_X1 port map( B1 => n556, B2 => n2140, C1 => n1875, C2 => n2130
                           , A => n762, ZN => n1609);
   U201 : AOI222_X1 port map( A1 => n2128, A2 => n54, B1 => n2122, B2 => n182, 
                           C1 => n2116, C2 => n558, ZN => n762);
   U202 : OAI221_X1 port map( B1 => n559, B2 => n2140, C1 => n1874, C2 => n2130
                           , A => n764, ZN => n1607);
   U203 : AOI222_X1 port map( A1 => n2128, A2 => n53, B1 => n2122, B2 => n181, 
                           C1 => n2116, C2 => n561, ZN => n764);
   U204 : OAI221_X1 port map( B1 => n562, B2 => n2140, C1 => n1873, C2 => n2131
                           , A => n766, ZN => n1605);
   U205 : AOI222_X1 port map( A1 => n2128, A2 => n52, B1 => n2122, B2 => n180, 
                           C1 => n2116, C2 => n564, ZN => n766);
   U206 : OAI221_X1 port map( B1 => n565, B2 => n2140, C1 => n1872, C2 => n2131
                           , A => n768, ZN => n1603);
   U207 : AOI222_X1 port map( A1 => n2128, A2 => n51, B1 => n2122, B2 => n179, 
                           C1 => n2116, C2 => n567, ZN => n768);
   U208 : OAI221_X1 port map( B1 => n568, B2 => n2140, C1 => n1871, C2 => n2131
                           , A => n770, ZN => n1601);
   U209 : AOI222_X1 port map( A1 => n2128, A2 => n50, B1 => n2122, B2 => n178, 
                           C1 => n2116, C2 => n570, ZN => n770);
   U210 : OAI221_X1 port map( B1 => n571, B2 => n2140, C1 => n1870, C2 => n2132
                           , A => n772, ZN => n1599);
   U211 : AOI222_X1 port map( A1 => n2128, A2 => n49, B1 => n2122, B2 => n177, 
                           C1 => n2116, C2 => n573, ZN => n772);
   U212 : OAI221_X1 port map( B1 => n574, B2 => n2139, C1 => n1869, C2 => n2131
                           , A => n774, ZN => n1597);
   U213 : AOI222_X1 port map( A1 => n2127, A2 => n48, B1 => n2121, B2 => n176, 
                           C1 => n2115, C2 => n576, ZN => n774);
   U214 : OAI221_X1 port map( B1 => n577, B2 => n2139, C1 => n1868, C2 => n2131
                           , A => n776, ZN => n1595);
   U215 : AOI222_X1 port map( A1 => n2127, A2 => n47, B1 => n2121, B2 => n175, 
                           C1 => n2115, C2 => n579, ZN => n776);
   U216 : OAI221_X1 port map( B1 => n580, B2 => n2139, C1 => n1867, C2 => n2131
                           , A => n778, ZN => n1593);
   U217 : AOI222_X1 port map( A1 => n2127, A2 => n46, B1 => n2121, B2 => n174, 
                           C1 => n2115, C2 => n582, ZN => n778);
   U218 : OAI221_X1 port map( B1 => n2166, B2 => n656, C1 => n1909, C2 => n2162
                           , A => n657, ZN => n1653);
   U219 : AOI222_X1 port map( A1 => n24, A2 => n2156, B1 => n2151, B2 => n658, 
                           C1 => n88, C2 => n2143, ZN => n657);
   U220 : OAI221_X1 port map( B1 => n2166, B2 => n659, C1 => n1908, C2 => n2162
                           , A => n660, ZN => n1652);
   U221 : AOI222_X1 port map( A1 => n23, A2 => n2156, B1 => n2151, B2 => n661, 
                           C1 => n87, C2 => n2143, ZN => n660);
   U222 : OAI221_X1 port map( B1 => n2166, B2 => n662, C1 => n1907, C2 => n2162
                           , A => n663, ZN => n1651);
   U223 : AOI222_X1 port map( A1 => n22, A2 => n2156, B1 => n2151, B2 => n664, 
                           C1 => n86, C2 => n2143, ZN => n663);
   U224 : OAI221_X1 port map( B1 => n2166, B2 => n665, C1 => n1906, C2 => n2162
                           , A => n666, ZN => n1650);
   U225 : AOI222_X1 port map( A1 => n21, A2 => n2156, B1 => n2151, B2 => n667, 
                           C1 => n85, C2 => n2143, ZN => n666);
   U226 : OAI221_X1 port map( B1 => n2166, B2 => n668, C1 => n1905, C2 => n2162
                           , A => n669, ZN => n1649);
   U227 : AOI222_X1 port map( A1 => n20, A2 => n2156, B1 => n2151, B2 => n670, 
                           C1 => n84, C2 => n2143, ZN => n669);
   U228 : OAI221_X1 port map( B1 => n2166, B2 => n671, C1 => n1904, C2 => n2162
                           , A => n672, ZN => n1648);
   U229 : AOI222_X1 port map( A1 => n19, A2 => n2156, B1 => n2151, B2 => n673, 
                           C1 => n83, C2 => n2143, ZN => n672);
   U230 : OAI221_X1 port map( B1 => n2166, B2 => n674, C1 => n1903, C2 => n2162
                           , A => n675, ZN => n1647);
   U231 : AOI222_X1 port map( A1 => n18, A2 => n2156, B1 => n2151, B2 => n676, 
                           C1 => n82, C2 => n2143, ZN => n675);
   U232 : OAI221_X1 port map( B1 => n2166, B2 => n677, C1 => n1902, C2 => n2162
                           , A => n678, ZN => n1646);
   U233 : AOI222_X1 port map( A1 => n17, A2 => n2156, B1 => n2151, B2 => n679, 
                           C1 => n81, C2 => n2143, ZN => n678);
   U234 : OAI221_X1 port map( B1 => n2166, B2 => n680, C1 => n1901, C2 => n2163
                           , A => n681, ZN => n1645);
   U235 : AOI222_X1 port map( A1 => n16, A2 => n2157, B1 => n2151, B2 => n682, 
                           C1 => n80, C2 => n2143, ZN => n681);
   U236 : OAI221_X1 port map( B1 => n2166, B2 => n683, C1 => n1900, C2 => n2163
                           , A => n684, ZN => n1644);
   U237 : AOI222_X1 port map( A1 => n15, A2 => n2157, B1 => n2151, B2 => n685, 
                           C1 => n79, C2 => n2143, ZN => n684);
   U238 : OAI221_X1 port map( B1 => n2166, B2 => n686, C1 => n1899, C2 => n2163
                           , A => n687, ZN => n1643);
   U239 : AOI222_X1 port map( A1 => n14, A2 => n2157, B1 => n2152, B2 => n688, 
                           C1 => n78, C2 => n2143, ZN => n687);
   U240 : OAI221_X1 port map( B1 => n2166, B2 => n689, C1 => n1898, C2 => n2163
                           , A => n690, ZN => n1642);
   U241 : AOI222_X1 port map( A1 => n13, A2 => n2157, B1 => n2152, B2 => n691, 
                           C1 => n77, C2 => n2143, ZN => n690);
   U242 : OAI221_X1 port map( B1 => n2165, B2 => n692, C1 => n1897, C2 => n2163
                           , A => n693, ZN => n1641);
   U243 : AOI222_X1 port map( A1 => n2158, A2 => n694, B1 => n2152, B2 => n695,
                           C1 => n76, C2 => n2142, ZN => n693);
   U244 : OAI221_X1 port map( B1 => n2165, B2 => n696, C1 => n1896, C2 => n2163
                           , A => n697, ZN => n1640);
   U245 : AOI222_X1 port map( A1 => n2158, A2 => n698, B1 => n2152, B2 => n699,
                           C1 => n75, C2 => n2142, ZN => n697);
   U246 : OAI221_X1 port map( B1 => n2165, B2 => n700, C1 => n1895, C2 => n2163
                           , A => n701, ZN => n1639);
   U247 : AOI222_X1 port map( A1 => n2158, A2 => n702, B1 => n2152, B2 => n703,
                           C1 => n74, C2 => n2142, ZN => n701);
   U248 : OAI221_X1 port map( B1 => n2165, B2 => n704, C1 => n1894, C2 => n2163
                           , A => n705, ZN => n1638);
   U249 : AOI222_X1 port map( A1 => n9, A2 => n2157, B1 => n2152, B2 => n706, 
                           C1 => n73, C2 => n2142, ZN => n705);
   U250 : OAI221_X1 port map( B1 => n2165, B2 => n707, C1 => n1893, C2 => n2163
                           , A => n708, ZN => n1637);
   U251 : AOI222_X1 port map( A1 => n8, A2 => n2157, B1 => n2152, B2 => n709, 
                           C1 => n72, C2 => n2142, ZN => n708);
   U252 : OAI221_X1 port map( B1 => n2165, B2 => n710, C1 => n1892, C2 => n2163
                           , A => n711, ZN => n1636);
   U253 : AOI222_X1 port map( A1 => n7, A2 => n2157, B1 => n2152, B2 => n712, 
                           C1 => n71, C2 => n2142, ZN => n711);
   U254 : OAI221_X1 port map( B1 => n2165, B2 => n713, C1 => n1891, C2 => n2163
                           , A => n714, ZN => n1635);
   U255 : AOI222_X1 port map( A1 => n6, A2 => n2157, B1 => n2152, B2 => n715, 
                           C1 => n70, C2 => n2142, ZN => n714);
   U256 : OAI221_X1 port map( B1 => n2165, B2 => n719, C1 => n1889, C2 => n2163
                           , A => n720, ZN => n1633);
   U257 : AOI222_X1 port map( A1 => n4, A2 => n2157, B1 => n2152, B2 => n721, 
                           C1 => n68, C2 => n2142, ZN => n720);
   U258 : OAI221_X1 port map( B1 => n2165, B2 => n728, C1 => n1886, C2 => n2164
                           , A => n729, ZN => n1630);
   U259 : AOI222_X1 port map( A1 => n2158, A2 => n730, B1 => n2148, B2 => n731,
                           C1 => n65, C2 => n2142, ZN => n729);
   U260 : OAI221_X1 port map( B1 => n623, B2 => n2138, C1 => n1856, C2 => n2132
                           , A => n800, ZN => n1571);
   U261 : AOI222_X1 port map( A1 => n2126, A2 => n35, B1 => n2120, B2 => n625, 
                           C1 => n2114, C2 => n99, ZN => n800);
   U262 : OAI221_X1 port map( B1 => n626, B2 => n2138, C1 => n1855, C2 => n2132
                           , A => n802, ZN => n1569);
   U263 : AOI222_X1 port map( A1 => n2126, A2 => n34, B1 => n2120, B2 => n628, 
                           C1 => n2114, C2 => n98, ZN => n802);
   U264 : OAI221_X1 port map( B1 => n629, B2 => n2138, C1 => n1854, C2 => n2132
                           , A => n804, ZN => n1567);
   U265 : AOI222_X1 port map( A1 => n2126, A2 => n33, B1 => n2120, B2 => n631, 
                           C1 => n2114, C2 => n97, ZN => n804);
   U266 : OAI221_X1 port map( B1 => n632, B2 => n2138, C1 => n1853, C2 => n2132
                           , A => n806, ZN => n1565);
   U267 : AOI222_X1 port map( A1 => n2126, A2 => n32, B1 => n2120, B2 => n634, 
                           C1 => n2114, C2 => n96, ZN => n806);
   U268 : OAI221_X1 port map( B1 => n635, B2 => n2138, C1 => n1852, C2 => n2132
                           , A => n808, ZN => n1563);
   U269 : AOI222_X1 port map( A1 => n2126, A2 => n31, B1 => n2120, B2 => n637, 
                           C1 => n2114, C2 => n95, ZN => n808);
   U270 : OAI221_X1 port map( B1 => n638, B2 => n2138, C1 => n1851, C2 => n2132
                           , A => n810, ZN => n1561);
   U271 : AOI222_X1 port map( A1 => n2126, A2 => n30, B1 => n2120, B2 => n640, 
                           C1 => n2114, C2 => n94, ZN => n810);
   U272 : OAI221_X1 port map( B1 => n641, B2 => n2138, C1 => n1850, C2 => n2132
                           , A => n812, ZN => n1559);
   U273 : AOI222_X1 port map( A1 => n2126, A2 => n29, B1 => n2120, B2 => n643, 
                           C1 => n2114, C2 => n93, ZN => n812);
   U274 : OAI221_X1 port map( B1 => n644, B2 => n2138, C1 => n1849, C2 => n2133
                           , A => n814, ZN => n1557);
   U275 : AOI222_X1 port map( A1 => n2126, A2 => n28, B1 => n2120, B2 => n646, 
                           C1 => n2114, C2 => n92, ZN => n814);
   U276 : OAI221_X1 port map( B1 => n647, B2 => n2138, C1 => n1848, C2 => n2133
                           , A => n816, ZN => n1555);
   U277 : AOI222_X1 port map( A1 => n2126, A2 => n27, B1 => n2120, B2 => n649, 
                           C1 => n2114, C2 => n91, ZN => n816);
   U278 : OAI221_X1 port map( B1 => n650, B2 => n2138, C1 => n1847, C2 => n2133
                           , A => n818, ZN => n1553);
   U279 : AOI222_X1 port map( A1 => n2126, A2 => n26, B1 => n2120, B2 => n652, 
                           C1 => n2114, C2 => n90, ZN => n818);
   U280 : OAI221_X1 port map( B1 => n653, B2 => n2138, C1 => n1846, C2 => n2133
                           , A => n820, ZN => n1551);
   U281 : AOI222_X1 port map( A1 => n2126, A2 => n25, B1 => n2120, B2 => n655, 
                           C1 => n2114, C2 => n89, ZN => n820);
   U282 : OAI221_X1 port map( B1 => n656, B2 => n2137, C1 => n1845, C2 => n2133
                           , A => n822, ZN => n1549);
   U283 : AOI222_X1 port map( A1 => n2125, A2 => n24, B1 => n2119, B2 => n658, 
                           C1 => n2113, C2 => n88, ZN => n822);
   U284 : OAI221_X1 port map( B1 => n659, B2 => n2137, C1 => n1844, C2 => n2133
                           , A => n824, ZN => n1547);
   U285 : AOI222_X1 port map( A1 => n2125, A2 => n23, B1 => n2119, B2 => n661, 
                           C1 => n2113, C2 => n87, ZN => n824);
   U286 : OAI221_X1 port map( B1 => n662, B2 => n2137, C1 => n1843, C2 => n2133
                           , A => n826, ZN => n1545);
   U287 : AOI222_X1 port map( A1 => n2125, A2 => n22, B1 => n2119, B2 => n664, 
                           C1 => n2113, C2 => n86, ZN => n826);
   U288 : OAI221_X1 port map( B1 => n665, B2 => n2137, C1 => n1842, C2 => n2133
                           , A => n828, ZN => n1543);
   U289 : AOI222_X1 port map( A1 => n2125, A2 => n21, B1 => n2119, B2 => n667, 
                           C1 => n2113, C2 => n85, ZN => n828);
   U290 : OAI221_X1 port map( B1 => n668, B2 => n2137, C1 => n1841, C2 => n2133
                           , A => n830, ZN => n1541);
   U291 : AOI222_X1 port map( A1 => n2125, A2 => n20, B1 => n2119, B2 => n670, 
                           C1 => n2113, C2 => n84, ZN => n830);
   U292 : OAI221_X1 port map( B1 => n671, B2 => n2137, C1 => n1840, C2 => n2133
                           , A => n832, ZN => n1539);
   U293 : AOI222_X1 port map( A1 => n2125, A2 => n19, B1 => n2119, B2 => n673, 
                           C1 => n2113, C2 => n83, ZN => n832);
   U294 : OAI221_X1 port map( B1 => n674, B2 => n2137, C1 => n1839, C2 => n2133
                           , A => n834, ZN => n1537);
   U295 : AOI222_X1 port map( A1 => n2125, A2 => n18, B1 => n2119, B2 => n676, 
                           C1 => n2113, C2 => n82, ZN => n834);
   U296 : OAI221_X1 port map( B1 => n677, B2 => n2137, C1 => n1838, C2 => n2133
                           , A => n836, ZN => n1535);
   U297 : AOI222_X1 port map( A1 => n2125, A2 => n17, B1 => n2119, B2 => n679, 
                           C1 => n2113, C2 => n81, ZN => n836);
   U298 : OAI221_X1 port map( B1 => n680, B2 => n2137, C1 => n1837, C2 => n2134
                           , A => n838, ZN => n1533);
   U299 : AOI222_X1 port map( A1 => n2125, A2 => n16, B1 => n2119, B2 => n682, 
                           C1 => n2113, C2 => n80, ZN => n838);
   U300 : OAI221_X1 port map( B1 => n683, B2 => n2137, C1 => n1836, C2 => n2134
                           , A => n840, ZN => n1531);
   U301 : AOI222_X1 port map( A1 => n2125, A2 => n15, B1 => n2119, B2 => n685, 
                           C1 => n2113, C2 => n79, ZN => n840);
   U302 : OAI221_X1 port map( B1 => n686, B2 => n2137, C1 => n1835, C2 => n2134
                           , A => n842, ZN => n1529);
   U303 : AOI222_X1 port map( A1 => n2125, A2 => n14, B1 => n2119, B2 => n688, 
                           C1 => n2113, C2 => n78, ZN => n842);
   U304 : OAI221_X1 port map( B1 => n689, B2 => n2137, C1 => n1834, C2 => n2134
                           , A => n844, ZN => n1527);
   U305 : AOI222_X1 port map( A1 => n2125, A2 => n13, B1 => n2119, B2 => n691, 
                           C1 => n2113, C2 => n77, ZN => n844);
   U306 : OAI221_X1 port map( B1 => n692, B2 => n2136, C1 => n1833, C2 => n2134
                           , A => n846, ZN => n1525);
   U307 : AOI222_X1 port map( A1 => n2124, A2 => n694, B1 => n2118, B2 => n695,
                           C1 => n2112, C2 => n76, ZN => n846);
   U308 : OAI221_X1 port map( B1 => n696, B2 => n2136, C1 => n1832, C2 => n2134
                           , A => n848, ZN => n1523);
   U309 : AOI222_X1 port map( A1 => n2124, A2 => n698, B1 => n2118, B2 => n699,
                           C1 => n2112, C2 => n75, ZN => n848);
   U310 : OAI221_X1 port map( B1 => n700, B2 => n2136, C1 => n1831, C2 => n2134
                           , A => n850, ZN => n1521);
   U311 : AOI222_X1 port map( A1 => n2124, A2 => n702, B1 => n2118, B2 => n703,
                           C1 => n2112, C2 => n74, ZN => n850);
   U312 : OAI221_X1 port map( B1 => n704, B2 => n2136, C1 => n1830, C2 => n2134
                           , A => n852, ZN => n1519);
   U313 : AOI222_X1 port map( A1 => n2124, A2 => n9, B1 => n2118, B2 => n706, 
                           C1 => n2112, C2 => n73, ZN => n852);
   U314 : OAI221_X1 port map( B1 => n707, B2 => n2136, C1 => n1829, C2 => n2134
                           , A => n854, ZN => n1517);
   U315 : AOI222_X1 port map( A1 => n2124, A2 => n8, B1 => n2118, B2 => n709, 
                           C1 => n2112, C2 => n72, ZN => n854);
   U316 : OAI221_X1 port map( B1 => n710, B2 => n2136, C1 => n1828, C2 => n2134
                           , A => n856, ZN => n1515);
   U317 : AOI222_X1 port map( A1 => n2124, A2 => n7, B1 => n2118, B2 => n712, 
                           C1 => n2112, C2 => n71, ZN => n856);
   U318 : OAI221_X1 port map( B1 => n713, B2 => n2136, C1 => n1827, C2 => n2134
                           , A => n858, ZN => n1513);
   U319 : AOI222_X1 port map( A1 => n2124, A2 => n6, B1 => n2118, B2 => n715, 
                           C1 => n2112, C2 => n70, ZN => n858);
   U320 : OAI221_X1 port map( B1 => n716, B2 => n2136, C1 => n1826, C2 => n2135
                           , A => n860, ZN => n1511);
   U321 : AOI222_X1 port map( A1 => n2124, A2 => n5, B1 => n2118, B2 => n718, 
                           C1 => n2112, C2 => n69, ZN => n860);
   U322 : OAI221_X1 port map( B1 => n719, B2 => n2136, C1 => n1825, C2 => n2134
                           , A => n862, ZN => n1509);
   U323 : AOI222_X1 port map( A1 => n2124, A2 => n4, B1 => n2118, B2 => n721, 
                           C1 => n2112, C2 => n68, ZN => n862);
   U324 : OAI221_X1 port map( B1 => n722, B2 => n2136, C1 => n1824, C2 => n2135
                           , A => n864, ZN => n1507);
   U325 : AOI222_X1 port map( A1 => n2124, A2 => n3, B1 => n2118, B2 => n724, 
                           C1 => n2112, C2 => n67, ZN => n864);
   U326 : OAI221_X1 port map( B1 => n725, B2 => n2136, C1 => n1823, C2 => n2135
                           , A => n866, ZN => n1505);
   U327 : AOI222_X1 port map( A1 => n2124, A2 => n2, B1 => n2118, B2 => n727, 
                           C1 => n2112, C2 => n66, ZN => n866);
   U328 : OAI221_X1 port map( B1 => n728, B2 => n2136, C1 => n1822, C2 => n2135
                           , A => n868, ZN => n1503);
   U329 : AOI222_X1 port map( A1 => n2124, A2 => n730, B1 => n2118, B2 => n731,
                           C1 => n2112, C2 => n65, ZN => n868);
   U330 : INV_X1 port map( A => RESET, ZN => n734);
   U331 : OAI221_X1 port map( B1 => n2170, B2 => n522, C1 => n1949, C2 => n2159
                           , A => n524, ZN => n1693);
   U332 : AOI222_X1 port map( A1 => n64, A2 => n2155, B1 => n192, B2 => n2148, 
                           C1 => n2147, C2 => n528, ZN => n524);
   U333 : OAI221_X1 port map( B1 => n2170, B2 => n529, C1 => n1948, C2 => n2159
                           , A => n530, ZN => n1692);
   U334 : AOI222_X1 port map( A1 => n63, A2 => n2153, B1 => n191, B2 => n2148, 
                           C1 => n2147, C2 => n531, ZN => n530);
   U335 : OAI221_X1 port map( B1 => n2170, B2 => n532, C1 => n1947, C2 => n2159
                           , A => n533, ZN => n1691);
   U336 : AOI222_X1 port map( A1 => n62, A2 => n2153, B1 => n190, B2 => n2148, 
                           C1 => n2146, C2 => n534, ZN => n533);
   U337 : OAI221_X1 port map( B1 => n2170, B2 => n535, C1 => n1946, C2 => n2159
                           , A => n536, ZN => n1690);
   U338 : AOI222_X1 port map( A1 => n61, A2 => n2153, B1 => n189, B2 => n2148, 
                           C1 => n2146, C2 => n537, ZN => n536);
   U339 : OAI221_X1 port map( B1 => n2167, B2 => n619, C1 => n1921, C2 => n2161
                           , A => n620, ZN => n1665);
   U340 : AOI222_X1 port map( A1 => n36, A2 => n2155, B1 => n2150, B2 => n621, 
                           C1 => n2144, C2 => n622, ZN => n620);
   U341 : OAI221_X1 port map( B1 => n2167, B2 => n623, C1 => n1920, C2 => n2161
                           , A => n624, ZN => n1664);
   U342 : AOI222_X1 port map( A1 => n35, A2 => n2155, B1 => n2150, B2 => n625, 
                           C1 => n99, C2 => n2144, ZN => n624);
   U343 : OAI221_X1 port map( B1 => n2167, B2 => n626, C1 => n1919, C2 => n2161
                           , A => n627, ZN => n1663);
   U344 : AOI222_X1 port map( A1 => n34, A2 => n2155, B1 => n2150, B2 => n628, 
                           C1 => n98, C2 => n2144, ZN => n627);
   U345 : OAI221_X1 port map( B1 => n2167, B2 => n629, C1 => n1918, C2 => n2161
                           , A => n630, ZN => n1662);
   U346 : AOI222_X1 port map( A1 => n33, A2 => n2155, B1 => n2150, B2 => n631, 
                           C1 => n97, C2 => n2144, ZN => n630);
   U347 : OAI221_X1 port map( B1 => n2167, B2 => n632, C1 => n1917, C2 => n2161
                           , A => n633, ZN => n1661);
   U348 : AOI222_X1 port map( A1 => n32, A2 => n2155, B1 => n2150, B2 => n634, 
                           C1 => n96, C2 => n2144, ZN => n633);
   U349 : OAI221_X1 port map( B1 => n2167, B2 => n635, C1 => n1916, C2 => n2161
                           , A => n636, ZN => n1660);
   U350 : AOI222_X1 port map( A1 => n31, A2 => n2155, B1 => n2150, B2 => n637, 
                           C1 => n95, C2 => n2144, ZN => n636);
   U351 : OAI221_X1 port map( B1 => n2167, B2 => n638, C1 => n1915, C2 => n2161
                           , A => n639, ZN => n1659);
   U352 : AOI222_X1 port map( A1 => n30, A2 => n2155, B1 => n2150, B2 => n640, 
                           C1 => n94, C2 => n2144, ZN => n639);
   U353 : OAI221_X1 port map( B1 => n2167, B2 => n641, C1 => n1914, C2 => n2161
                           , A => n642, ZN => n1658);
   U354 : AOI222_X1 port map( A1 => n29, A2 => n2155, B1 => n2150, B2 => n643, 
                           C1 => n93, C2 => n2144, ZN => n642);
   U355 : OAI221_X1 port map( B1 => n2167, B2 => n644, C1 => n1913, C2 => n2162
                           , A => n645, ZN => n1657);
   U356 : AOI222_X1 port map( A1 => n28, A2 => n2156, B1 => n2150, B2 => n646, 
                           C1 => n92, C2 => n2144, ZN => n645);
   U357 : OAI221_X1 port map( B1 => n2167, B2 => n647, C1 => n1912, C2 => n2162
                           , A => n648, ZN => n1656);
   U358 : AOI222_X1 port map( A1 => n27, A2 => n2156, B1 => n2151, B2 => n649, 
                           C1 => n91, C2 => n2144, ZN => n648);
   U359 : OAI221_X1 port map( B1 => n2167, B2 => n650, C1 => n1911, C2 => n2162
                           , A => n651, ZN => n1655);
   U360 : AOI222_X1 port map( A1 => n26, A2 => n2156, B1 => n2151, B2 => n652, 
                           C1 => n90, C2 => n2144, ZN => n651);
   U361 : OAI221_X1 port map( B1 => n2167, B2 => n653, C1 => n1910, C2 => n2162
                           , A => n654, ZN => n1654);
   U362 : AOI222_X1 port map( A1 => n25, A2 => n2156, B1 => n2151, B2 => n655, 
                           C1 => n89, C2 => n2144, ZN => n654);
   U363 : OAI221_X1 port map( B1 => n2165, B2 => n716, C1 => n1890, C2 => n2164
                           , A => n717, ZN => n1634);
   U364 : AOI222_X1 port map( A1 => n5, A2 => n2157, B1 => n2152, B2 => n718, 
                           C1 => n69, C2 => n2142, ZN => n717);
   U365 : OAI221_X1 port map( B1 => n2165, B2 => n722, C1 => n1888, C2 => n2164
                           , A => n723, ZN => n1632);
   U366 : AOI222_X1 port map( A1 => n3, A2 => n2157, B1 => n2152, B2 => n724, 
                           C1 => n67, C2 => n2142, ZN => n723);
   U367 : OAI221_X1 port map( B1 => n2165, B2 => n725, C1 => n1887, C2 => n2164
                           , A => n726, ZN => n1631);
   U368 : AOI222_X1 port map( A1 => n2, A2 => n2157, B1 => n2152, B2 => n727, 
                           C1 => n66, C2 => n2142, ZN => n726);
   U369 : OAI221_X1 port map( B1 => n522, B2 => n2141, C1 => n1885, C2 => n2130
                           , A => n737, ZN => n1629);
   U370 : AOI222_X1 port map( A1 => n2129, A2 => n64, B1 => n2123, B2 => n192, 
                           C1 => n2117, C2 => n528, ZN => n737);
   U371 : OAI221_X1 port map( B1 => n529, B2 => n2141, C1 => n1884, C2 => n2130
                           , A => n744, ZN => n1627);
   U372 : AOI222_X1 port map( A1 => n2129, A2 => n63, B1 => n2123, B2 => n191, 
                           C1 => n2117, C2 => n531, ZN => n744);
   U373 : OAI221_X1 port map( B1 => n532, B2 => n2141, C1 => n1883, C2 => n2130
                           , A => n746, ZN => n1625);
   U374 : AOI222_X1 port map( A1 => n2129, A2 => n62, B1 => n2123, B2 => n190, 
                           C1 => n2117, C2 => n534, ZN => n746);
   U375 : OAI221_X1 port map( B1 => n535, B2 => n2141, C1 => n1882, C2 => n2130
                           , A => n748, ZN => n1623);
   U376 : AOI222_X1 port map( A1 => n2129, A2 => n61, B1 => n2123, B2 => n189, 
                           C1 => n2117, C2 => n537, ZN => n748);
   U377 : OAI221_X1 port map( B1 => n583, B2 => n2139, C1 => n1866, C2 => n2131
                           , A => n780, ZN => n1591);
   U378 : AOI222_X1 port map( A1 => n2127, A2 => n45, B1 => n2121, B2 => n585, 
                           C1 => n2115, C2 => n586, ZN => n780);
   U379 : OAI221_X1 port map( B1 => n587, B2 => n2139, C1 => n1865, C2 => n2131
                           , A => n782, ZN => n1589);
   U380 : AOI222_X1 port map( A1 => n2127, A2 => n44, B1 => n2121, B2 => n589, 
                           C1 => n2115, C2 => n590, ZN => n782);
   U381 : OAI221_X1 port map( B1 => n591, B2 => n2139, C1 => n1864, C2 => n2131
                           , A => n784, ZN => n1587);
   U382 : AOI222_X1 port map( A1 => n2127, A2 => n43, B1 => n2121, B2 => n593, 
                           C1 => n2115, C2 => n594, ZN => n784);
   U383 : OAI221_X1 port map( B1 => n595, B2 => n2139, C1 => n1863, C2 => n2131
                           , A => n786, ZN => n1585);
   U384 : AOI222_X1 port map( A1 => n2127, A2 => n42, B1 => n2121, B2 => n597, 
                           C1 => n2115, C2 => n598, ZN => n786);
   U385 : OAI221_X1 port map( B1 => n599, B2 => n2139, C1 => n1862, C2 => n2131
                           , A => n788, ZN => n1583);
   U386 : AOI222_X1 port map( A1 => n2127, A2 => n41, B1 => n2121, B2 => n601, 
                           C1 => n2115, C2 => n602, ZN => n788);
   U387 : OAI221_X1 port map( B1 => n603, B2 => n2139, C1 => n1861, C2 => n2131
                           , A => n790, ZN => n1581);
   U388 : AOI222_X1 port map( A1 => n2127, A2 => n40, B1 => n2121, B2 => n605, 
                           C1 => n2115, C2 => n606, ZN => n790);
   U389 : OAI221_X1 port map( B1 => n607, B2 => n2139, C1 => n1860, C2 => n2132
                           , A => n792, ZN => n1579);
   U390 : AOI222_X1 port map( A1 => n2127, A2 => n39, B1 => n2121, B2 => n609, 
                           C1 => n2115, C2 => n610, ZN => n792);
   U391 : OAI221_X1 port map( B1 => n611, B2 => n2139, C1 => n1859, C2 => n2132
                           , A => n794, ZN => n1577);
   U392 : AOI222_X1 port map( A1 => n2127, A2 => n38, B1 => n2121, B2 => n613, 
                           C1 => n2115, C2 => n614, ZN => n794);
   U393 : OAI221_X1 port map( B1 => n615, B2 => n2139, C1 => n1858, C2 => n2132
                           , A => n796, ZN => n1575);
   U394 : AOI222_X1 port map( A1 => n2127, A2 => n37, B1 => n2121, B2 => n617, 
                           C1 => n2115, C2 => n618, ZN => n796);
   U395 : OAI221_X1 port map( B1 => n619, B2 => n2138, C1 => n1857, C2 => n2132
                           , A => n798, ZN => n1573);
   U396 : AOI222_X1 port map( A1 => n2126, A2 => n36, B1 => n2120, B2 => n621, 
                           C1 => n2114, C2 => n622, ZN => n798);
   U397 : OAI221_X1 port map( B1 => n2169, B2 => n538, C1 => n1945, C2 => n2159
                           , A => n539, ZN => n1689);
   U398 : AOI222_X1 port map( A1 => n60, A2 => n2153, B1 => n188, B2 => n2148, 
                           C1 => n2146, C2 => n540, ZN => n539);
   U399 : OAI221_X1 port map( B1 => n2169, B2 => n541, C1 => n1944, C2 => n2159
                           , A => n542, ZN => n1688);
   U400 : AOI222_X1 port map( A1 => n59, A2 => n2153, B1 => n187, B2 => n2148, 
                           C1 => n2146, C2 => n543, ZN => n542);
   U401 : OAI221_X1 port map( B1 => n2169, B2 => n544, C1 => n1943, C2 => n2159
                           , A => n545, ZN => n1687);
   U402 : AOI222_X1 port map( A1 => n58, A2 => n2153, B1 => n186, B2 => n2148, 
                           C1 => n2146, C2 => n546, ZN => n545);
   U403 : OAI221_X1 port map( B1 => n2169, B2 => n547, C1 => n1942, C2 => n2159
                           , A => n548, ZN => n1686);
   U404 : AOI222_X1 port map( A1 => n57, A2 => n2153, B1 => n185, B2 => n2148, 
                           C1 => n2146, C2 => n549, ZN => n548);
   U405 : OAI221_X1 port map( B1 => n2169, B2 => n550, C1 => n1941, C2 => n2159
                           , A => n551, ZN => n1685);
   U406 : AOI222_X1 port map( A1 => n56, A2 => n2153, B1 => n184, B2 => n2148, 
                           C1 => n2146, C2 => n552, ZN => n551);
   U407 : OAI221_X1 port map( B1 => n2169, B2 => n553, C1 => n1940, C2 => n2159
                           , A => n554, ZN => n1684);
   U408 : AOI222_X1 port map( A1 => n55, A2 => n2153, B1 => n183, B2 => n2148, 
                           C1 => n2146, C2 => n555, ZN => n554);
   U409 : OAI221_X1 port map( B1 => n2169, B2 => n556, C1 => n1939, C2 => n2159
                           , A => n557, ZN => n1683);
   U410 : AOI222_X1 port map( A1 => n54, A2 => n2153, B1 => n182, B2 => n2148, 
                           C1 => n2146, C2 => n558, ZN => n557);
   U411 : OAI221_X1 port map( B1 => n2169, B2 => n559, C1 => n1938, C2 => n2159
                           , A => n560, ZN => n1682);
   U412 : AOI222_X1 port map( A1 => n53, A2 => n2153, B1 => n181, B2 => n2148, 
                           C1 => n2146, C2 => n561, ZN => n560);
   U413 : OAI221_X1 port map( B1 => n2168, B2 => n583, C1 => n1930, C2 => n2160
                           , A => n584, ZN => n1674);
   U414 : AOI222_X1 port map( A1 => n45, A2 => n2154, B1 => n2149, B2 => n585, 
                           C1 => n2145, C2 => n586, ZN => n584);
   U415 : OAI221_X1 port map( B1 => n2168, B2 => n587, C1 => n1929, C2 => n2160
                           , A => n588, ZN => n1673);
   U416 : AOI222_X1 port map( A1 => n44, A2 => n2154, B1 => n2149, B2 => n589, 
                           C1 => n2145, C2 => n590, ZN => n588);
   U417 : OAI221_X1 port map( B1 => n2168, B2 => n591, C1 => n1928, C2 => n2160
                           , A => n592, ZN => n1672);
   U418 : AOI222_X1 port map( A1 => n43, A2 => n2154, B1 => n2149, B2 => n593, 
                           C1 => n2145, C2 => n594, ZN => n592);
   U419 : OAI221_X1 port map( B1 => n2168, B2 => n595, C1 => n1927, C2 => n2160
                           , A => n596, ZN => n1671);
   U420 : AOI222_X1 port map( A1 => n42, A2 => n2154, B1 => n2149, B2 => n597, 
                           C1 => n2145, C2 => n598, ZN => n596);
   U421 : OAI221_X1 port map( B1 => n2168, B2 => n599, C1 => n1926, C2 => n2160
                           , A => n600, ZN => n1670);
   U422 : AOI222_X1 port map( A1 => n41, A2 => n2154, B1 => n2149, B2 => n601, 
                           C1 => n2145, C2 => n602, ZN => n600);
   U423 : OAI221_X1 port map( B1 => n2168, B2 => n603, C1 => n1925, C2 => n2160
                           , A => n604, ZN => n1669);
   U424 : AOI222_X1 port map( A1 => n40, A2 => n2154, B1 => n2150, B2 => n605, 
                           C1 => n2145, C2 => n606, ZN => n604);
   U425 : OAI221_X1 port map( B1 => n2168, B2 => n607, C1 => n1924, C2 => n2161
                           , A => n608, ZN => n1668);
   U426 : AOI222_X1 port map( A1 => n39, A2 => n2155, B1 => n2150, B2 => n609, 
                           C1 => n2145, C2 => n610, ZN => n608);
   U427 : OAI221_X1 port map( B1 => n2168, B2 => n611, C1 => n1923, C2 => n2161
                           , A => n612, ZN => n1667);
   U428 : AOI222_X1 port map( A1 => n38, A2 => n2155, B1 => n2150, B2 => n613, 
                           C1 => n2145, C2 => n614, ZN => n612);
   U429 : OAI221_X1 port map( B1 => n2168, B2 => n615, C1 => n1922, C2 => n2161
                           , A => n616, ZN => n1666);
   U430 : AOI222_X1 port map( A1 => n37, A2 => n2155, B1 => n2150, B2 => n617, 
                           C1 => n2145, C2 => n618, ZN => n616);
   U431 : OAI22_X1 port map( A1 => n1950, A2 => n2099, B1 => n743, B2 => n2093,
                           ZN => n1501);
   U432 : OAI22_X1 port map( A1 => n1951, A2 => n2099, B1 => n745, B2 => n2093,
                           ZN => n1500);
   U433 : OAI22_X1 port map( A1 => n1952, A2 => n2099, B1 => n747, B2 => n2093,
                           ZN => n1499);
   U434 : OAI22_X1 port map( A1 => n1953, A2 => n2099, B1 => n749, B2 => n2093,
                           ZN => n1498);
   U435 : OAI22_X1 port map( A1 => n1821, A2 => n2087, B1 => n743, B2 => n2081,
                           ZN => n1437);
   U436 : OAI22_X1 port map( A1 => n1820, A2 => n2087, B1 => n745, B2 => n2081,
                           ZN => n1436);
   U437 : OAI22_X1 port map( A1 => n1819, A2 => n2087, B1 => n747, B2 => n2081,
                           ZN => n1435);
   U438 : OAI22_X1 port map( A1 => n1818, A2 => n2087, B1 => n749, B2 => n2081,
                           ZN => n1434);
   U439 : OAI22_X1 port map( A1 => n2010, A2 => n2075, B1 => n743, B2 => n2069,
                           ZN => n1373);
   U440 : OAI22_X1 port map( A1 => n2011, A2 => n2075, B1 => n745, B2 => n2069,
                           ZN => n1372);
   U441 : OAI22_X1 port map( A1 => n2012, A2 => n2075, B1 => n747, B2 => n2069,
                           ZN => n1371);
   U442 : OAI22_X1 port map( A1 => n2013, A2 => n2075, B1 => n749, B2 => n2069,
                           ZN => n1370);
   U443 : OAI22_X1 port map( A1 => n1954, A2 => n2099, B1 => n751, B2 => n2092,
                           ZN => n1497);
   U444 : OAI22_X1 port map( A1 => n1955, A2 => n2098, B1 => n753, B2 => n2092,
                           ZN => n1496);
   U445 : OAI22_X1 port map( A1 => n1956, A2 => n2098, B1 => n755, B2 => n2092,
                           ZN => n1495);
   U446 : OAI22_X1 port map( A1 => n1957, A2 => n2098, B1 => n757, B2 => n2092,
                           ZN => n1494);
   U447 : OAI22_X1 port map( A1 => n1958, A2 => n2098, B1 => n759, B2 => n2092,
                           ZN => n1493);
   U448 : OAI22_X1 port map( A1 => n1959, A2 => n2098, B1 => n761, B2 => n2092,
                           ZN => n1492);
   U449 : OAI22_X1 port map( A1 => n1960, A2 => n2098, B1 => n763, B2 => n2092,
                           ZN => n1491);
   U450 : OAI22_X1 port map( A1 => n1961, A2 => n2098, B1 => n765, B2 => n2092,
                           ZN => n1490);
   U451 : OAI22_X1 port map( A1 => n1962, A2 => n2098, B1 => n767, B2 => n2092,
                           ZN => n1489);
   U452 : OAI22_X1 port map( A1 => n1963, A2 => n2098, B1 => n769, B2 => n2092,
                           ZN => n1488);
   U453 : OAI22_X1 port map( A1 => n1964, A2 => n2098, B1 => n771, B2 => n2092,
                           ZN => n1487);
   U454 : OAI22_X1 port map( A1 => n1965, A2 => n2098, B1 => n773, B2 => n2092,
                           ZN => n1486);
   U455 : OAI22_X1 port map( A1 => n1966, A2 => n2098, B1 => n775, B2 => n2091,
                           ZN => n1485);
   U456 : OAI22_X1 port map( A1 => n1967, A2 => n2097, B1 => n777, B2 => n2091,
                           ZN => n1484);
   U457 : OAI22_X1 port map( A1 => n1968, A2 => n2097, B1 => n779, B2 => n2091,
                           ZN => n1483);
   U458 : OAI22_X1 port map( A1 => n1969, A2 => n2097, B1 => n781, B2 => n2091,
                           ZN => n1482);
   U459 : OAI22_X1 port map( A1 => n1970, A2 => n2097, B1 => n783, B2 => n2091,
                           ZN => n1481);
   U460 : OAI22_X1 port map( A1 => n1971, A2 => n2097, B1 => n785, B2 => n2091,
                           ZN => n1480);
   U461 : OAI22_X1 port map( A1 => n1972, A2 => n2097, B1 => n787, B2 => n2091,
                           ZN => n1479);
   U462 : OAI22_X1 port map( A1 => n1973, A2 => n2097, B1 => n789, B2 => n2091,
                           ZN => n1478);
   U463 : OAI22_X1 port map( A1 => n1974, A2 => n2097, B1 => n791, B2 => n2091,
                           ZN => n1477);
   U464 : OAI22_X1 port map( A1 => n1975, A2 => n2097, B1 => n793, B2 => n2091,
                           ZN => n1476);
   U465 : OAI22_X1 port map( A1 => n1976, A2 => n2097, B1 => n795, B2 => n2091,
                           ZN => n1475);
   U466 : OAI22_X1 port map( A1 => n1977, A2 => n2097, B1 => n797, B2 => n2091,
                           ZN => n1474);
   U467 : OAI22_X1 port map( A1 => n1978, A2 => n2097, B1 => n799, B2 => n2090,
                           ZN => n1473);
   U468 : OAI22_X1 port map( A1 => n1979, A2 => n2096, B1 => n801, B2 => n2090,
                           ZN => n1472);
   U469 : OAI22_X1 port map( A1 => n1980, A2 => n2096, B1 => n803, B2 => n2090,
                           ZN => n1471);
   U470 : OAI22_X1 port map( A1 => n1981, A2 => n2096, B1 => n805, B2 => n2090,
                           ZN => n1470);
   U471 : OAI22_X1 port map( A1 => n1982, A2 => n2096, B1 => n807, B2 => n2090,
                           ZN => n1469);
   U472 : OAI22_X1 port map( A1 => n1983, A2 => n2096, B1 => n809, B2 => n2090,
                           ZN => n1468);
   U473 : OAI22_X1 port map( A1 => n1984, A2 => n2096, B1 => n811, B2 => n2090,
                           ZN => n1467);
   U474 : OAI22_X1 port map( A1 => n1985, A2 => n2096, B1 => n813, B2 => n2090,
                           ZN => n1466);
   U475 : OAI22_X1 port map( A1 => n1986, A2 => n2096, B1 => n815, B2 => n2090,
                           ZN => n1465);
   U476 : OAI22_X1 port map( A1 => n1987, A2 => n2096, B1 => n817, B2 => n2090,
                           ZN => n1464);
   U477 : OAI22_X1 port map( A1 => n1988, A2 => n2096, B1 => n819, B2 => n2090,
                           ZN => n1463);
   U478 : OAI22_X1 port map( A1 => n1989, A2 => n2096, B1 => n821, B2 => n2090,
                           ZN => n1462);
   U479 : OAI22_X1 port map( A1 => n1990, A2 => n2096, B1 => n823, B2 => n2089,
                           ZN => n1461);
   U480 : OAI22_X1 port map( A1 => n1991, A2 => n2095, B1 => n825, B2 => n2089,
                           ZN => n1460);
   U481 : OAI22_X1 port map( A1 => n1992, A2 => n2095, B1 => n827, B2 => n2089,
                           ZN => n1459);
   U482 : OAI22_X1 port map( A1 => n1993, A2 => n2095, B1 => n829, B2 => n2089,
                           ZN => n1458);
   U483 : OAI22_X1 port map( A1 => n1994, A2 => n2095, B1 => n831, B2 => n2089,
                           ZN => n1457);
   U484 : OAI22_X1 port map( A1 => n1995, A2 => n2095, B1 => n833, B2 => n2089,
                           ZN => n1456);
   U485 : OAI22_X1 port map( A1 => n1996, A2 => n2095, B1 => n835, B2 => n2089,
                           ZN => n1455);
   U486 : OAI22_X1 port map( A1 => n1997, A2 => n2095, B1 => n837, B2 => n2089,
                           ZN => n1454);
   U487 : OAI22_X1 port map( A1 => n1998, A2 => n2095, B1 => n839, B2 => n2089,
                           ZN => n1453);
   U488 : OAI22_X1 port map( A1 => n1999, A2 => n2095, B1 => n841, B2 => n2089,
                           ZN => n1452);
   U489 : OAI22_X1 port map( A1 => n2000, A2 => n2095, B1 => n843, B2 => n2089,
                           ZN => n1451);
   U490 : OAI22_X1 port map( A1 => n2001, A2 => n2095, B1 => n845, B2 => n2089,
                           ZN => n1450);
   U491 : OAI22_X1 port map( A1 => n1204, A2 => n2095, B1 => n847, B2 => n2088,
                           ZN => n1449);
   U492 : OAI22_X1 port map( A1 => n1202, A2 => n2094, B1 => n849, B2 => n2088,
                           ZN => n1448);
   U493 : OAI22_X1 port map( A1 => n1200, A2 => n2094, B1 => n851, B2 => n2088,
                           ZN => n1447);
   U494 : OAI22_X1 port map( A1 => n2002, A2 => n2094, B1 => n853, B2 => n2088,
                           ZN => n1446);
   U495 : OAI22_X1 port map( A1 => n2003, A2 => n2094, B1 => n855, B2 => n2088,
                           ZN => n1445);
   U496 : OAI22_X1 port map( A1 => n2004, A2 => n2094, B1 => n857, B2 => n2088,
                           ZN => n1444);
   U497 : OAI22_X1 port map( A1 => n2005, A2 => n2094, B1 => n859, B2 => n2088,
                           ZN => n1443);
   U498 : OAI22_X1 port map( A1 => n2006, A2 => n2094, B1 => n861, B2 => n2088,
                           ZN => n1442);
   U499 : OAI22_X1 port map( A1 => n2007, A2 => n2094, B1 => n863, B2 => n2088,
                           ZN => n1441);
   U500 : OAI22_X1 port map( A1 => n2008, A2 => n2094, B1 => n865, B2 => n2088,
                           ZN => n1440);
   U501 : OAI22_X1 port map( A1 => n2009, A2 => n2094, B1 => n867, B2 => n2088,
                           ZN => n1439);
   U502 : OAI22_X1 port map( A1 => n415, A2 => n2094, B1 => n871, B2 => n2088, 
                           ZN => n1438);
   U503 : OAI22_X1 port map( A1 => n1817, A2 => n2087, B1 => n751, B2 => n2080,
                           ZN => n1433);
   U504 : OAI22_X1 port map( A1 => n1816, A2 => n2086, B1 => n753, B2 => n2080,
                           ZN => n1432);
   U505 : OAI22_X1 port map( A1 => n1815, A2 => n2086, B1 => n755, B2 => n2080,
                           ZN => n1431);
   U506 : OAI22_X1 port map( A1 => n1814, A2 => n2086, B1 => n757, B2 => n2080,
                           ZN => n1430);
   U507 : OAI22_X1 port map( A1 => n1813, A2 => n2086, B1 => n759, B2 => n2080,
                           ZN => n1429);
   U508 : OAI22_X1 port map( A1 => n1812, A2 => n2086, B1 => n761, B2 => n2080,
                           ZN => n1428);
   U509 : OAI22_X1 port map( A1 => n1811, A2 => n2086, B1 => n763, B2 => n2080,
                           ZN => n1427);
   U510 : OAI22_X1 port map( A1 => n1810, A2 => n2086, B1 => n765, B2 => n2080,
                           ZN => n1426);
   U511 : OAI22_X1 port map( A1 => n1809, A2 => n2086, B1 => n767, B2 => n2080,
                           ZN => n1425);
   U512 : OAI22_X1 port map( A1 => n1808, A2 => n2086, B1 => n769, B2 => n2080,
                           ZN => n1424);
   U513 : OAI22_X1 port map( A1 => n1807, A2 => n2086, B1 => n771, B2 => n2080,
                           ZN => n1423);
   U514 : OAI22_X1 port map( A1 => n1806, A2 => n2086, B1 => n773, B2 => n2080,
                           ZN => n1422);
   U515 : OAI22_X1 port map( A1 => n1805, A2 => n2086, B1 => n775, B2 => n2079,
                           ZN => n1421);
   U516 : OAI22_X1 port map( A1 => n1804, A2 => n2085, B1 => n777, B2 => n2079,
                           ZN => n1420);
   U517 : OAI22_X1 port map( A1 => n1803, A2 => n2085, B1 => n779, B2 => n2079,
                           ZN => n1419);
   U518 : OAI22_X1 port map( A1 => n1802, A2 => n2085, B1 => n781, B2 => n2079,
                           ZN => n1418);
   U519 : OAI22_X1 port map( A1 => n1801, A2 => n2085, B1 => n783, B2 => n2079,
                           ZN => n1417);
   U520 : OAI22_X1 port map( A1 => n1800, A2 => n2085, B1 => n785, B2 => n2079,
                           ZN => n1416);
   U521 : OAI22_X1 port map( A1 => n1799, A2 => n2085, B1 => n787, B2 => n2079,
                           ZN => n1415);
   U522 : OAI22_X1 port map( A1 => n1798, A2 => n2085, B1 => n789, B2 => n2079,
                           ZN => n1414);
   U523 : OAI22_X1 port map( A1 => n1797, A2 => n2085, B1 => n791, B2 => n2079,
                           ZN => n1413);
   U524 : OAI22_X1 port map( A1 => n1796, A2 => n2085, B1 => n793, B2 => n2079,
                           ZN => n1412);
   U525 : OAI22_X1 port map( A1 => n1795, A2 => n2085, B1 => n795, B2 => n2079,
                           ZN => n1411);
   U526 : OAI22_X1 port map( A1 => n1794, A2 => n2085, B1 => n797, B2 => n2079,
                           ZN => n1410);
   U527 : OAI22_X1 port map( A1 => n1793, A2 => n2085, B1 => n799, B2 => n2078,
                           ZN => n1409);
   U528 : OAI22_X1 port map( A1 => n2029, A2 => n2084, B1 => n801, B2 => n2078,
                           ZN => n1408);
   U529 : OAI22_X1 port map( A1 => n2030, A2 => n2084, B1 => n803, B2 => n2078,
                           ZN => n1407);
   U530 : OAI22_X1 port map( A1 => n2031, A2 => n2084, B1 => n805, B2 => n2078,
                           ZN => n1406);
   U531 : OAI22_X1 port map( A1 => n2032, A2 => n2084, B1 => n807, B2 => n2078,
                           ZN => n1405);
   U532 : OAI22_X1 port map( A1 => n2033, A2 => n2084, B1 => n809, B2 => n2078,
                           ZN => n1404);
   U533 : OAI22_X1 port map( A1 => n2034, A2 => n2084, B1 => n811, B2 => n2078,
                           ZN => n1403);
   U534 : OAI22_X1 port map( A1 => n2035, A2 => n2084, B1 => n813, B2 => n2078,
                           ZN => n1402);
   U535 : OAI22_X1 port map( A1 => n2036, A2 => n2084, B1 => n815, B2 => n2078,
                           ZN => n1401);
   U536 : OAI22_X1 port map( A1 => n2037, A2 => n2084, B1 => n817, B2 => n2078,
                           ZN => n1400);
   U537 : OAI22_X1 port map( A1 => n2038, A2 => n2084, B1 => n819, B2 => n2078,
                           ZN => n1399);
   U538 : OAI22_X1 port map( A1 => n2039, A2 => n2084, B1 => n821, B2 => n2078,
                           ZN => n1398);
   U539 : OAI22_X1 port map( A1 => n2040, A2 => n2084, B1 => n823, B2 => n2077,
                           ZN => n1397);
   U540 : OAI22_X1 port map( A1 => n2041, A2 => n2083, B1 => n825, B2 => n2077,
                           ZN => n1396);
   U541 : OAI22_X1 port map( A1 => n2042, A2 => n2083, B1 => n827, B2 => n2077,
                           ZN => n1395);
   U542 : OAI22_X1 port map( A1 => n2043, A2 => n2083, B1 => n829, B2 => n2077,
                           ZN => n1394);
   U543 : OAI22_X1 port map( A1 => n2044, A2 => n2083, B1 => n831, B2 => n2077,
                           ZN => n1393);
   U544 : OAI22_X1 port map( A1 => n2045, A2 => n2083, B1 => n833, B2 => n2077,
                           ZN => n1392);
   U545 : OAI22_X1 port map( A1 => n2046, A2 => n2083, B1 => n835, B2 => n2077,
                           ZN => n1391);
   U546 : OAI22_X1 port map( A1 => n2047, A2 => n2083, B1 => n837, B2 => n2077,
                           ZN => n1390);
   U547 : OAI22_X1 port map( A1 => n2048, A2 => n2083, B1 => n839, B2 => n2077,
                           ZN => n1389);
   U548 : OAI22_X1 port map( A1 => n2049, A2 => n2083, B1 => n841, B2 => n2077,
                           ZN => n1388);
   U549 : OAI22_X1 port map( A1 => n2050, A2 => n2083, B1 => n843, B2 => n2077,
                           ZN => n1387);
   U550 : OAI22_X1 port map( A1 => n2051, A2 => n2083, B1 => n845, B2 => n2077,
                           ZN => n1386);
   U551 : OAI22_X1 port map( A1 => n2052, A2 => n2083, B1 => n847, B2 => n2076,
                           ZN => n1385);
   U552 : OAI22_X1 port map( A1 => n2053, A2 => n2082, B1 => n849, B2 => n2076,
                           ZN => n1384);
   U553 : OAI22_X1 port map( A1 => n2054, A2 => n2082, B1 => n851, B2 => n2076,
                           ZN => n1383);
   U554 : OAI22_X1 port map( A1 => n2055, A2 => n2082, B1 => n853, B2 => n2076,
                           ZN => n1382);
   U555 : OAI22_X1 port map( A1 => n2056, A2 => n2082, B1 => n855, B2 => n2076,
                           ZN => n1381);
   U556 : OAI22_X1 port map( A1 => n2057, A2 => n2082, B1 => n857, B2 => n2076,
                           ZN => n1380);
   U557 : OAI22_X1 port map( A1 => n2058, A2 => n2082, B1 => n859, B2 => n2076,
                           ZN => n1379);
   U558 : OAI22_X1 port map( A1 => n2059, A2 => n2082, B1 => n861, B2 => n2076,
                           ZN => n1378);
   U559 : OAI22_X1 port map( A1 => n2060, A2 => n2082, B1 => n863, B2 => n2076,
                           ZN => n1377);
   U560 : OAI22_X1 port map( A1 => n2061, A2 => n2082, B1 => n865, B2 => n2076,
                           ZN => n1376);
   U561 : OAI22_X1 port map( A1 => n2062, A2 => n2082, B1 => n867, B2 => n2076,
                           ZN => n1375);
   U562 : OAI22_X1 port map( A1 => n2063, A2 => n2082, B1 => n871, B2 => n2076,
                           ZN => n1374);
   U563 : OAI22_X1 port map( A1 => n2014, A2 => n2075, B1 => n751, B2 => n2068,
                           ZN => n1369);
   U564 : OAI22_X1 port map( A1 => n2015, A2 => n2074, B1 => n753, B2 => n2068,
                           ZN => n1368);
   U565 : OAI22_X1 port map( A1 => n2016, A2 => n2074, B1 => n755, B2 => n2068,
                           ZN => n1367);
   U566 : OAI22_X1 port map( A1 => n2017, A2 => n2074, B1 => n757, B2 => n2068,
                           ZN => n1366);
   U567 : OAI22_X1 port map( A1 => n2018, A2 => n2074, B1 => n759, B2 => n2068,
                           ZN => n1365);
   U568 : OAI22_X1 port map( A1 => n2019, A2 => n2074, B1 => n761, B2 => n2068,
                           ZN => n1364);
   U569 : OAI22_X1 port map( A1 => n2020, A2 => n2074, B1 => n763, B2 => n2068,
                           ZN => n1363);
   U570 : OAI22_X1 port map( A1 => n2021, A2 => n2074, B1 => n765, B2 => n2068,
                           ZN => n1362);
   U571 : OAI22_X1 port map( A1 => n2022, A2 => n2074, B1 => n767, B2 => n2068,
                           ZN => n1361);
   U572 : OAI22_X1 port map( A1 => n2023, A2 => n2074, B1 => n769, B2 => n2068,
                           ZN => n1360);
   U573 : OAI22_X1 port map( A1 => n2024, A2 => n2074, B1 => n771, B2 => n2068,
                           ZN => n1359);
   U574 : OAI22_X1 port map( A1 => n2025, A2 => n2074, B1 => n773, B2 => n2068,
                           ZN => n1358);
   U575 : OAI22_X1 port map( A1 => n2026, A2 => n2074, B1 => n775, B2 => n2067,
                           ZN => n1357);
   U576 : OAI22_X1 port map( A1 => n2027, A2 => n2073, B1 => n777, B2 => n2067,
                           ZN => n1356);
   U577 : OAI22_X1 port map( A1 => n2028, A2 => n2073, B1 => n779, B2 => n2067,
                           ZN => n1355);
   U578 : OAI22_X1 port map( A1 => n1738, A2 => n2073, B1 => n781, B2 => n2067,
                           ZN => n1354);
   U579 : OAI22_X1 port map( A1 => n1737, A2 => n2073, B1 => n783, B2 => n2067,
                           ZN => n1353);
   U580 : OAI22_X1 port map( A1 => n1736, A2 => n2073, B1 => n785, B2 => n2067,
                           ZN => n1352);
   U581 : OAI22_X1 port map( A1 => n1735, A2 => n2073, B1 => n787, B2 => n2067,
                           ZN => n1351);
   U582 : OAI22_X1 port map( A1 => n1734, A2 => n2073, B1 => n789, B2 => n2067,
                           ZN => n1350);
   U583 : OAI22_X1 port map( A1 => n1733, A2 => n2073, B1 => n791, B2 => n2067,
                           ZN => n1349);
   U584 : OAI22_X1 port map( A1 => n1732, A2 => n2073, B1 => n793, B2 => n2067,
                           ZN => n1348);
   U585 : OAI22_X1 port map( A1 => n1731, A2 => n2073, B1 => n795, B2 => n2067,
                           ZN => n1347);
   U586 : OAI22_X1 port map( A1 => n1730, A2 => n2073, B1 => n797, B2 => n2067,
                           ZN => n1346);
   U587 : OAI22_X1 port map( A1 => n1729, A2 => n2073, B1 => n799, B2 => n2066,
                           ZN => n1345);
   U588 : OAI22_X1 port map( A1 => n1728, A2 => n2072, B1 => n801, B2 => n2066,
                           ZN => n1344);
   U589 : OAI22_X1 port map( A1 => n1727, A2 => n2072, B1 => n803, B2 => n2066,
                           ZN => n1343);
   U590 : OAI22_X1 port map( A1 => n1726, A2 => n2072, B1 => n805, B2 => n2066,
                           ZN => n1342);
   U591 : OAI22_X1 port map( A1 => n1725, A2 => n2072, B1 => n807, B2 => n2066,
                           ZN => n1341);
   U592 : OAI22_X1 port map( A1 => n1724, A2 => n2072, B1 => n809, B2 => n2066,
                           ZN => n1340);
   U593 : OAI22_X1 port map( A1 => n1723, A2 => n2072, B1 => n811, B2 => n2066,
                           ZN => n1339);
   U594 : OAI22_X1 port map( A1 => n1722, A2 => n2072, B1 => n813, B2 => n2066,
                           ZN => n1338);
   U595 : OAI22_X1 port map( A1 => n1721, A2 => n2072, B1 => n815, B2 => n2066,
                           ZN => n1337);
   U596 : OAI22_X1 port map( A1 => n1720, A2 => n2072, B1 => n817, B2 => n2066,
                           ZN => n1336);
   U597 : OAI22_X1 port map( A1 => n1719, A2 => n2072, B1 => n819, B2 => n2066,
                           ZN => n1335);
   U598 : OAI22_X1 port map( A1 => n1718, A2 => n2072, B1 => n821, B2 => n2066,
                           ZN => n1334);
   U599 : OAI22_X1 port map( A1 => n1717, A2 => n2072, B1 => n823, B2 => n2065,
                           ZN => n1333);
   U600 : OAI22_X1 port map( A1 => n1716, A2 => n2071, B1 => n825, B2 => n2065,
                           ZN => n1332);
   U601 : OAI22_X1 port map( A1 => n1715, A2 => n2071, B1 => n827, B2 => n2065,
                           ZN => n1331);
   U602 : OAI22_X1 port map( A1 => n1714, A2 => n2071, B1 => n829, B2 => n2065,
                           ZN => n1330);
   U603 : OAI22_X1 port map( A1 => n1713, A2 => n2071, B1 => n831, B2 => n2065,
                           ZN => n1329);
   U604 : OAI22_X1 port map( A1 => n1712, A2 => n2071, B1 => n833, B2 => n2065,
                           ZN => n1328);
   U605 : OAI22_X1 port map( A1 => n1711, A2 => n2071, B1 => n835, B2 => n2065,
                           ZN => n1327);
   U606 : OAI22_X1 port map( A1 => n1710, A2 => n2071, B1 => n837, B2 => n2065,
                           ZN => n1326);
   U607 : OAI22_X1 port map( A1 => n1709, A2 => n2071, B1 => n839, B2 => n2065,
                           ZN => n1325);
   U608 : OAI22_X1 port map( A1 => n1708, A2 => n2071, B1 => n841, B2 => n2065,
                           ZN => n1324);
   U609 : OAI22_X1 port map( A1 => n1707, A2 => n2071, B1 => n843, B2 => n2065,
                           ZN => n1323);
   U610 : OAI22_X1 port map( A1 => n1706, A2 => n2071, B1 => n845, B2 => n2065,
                           ZN => n1322);
   U611 : OAI22_X1 port map( A1 => n1705, A2 => n2071, B1 => n847, B2 => n2064,
                           ZN => n1321);
   U612 : OAI22_X1 port map( A1 => n1704, A2 => n2070, B1 => n849, B2 => n2064,
                           ZN => n1320);
   U613 : OAI22_X1 port map( A1 => n1703, A2 => n2070, B1 => n851, B2 => n2064,
                           ZN => n1319);
   U614 : OAI22_X1 port map( A1 => n1702, A2 => n2070, B1 => n853, B2 => n2064,
                           ZN => n1318);
   U615 : OAI22_X1 port map( A1 => n1701, A2 => n2070, B1 => n855, B2 => n2064,
                           ZN => n1317);
   U616 : OAI22_X1 port map( A1 => n1700, A2 => n2070, B1 => n857, B2 => n2064,
                           ZN => n1316);
   U617 : OAI22_X1 port map( A1 => n1699, A2 => n2070, B1 => n859, B2 => n2064,
                           ZN => n1315);
   U618 : OAI22_X1 port map( A1 => n1698, A2 => n2070, B1 => n861, B2 => n2064,
                           ZN => n1314);
   U619 : OAI22_X1 port map( A1 => n1697, A2 => n2070, B1 => n863, B2 => n2064,
                           ZN => n1313);
   U620 : OAI22_X1 port map( A1 => n1696, A2 => n2070, B1 => n865, B2 => n2064,
                           ZN => n1312);
   U621 : OAI22_X1 port map( A1 => n1695, A2 => n2070, B1 => n867, B2 => n2064,
                           ZN => n1311);
   U622 : OAI22_X1 port map( A1 => n1694, A2 => n2070, B1 => n871, B2 => n2064,
                           ZN => n1310);
   U623 : INV_X1 port map( A => DATAIN(0), ZN => n743);
   U624 : INV_X1 port map( A => DATAIN(1), ZN => n745);
   U625 : INV_X1 port map( A => DATAIN(2), ZN => n747);
   U626 : INV_X1 port map( A => DATAIN(3), ZN => n749);
   U627 : INV_X1 port map( A => DATAIN(4), ZN => n751);
   U628 : INV_X1 port map( A => DATAIN(5), ZN => n753);
   U629 : INV_X1 port map( A => DATAIN(6), ZN => n755);
   U630 : INV_X1 port map( A => DATAIN(7), ZN => n757);
   U631 : INV_X1 port map( A => DATAIN(8), ZN => n759);
   U632 : INV_X1 port map( A => DATAIN(9), ZN => n761);
   U633 : INV_X1 port map( A => DATAIN(10), ZN => n763);
   U634 : INV_X1 port map( A => DATAIN(11), ZN => n765);
   U635 : INV_X1 port map( A => DATAIN(12), ZN => n767);
   U636 : INV_X1 port map( A => DATAIN(13), ZN => n769);
   U637 : INV_X1 port map( A => DATAIN(14), ZN => n771);
   U638 : INV_X1 port map( A => DATAIN(15), ZN => n773);
   U639 : INV_X1 port map( A => DATAIN(16), ZN => n775);
   U640 : INV_X1 port map( A => DATAIN(17), ZN => n777);
   U641 : INV_X1 port map( A => DATAIN(18), ZN => n779);
   U642 : INV_X1 port map( A => DATAIN(19), ZN => n781);
   U643 : INV_X1 port map( A => DATAIN(20), ZN => n783);
   U644 : INV_X1 port map( A => DATAIN(21), ZN => n785);
   U645 : INV_X1 port map( A => DATAIN(22), ZN => n787);
   U646 : INV_X1 port map( A => DATAIN(23), ZN => n789);
   U647 : INV_X1 port map( A => DATAIN(24), ZN => n791);
   U648 : INV_X1 port map( A => DATAIN(25), ZN => n793);
   U649 : INV_X1 port map( A => DATAIN(26), ZN => n795);
   U650 : INV_X1 port map( A => DATAIN(27), ZN => n797);
   U651 : INV_X1 port map( A => DATAIN(28), ZN => n799);
   U652 : INV_X1 port map( A => DATAIN(29), ZN => n801);
   U653 : INV_X1 port map( A => DATAIN(30), ZN => n803);
   U654 : INV_X1 port map( A => DATAIN(31), ZN => n805);
   U655 : INV_X1 port map( A => DATAIN(32), ZN => n807);
   U656 : INV_X1 port map( A => DATAIN(33), ZN => n809);
   U657 : INV_X1 port map( A => DATAIN(34), ZN => n811);
   U658 : INV_X1 port map( A => DATAIN(35), ZN => n813);
   U659 : INV_X1 port map( A => DATAIN(36), ZN => n815);
   U660 : INV_X1 port map( A => DATAIN(37), ZN => n817);
   U661 : INV_X1 port map( A => DATAIN(38), ZN => n819);
   U662 : INV_X1 port map( A => DATAIN(39), ZN => n821);
   U663 : INV_X1 port map( A => DATAIN(40), ZN => n823);
   U664 : INV_X1 port map( A => DATAIN(41), ZN => n825);
   U665 : INV_X1 port map( A => DATAIN(42), ZN => n827);
   U666 : INV_X1 port map( A => DATAIN(43), ZN => n829);
   U667 : INV_X1 port map( A => DATAIN(44), ZN => n831);
   U668 : INV_X1 port map( A => DATAIN(45), ZN => n833);
   U669 : INV_X1 port map( A => DATAIN(46), ZN => n835);
   U670 : INV_X1 port map( A => DATAIN(47), ZN => n837);
   U671 : INV_X1 port map( A => DATAIN(48), ZN => n839);
   U672 : INV_X1 port map( A => DATAIN(49), ZN => n841);
   U673 : INV_X1 port map( A => DATAIN(50), ZN => n843);
   U674 : INV_X1 port map( A => DATAIN(51), ZN => n845);
   U675 : INV_X1 port map( A => DATAIN(52), ZN => n847);
   U676 : INV_X1 port map( A => DATAIN(53), ZN => n849);
   U677 : INV_X1 port map( A => DATAIN(54), ZN => n851);
   U678 : INV_X1 port map( A => DATAIN(55), ZN => n853);
   U679 : INV_X1 port map( A => DATAIN(56), ZN => n855);
   U680 : INV_X1 port map( A => DATAIN(57), ZN => n857);
   U681 : INV_X1 port map( A => DATAIN(58), ZN => n859);
   U682 : INV_X1 port map( A => DATAIN(59), ZN => n861);
   U683 : INV_X1 port map( A => DATAIN(60), ZN => n863);
   U684 : INV_X1 port map( A => DATAIN(61), ZN => n865);
   U685 : INV_X1 port map( A => DATAIN(62), ZN => n867);
   U686 : INV_X1 port map( A => DATAIN(63), ZN => n871);
   U687 : CLKBUF_X1 port map( A => n979, Z => n2069);
   U688 : CLKBUF_X1 port map( A => n978, Z => n2075);
   U689 : CLKBUF_X1 port map( A => n939, Z => n2081);
   U690 : CLKBUF_X1 port map( A => n938, Z => n2087);
   U691 : CLKBUF_X1 port map( A => n876, Z => n2093);
   U692 : CLKBUF_X1 port map( A => n875, Z => n2099);
   U693 : CLKBUF_X1 port map( A => n742, Z => n2105);
   U694 : CLKBUF_X1 port map( A => n741, Z => n2111);
   U695 : CLKBUF_X1 port map( A => n740, Z => n2117);
   U696 : CLKBUF_X1 port map( A => n739, Z => n2123);
   U697 : CLKBUF_X1 port map( A => n738, Z => n2129);
   U698 : CLKBUF_X1 port map( A => n736, Z => n2135);
   U699 : CLKBUF_X1 port map( A => n735, Z => n2141);
   U700 : CLKBUF_X1 port map( A => n527, Z => n2147);
   U701 : CLKBUF_X1 port map( A => n525, Z => n2158);
   U702 : CLKBUF_X1 port map( A => n523, Z => n2164);
   U703 : CLKBUF_X1 port map( A => n521, Z => n2170);
   U704 : INV_X1 port map( A => ADD_RD2(0), ZN => n2171);
   U705 : INV_X1 port map( A => ADD_RD2(1), ZN => n2172);
   U706 : INV_X1 port map( A => ADD_RD1(0), ZN => n2173);
   U707 : INV_X1 port map( A => ADD_RD1(1), ZN => n2174);
   U708 : INV_X1 port map( A => ADD_WR(0), ZN => n2175);
   U709 : INV_X1 port map( A => ADD_WR(1), ZN => n2176);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4.all;

entity register_file_reg_size64_file_size4_6 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_reg_size64_file_size4_6;

architecture SYN_BEHAVIORAL of register_file_reg_size64_file_size4_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n415, n1200, n1202, n1204, n1310, n1311, n1312, n1313, n1314, n1315
      , n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n871, n872, 
      n873, n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, 
      n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, 
      n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, 
      n909, n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, 
      n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, 
      n933, n934, n935, n936, n938, n939, n940, n941, n942, n943, n944, n945, 
      n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, 
      n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, 
      n970, n971, n972, n973, n974, n975, n977, n978, n979, n980, n981, n982, 
      n983, n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, 
      n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, 
      n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, 
      n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, 
      n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, 
      n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, 
      n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, 
      n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1950, n1951, n1952, 
      n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, 
      n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, 
      n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, 
      n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, 
      n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, 
      n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, 
      n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, 
      n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, 
      n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, 
      n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, 
      n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062 : 
      std_logic;

begin
   
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => n174,
                           QN => n997);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => n175,
                           QN => n996);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => n176,
                           QN => n995);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => n177,
                           QN => n994);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => n178,
                           QN => n993);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => n179,
                           QN => n992);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => n180,
                           QN => n991);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => n181,
                           QN => n990);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => n182,
                           QN => n989);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => n183, 
                           QN => n988);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => n184, 
                           QN => n987);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => n185, 
                           QN => n986);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => n186, 
                           QN => n985);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => n187, 
                           QN => n984);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => n188, 
                           QN => n983);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => n189, 
                           QN => n982);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => n190, 
                           QN => n981);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => n191, 
                           QN => n980);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => n192, 
                           QN => n977);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => n65, 
                           QN => n974);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => n66, 
                           QN => n973);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n67, 
                           QN => n972);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => n68, 
                           QN => n971);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => n69, 
                           QN => n970);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => n70, 
                           QN => n969);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => n71, 
                           QN => n968);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => n72, 
                           QN => n967);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => n73, 
                           QN => n966);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => n74, 
                           QN => n965);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => n75, 
                           QN => n964);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => n76, 
                           QN => n963);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => n77, 
                           QN => n962);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => n78, 
                           QN => n961);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => n79, 
                           QN => n960);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => n80, 
                           QN => n959);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => n81, 
                           QN => n958);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => n82, 
                           QN => n957);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => n83, 
                           QN => n956);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => n84, 
                           QN => n955);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => n85, 
                           QN => n954);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => n86, 
                           QN => n953);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => n87, 
                           QN => n952);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => n88, 
                           QN => n951);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => n89, 
                           QN => n950);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => n90, 
                           QN => n949);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => n91, 
                           QN => n948);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => n92, 
                           QN => n947);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => n93, 
                           QN => n946);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => n94, 
                           QN => n945);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => n95, 
                           QN => n944);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => n96, 
                           QN => n943);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => n97, 
                           QN => n942);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => n98, 
                           QN => n941);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => n99, 
                           QN => n940);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => n2, 
                           QN => n935);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => n3, 
                           QN => n934);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => n4, 
                           QN => n933);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => n5, 
                           QN => n932);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => n6, 
                           QN => n931);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => n7, 
                           QN => n930);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => n8, 
                           QN => n929);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => n9, 
                           QN => n928);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => n13, 
                           QN => n927);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => n14, 
                           QN => n926);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => n15, 
                           QN => n925);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => n16, 
                           QN => n924);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => n17, 
                           QN => n923);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => n18, 
                           QN => n922);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => n19, 
                           QN => n921);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => n20, 
                           QN => n920);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => n21, 
                           QN => n919);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => n22, 
                           QN => n918);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => n23, 
                           QN => n917);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => n24, 
                           QN => n916);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => n25, 
                           QN => n915);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => n26, 
                           QN => n914);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n27, 
                           QN => n913);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => n28, 
                           QN => n912);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n29, 
                           QN => n911);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => n30, 
                           QN => n910);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n31, 
                           QN => n909);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => n32, 
                           QN => n908);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n33, 
                           QN => n907);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => n34, 
                           QN => n906);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n35, 
                           QN => n905);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => n36, 
                           QN => n904);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => n37, 
                           QN => n903);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => n38, 
                           QN => n902);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => n39, 
                           QN => n901);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => n40, 
                           QN => n900);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => n41, 
                           QN => n899);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => n42, 
                           QN => n898);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => n43, 
                           QN => n897);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => n44, 
                           QN => n896);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => n45, 
                           QN => n895);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => n46, 
                           QN => n894);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => n47, 
                           QN => n893);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => n48, 
                           QN => n892);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => n49, 
                           QN => n891);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => n50, 
                           QN => n890);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => n51, 
                           QN => n889);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => n52, 
                           QN => n888);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => n53, 
                           QN => n887);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => n54, 
                           QN => n886);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n55, 
                           QN => n885);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => n56, 
                           QN => n884);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n57, 
                           QN => n883);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => n58, 
                           QN => n882);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n59, 
                           QN => n881);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => n60, 
                           QN => n880);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n61, 
                           QN => n879);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => n62, 
                           QN => n878);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n63, 
                           QN => n877);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => n64, 
                           QN => n874);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n999,
                           QN => n728);
   OUT2_reg_63_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => OUT2(63), QN
                           => n1822);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n1000
                           , QN => n725);
   OUT2_reg_62_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => OUT2(62), QN
                           => n1823);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n1001
                           , QN => n722);
   OUT2_reg_61_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => OUT2(61), QN
                           => n1824);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n1002
                           , QN => n719);
   OUT2_reg_60_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => OUT2(60), QN
                           => n1825);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n1003
                           , QN => n716);
   OUT2_reg_59_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => OUT2(59), QN
                           => n1826);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n1004
                           , QN => n713);
   OUT2_reg_58_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => OUT2(58), QN
                           => n1827);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n1005
                           , QN => n710);
   OUT2_reg_57_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => OUT2(57), QN
                           => n1828);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n1006
                           , QN => n707);
   OUT2_reg_56_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => OUT2(56), QN
                           => n1829);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n1007
                           , QN => n704);
   OUT2_reg_55_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => OUT2(55), QN
                           => n1830);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n1008
                           , QN => n700);
   OUT2_reg_54_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => OUT2(54), QN
                           => n1831);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n1009
                           , QN => n696);
   OUT2_reg_53_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => OUT2(53), QN
                           => n1832);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n1010
                           , QN => n692);
   OUT2_reg_52_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => OUT2(52), QN
                           => n1833);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n1011
                           , QN => n689);
   OUT2_reg_51_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => OUT2(51), QN
                           => n1834);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n1012
                           , QN => n686);
   OUT2_reg_50_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => OUT2(50), QN
                           => n1835);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n1013
                           , QN => n683);
   OUT2_reg_49_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => OUT2(49), QN
                           => n1836);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n1014
                           , QN => n680);
   OUT2_reg_48_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => OUT2(48), QN
                           => n1837);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n1015
                           , QN => n677);
   OUT2_reg_47_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => OUT2(47), QN
                           => n1838);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n1016
                           , QN => n674);
   OUT2_reg_46_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => OUT2(46), QN
                           => n1839);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n1017
                           , QN => n671);
   OUT2_reg_45_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => OUT2(45), QN
                           => n1840);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n1018
                           , QN => n668);
   OUT2_reg_44_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => OUT2(44), QN
                           => n1841);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n1019
                           , QN => n665);
   OUT2_reg_43_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => OUT2(43), QN
                           => n1842);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n1020
                           , QN => n662);
   OUT2_reg_42_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => OUT2(42), QN
                           => n1843);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n1021
                           , QN => n659);
   OUT2_reg_41_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => OUT2(41), QN
                           => n1844);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n1022
                           , QN => n656);
   OUT2_reg_40_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => OUT2(40), QN
                           => n1845);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n1023
                           , QN => n653);
   OUT2_reg_39_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => OUT2(39), QN
                           => n1846);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n1024
                           , QN => n650);
   OUT2_reg_38_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => OUT2(38), QN
                           => n1847);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n1025
                           , QN => n647);
   OUT2_reg_37_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => OUT2(37), QN
                           => n1848);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n1026
                           , QN => n644);
   OUT2_reg_36_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => OUT2(36), QN
                           => n1849);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n1027
                           , QN => n641);
   OUT2_reg_35_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => OUT2(35), QN
                           => n1850);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n1028
                           , QN => n638);
   OUT2_reg_34_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => OUT2(34), QN
                           => n1851);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n1029
                           , QN => n635);
   OUT2_reg_33_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => OUT2(33), QN
                           => n1852);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n1030
                           , QN => n632);
   OUT2_reg_32_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => OUT2(32), QN
                           => n1853);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n1031
                           , QN => n629);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => OUT2(31), QN
                           => n1854);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n1032
                           , QN => n626);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => OUT2(30), QN
                           => n1855);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n1033
                           , QN => n623);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => OUT2(29), QN
                           => n1856);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n1034
                           , QN => n619);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => OUT2(28), QN
                           => n1857);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n1035
                           , QN => n615);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => OUT2(27), QN
                           => n1858);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n1036
                           , QN => n611);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => OUT2(26), QN
                           => n1859);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n1037
                           , QN => n607);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => OUT2(25), QN
                           => n1860);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n1038
                           , QN => n603);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => OUT2(24), QN
                           => n1861);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n1039
                           , QN => n599);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => OUT2(23), QN
                           => n1862);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n1040
                           , QN => n595);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => OUT2(22), QN
                           => n1863);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n1041
                           , QN => n591);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => OUT2(21), QN
                           => n1864);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n1042
                           , QN => n587);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => OUT2(20), QN
                           => n1865);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n1043
                           , QN => n583);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => OUT2(19), QN
                           => n1866);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n1044
                           , QN => n580);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => OUT2(18), QN
                           => n1867);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n1045
                           , QN => n577);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => OUT2(17), QN
                           => n1868);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n1046
                           , QN => n574);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => OUT2(16), QN
                           => n1869);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n1047
                           , QN => n571);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => OUT2(15), QN
                           => n1870);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n1048
                           , QN => n568);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => OUT2(14), QN
                           => n1871);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n1049
                           , QN => n565);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => OUT2(13), QN
                           => n1872);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n1050
                           , QN => n562);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => OUT2(12), QN
                           => n1873);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n1051
                           , QN => n559);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => OUT2(11), QN
                           => n1874);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n1052
                           , QN => n556);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => OUT2(10), QN
                           => n1875);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n1053,
                           QN => n553);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => OUT2(9), QN 
                           => n1876);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => n1054,
                           QN => n550);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => OUT2(8), QN 
                           => n1877);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => n1055,
                           QN => n547);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => OUT2(7), QN 
                           => n1878);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => n1056,
                           QN => n544);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => OUT2(6), QN 
                           => n1879);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => n1057,
                           QN => n541);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => OUT2(5), QN 
                           => n1880);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => n1058,
                           QN => n538);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => OUT2(4), QN 
                           => n1881);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => n1059,
                           QN => n535);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => OUT2(3), QN 
                           => n1882);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n1060,
                           QN => n532);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => OUT2(2), QN 
                           => n1883);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n1061,
                           QN => n529);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => OUT2(1), QN 
                           => n1884);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n1062,
                           QN => n522);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => OUT2(0), QN 
                           => n1885);
   OUT1_reg_63_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => OUT1(63), QN
                           => n1886);
   OUT1_reg_62_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => OUT1(62), QN
                           => n1887);
   OUT1_reg_61_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => OUT1(61), QN
                           => n1888);
   OUT1_reg_60_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => OUT1(60), QN
                           => n1889);
   OUT1_reg_59_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => OUT1(59), QN
                           => n1890);
   OUT1_reg_58_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => OUT1(58), QN
                           => n1891);
   OUT1_reg_57_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => OUT1(57), QN
                           => n1892);
   OUT1_reg_56_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => OUT1(56), QN
                           => n1893);
   OUT1_reg_55_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => OUT1(55), QN
                           => n1894);
   OUT1_reg_54_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => OUT1(54), QN
                           => n1895);
   OUT1_reg_53_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => OUT1(53), QN
                           => n1896);
   OUT1_reg_52_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => OUT1(52), QN
                           => n1897);
   OUT1_reg_51_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => OUT1(51), QN
                           => n1898);
   OUT1_reg_50_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => OUT1(50), QN
                           => n1899);
   OUT1_reg_49_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => OUT1(49), QN
                           => n1900);
   OUT1_reg_48_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => OUT1(48), QN
                           => n1901);
   OUT1_reg_47_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => OUT1(47), QN
                           => n1902);
   OUT1_reg_46_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => OUT1(46), QN
                           => n1903);
   OUT1_reg_45_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => OUT1(45), QN
                           => n1904);
   OUT1_reg_44_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => OUT1(44), QN
                           => n1905);
   OUT1_reg_43_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => OUT1(43), QN
                           => n1906);
   OUT1_reg_42_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => OUT1(42), QN
                           => n1907);
   OUT1_reg_41_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => OUT1(41), QN
                           => n1908);
   OUT1_reg_40_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => OUT1(40), QN
                           => n1909);
   OUT1_reg_39_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => OUT1(39), QN
                           => n1910);
   OUT1_reg_38_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => OUT1(38), QN
                           => n1911);
   OUT1_reg_37_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => OUT1(37), QN
                           => n1912);
   OUT1_reg_36_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => OUT1(36), QN
                           => n1913);
   OUT1_reg_35_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => OUT1(35), QN
                           => n1914);
   OUT1_reg_34_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => OUT1(34), QN
                           => n1915);
   OUT1_reg_33_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => OUT1(33), QN
                           => n1916);
   OUT1_reg_32_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => OUT1(32), QN
                           => n1917);
   OUT1_reg_31_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => OUT1(31), QN
                           => n1918);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => OUT1(30), QN
                           => n1919);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => OUT1(29), QN
                           => n1920);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => OUT1(28), QN
                           => n1921);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => OUT1(27), QN
                           => n1922);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => OUT1(26), QN
                           => n1923);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => OUT1(25), QN
                           => n1924);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => OUT1(24), QN
                           => n1925);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => OUT1(23), QN
                           => n1926);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => OUT1(22), QN
                           => n1927);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => OUT1(21), QN
                           => n1928);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => OUT1(20), QN
                           => n1929);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => OUT1(19), QN
                           => n1930);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => OUT1(18), QN
                           => n1931);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => OUT1(17), QN
                           => n1932);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => OUT1(16), QN
                           => n1933);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => OUT1(15), QN
                           => n1934);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => OUT1(14), QN
                           => n1935);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => OUT1(13), QN
                           => n1936);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => OUT1(12), QN
                           => n1937);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => OUT1(11), QN
                           => n1938);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => OUT1(10), QN
                           => n1939);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => OUT1(9), QN 
                           => n1940);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => OUT1(8), QN 
                           => n1941);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => OUT1(7), QN 
                           => n1942);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => OUT1(6), QN 
                           => n1943);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => OUT1(5), QN 
                           => n1944);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => OUT1(4), QN 
                           => n1945);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => OUT1(3), QN 
                           => n1946);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => OUT1(2), QN 
                           => n1947);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => OUT1(1), QN 
                           => n1948);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => OUT1(0), QN 
                           => n1949);
   U859 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n2050, A3 => ADD_RD1(1), 
                           ZN => n521);
   U860 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n2021, A3 => ADD_RD2(1), 
                           ZN => n735);
   U861 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n873, A3 => ADD_WR(1), ZN 
                           => n872);
   U862 : NAND3_X1 port map( A1 => n873, A2 => n2061, A3 => ADD_WR(1), ZN => 
                           n936);
   U863 : NAND3_X1 port map( A1 => n873, A2 => n2062, A3 => ADD_WR(0), ZN => 
                           n975);
   U864 : NAND3_X1 port map( A1 => n2061, A2 => n2062, A3 => n873, ZN => n998);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => n537, 
                           QN => n1818);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => n534, 
                           QN => n1819);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => n531, 
                           QN => n1820);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => n528, 
                           QN => n1821);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => n730,
                           QN => n415);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => n702,
                           QN => n1200);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => n698,
                           QN => n1202);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => n694,
                           QN => n1204);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => n622,
                           QN => n1793);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => n618,
                           QN => n1794);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => n614,
                           QN => n1795);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => n610,
                           QN => n1796);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => n606,
                           QN => n1797);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => n602,
                           QN => n1798);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => n598,
                           QN => n1799);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => n594,
                           QN => n1800);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => n590,
                           QN => n1801);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => n586,
                           QN => n1802);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => n582,
                           QN => n1803);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => n579,
                           QN => n1804);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => n576,
                           QN => n1805);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => n573,
                           QN => n1806);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => n570,
                           QN => n1807);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => n567,
                           QN => n1808);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => n564,
                           QN => n1809);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => n561,
                           QN => n1810);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => n558,
                           QN => n1811);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => n555, 
                           QN => n1812);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => n552, 
                           QN => n1813);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => n549, 
                           QN => n1814);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => n546, 
                           QN => n1815);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => n543, 
                           QN => n1816);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => n540, 
                           QN => n1817);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => n731,
                           QN => n1694);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => n727,
                           QN => n1695);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => n724,
                           QN => n1696);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => n721,
                           QN => n1697);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => n718,
                           QN => n1698);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => n715,
                           QN => n1699);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => n712,
                           QN => n1700);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => n709,
                           QN => n1701);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => n706,
                           QN => n1702);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => n703,
                           QN => n1703);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => n699,
                           QN => n1704);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => n695,
                           QN => n1705);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => n691,
                           QN => n1706);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => n688,
                           QN => n1707);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => n685,
                           QN => n1708);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => n682,
                           QN => n1709);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => n679,
                           QN => n1710);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => n676,
                           QN => n1711);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => n673,
                           QN => n1712);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => n670,
                           QN => n1713);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => n667,
                           QN => n1714);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => n664,
                           QN => n1715);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => n661,
                           QN => n1716);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => n658,
                           QN => n1717);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => n655,
                           QN => n1718);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => n652,
                           QN => n1719);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => n649,
                           QN => n1720);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => n646,
                           QN => n1721);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => n643,
                           QN => n1722);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => n640,
                           QN => n1723);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => n637,
                           QN => n1724);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => n634,
                           QN => n1725);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => n631,
                           QN => n1726);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => n628,
                           QN => n1727);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n625,
                           QN => n1728);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => n621,
                           QN => n1729);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => n617,
                           QN => n1730);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => n613,
                           QN => n1731);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => n609,
                           QN => n1732);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => n605,
                           QN => n1733);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => n601,
                           QN => n1734);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => n597,
                           QN => n1735);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => n593,
                           QN => n1736);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => n589,
                           QN => n1737);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => n585,
                           QN => n1738);
   U3 : BUF_X1 port map( A => n521, Z => n2053);
   U4 : BUF_X1 port map( A => n521, Z => n2052);
   U5 : BUF_X1 port map( A => n521, Z => n2051);
   U6 : BUF_X1 port map( A => n735, Z => n2025);
   U7 : BUF_X1 port map( A => n735, Z => n2024);
   U8 : BUF_X1 port map( A => n735, Z => n2023);
   U9 : BUF_X1 port map( A => n735, Z => n2022);
   U10 : BUF_X1 port map( A => n521, Z => n2055);
   U11 : BUF_X1 port map( A => n521, Z => n2054);
   U12 : BUF_X1 port map( A => n735, Z => n2026);
   U13 : BUF_X1 port map( A => n742, Z => n1990);
   U14 : BUF_X1 port map( A => n742, Z => n1989);
   U15 : BUF_X1 port map( A => n742, Z => n1988);
   U16 : BUF_X1 port map( A => n742, Z => n1987);
   U17 : BUF_X1 port map( A => n741, Z => n1992);
   U18 : BUF_X1 port map( A => n875, Z => n1980);
   U19 : BUF_X1 port map( A => n938, Z => n1968);
   U20 : BUF_X1 port map( A => n978, Z => n1956);
   U21 : BUF_X1 port map( A => n876, Z => n1978);
   U22 : BUF_X1 port map( A => n876, Z => n1977);
   U23 : BUF_X1 port map( A => n876, Z => n1976);
   U24 : BUF_X1 port map( A => n876, Z => n1975);
   U25 : BUF_X1 port map( A => n876, Z => n1974);
   U26 : BUF_X1 port map( A => n939, Z => n1966);
   U27 : BUF_X1 port map( A => n939, Z => n1965);
   U28 : BUF_X1 port map( A => n939, Z => n1964);
   U29 : BUF_X1 port map( A => n939, Z => n1963);
   U30 : BUF_X1 port map( A => n939, Z => n1962);
   U31 : BUF_X1 port map( A => n979, Z => n1954);
   U32 : BUF_X1 port map( A => n979, Z => n1953);
   U33 : BUF_X1 port map( A => n979, Z => n1952);
   U34 : BUF_X1 port map( A => n979, Z => n1951);
   U35 : BUF_X1 port map( A => n979, Z => n1950);
   U36 : BUF_X1 port map( A => n742, Z => n1986);
   U37 : BUF_X1 port map( A => n526, Z => n2037);
   U38 : BUF_X1 port map( A => n526, Z => n2038);
   U39 : BUF_X1 port map( A => n527, Z => n2030);
   U40 : BUF_X1 port map( A => n527, Z => n2032);
   U41 : BUF_X1 port map( A => n527, Z => n2031);
   U42 : BUF_X1 port map( A => n523, Z => n2045);
   U43 : BUF_X1 port map( A => n523, Z => n2046);
   U44 : BUF_X1 port map( A => n523, Z => n2047);
   U45 : BUF_X1 port map( A => n523, Z => n2048);
   U46 : BUF_X1 port map( A => n523, Z => n2049);
   U47 : BUF_X1 port map( A => n736, Z => n2016);
   U48 : BUF_X1 port map( A => n736, Z => n2017);
   U49 : BUF_X1 port map( A => n736, Z => n2018);
   U50 : BUF_X1 port map( A => n736, Z => n2019);
   U51 : BUF_X1 port map( A => n736, Z => n2020);
   U52 : BUF_X1 port map( A => n525, Z => n2040);
   U53 : BUF_X1 port map( A => n525, Z => n2041);
   U54 : BUF_X1 port map( A => n525, Z => n2042);
   U55 : BUF_X1 port map( A => n525, Z => n2043);
   U56 : BUF_X1 port map( A => n738, Z => n2014);
   U57 : BUF_X1 port map( A => n738, Z => n2013);
   U58 : BUF_X1 port map( A => n738, Z => n2012);
   U59 : BUF_X1 port map( A => n738, Z => n2011);
   U60 : BUF_X1 port map( A => n738, Z => n2010);
   U61 : BUF_X1 port map( A => n739, Z => n2008);
   U62 : BUF_X1 port map( A => n739, Z => n2007);
   U63 : BUF_X1 port map( A => n739, Z => n2006);
   U64 : BUF_X1 port map( A => n739, Z => n2005);
   U65 : BUF_X1 port map( A => n739, Z => n2004);
   U66 : BUF_X1 port map( A => n740, Z => n2002);
   U67 : BUF_X1 port map( A => n740, Z => n2001);
   U68 : BUF_X1 port map( A => n740, Z => n2000);
   U69 : BUF_X1 port map( A => n740, Z => n1999);
   U70 : BUF_X1 port map( A => n740, Z => n1998);
   U71 : BUF_X1 port map( A => n741, Z => n1996);
   U72 : BUF_X1 port map( A => n741, Z => n1995);
   U73 : BUF_X1 port map( A => n741, Z => n1994);
   U74 : BUF_X1 port map( A => n741, Z => n1993);
   U75 : BUF_X1 port map( A => n875, Z => n1984);
   U76 : BUF_X1 port map( A => n875, Z => n1983);
   U77 : BUF_X1 port map( A => n875, Z => n1982);
   U78 : BUF_X1 port map( A => n875, Z => n1981);
   U79 : BUF_X1 port map( A => n938, Z => n1972);
   U80 : BUF_X1 port map( A => n938, Z => n1971);
   U81 : BUF_X1 port map( A => n938, Z => n1970);
   U82 : BUF_X1 port map( A => n938, Z => n1969);
   U83 : BUF_X1 port map( A => n978, Z => n1960);
   U84 : BUF_X1 port map( A => n978, Z => n1959);
   U85 : BUF_X1 port map( A => n978, Z => n1958);
   U86 : BUF_X1 port map( A => n978, Z => n1957);
   U87 : BUF_X1 port map( A => n526, Z => n2034);
   U88 : BUF_X1 port map( A => n526, Z => n2036);
   U89 : BUF_X1 port map( A => n527, Z => n2029);
   U90 : BUF_X1 port map( A => n527, Z => n2028);
   U91 : BUF_X1 port map( A => n526, Z => n2035);
   U92 : BUF_X1 port map( A => n525, Z => n2039);
   U93 : NAND2_X1 port map( A1 => n734, A2 => n872, ZN => n741);
   U94 : NAND2_X1 port map( A1 => n734, A2 => n936, ZN => n875);
   U95 : NAND2_X1 port map( A1 => n734, A2 => n1980, ZN => n876);
   U96 : NAND2_X1 port map( A1 => n734, A2 => n975, ZN => n938);
   U97 : NAND2_X1 port map( A1 => n734, A2 => n1968, ZN => n939);
   U98 : NAND2_X1 port map( A1 => n734, A2 => n998, ZN => n978);
   U99 : NAND2_X1 port map( A1 => n734, A2 => n1956, ZN => n979);
   U100 : OAI22_X1 port map( A1 => n538, A2 => n1997, B1 => n1990, B2 => n751, 
                           ZN => n1620);
   U101 : OAI22_X1 port map( A1 => n541, A2 => n1996, B1 => n1990, B2 => n753, 
                           ZN => n1618);
   U102 : OAI22_X1 port map( A1 => n544, A2 => n1996, B1 => n1990, B2 => n755, 
                           ZN => n1616);
   U103 : OAI22_X1 port map( A1 => n547, A2 => n1996, B1 => n1990, B2 => n757, 
                           ZN => n1614);
   U104 : OAI22_X1 port map( A1 => n550, A2 => n1996, B1 => n1990, B2 => n759, 
                           ZN => n1612);
   U105 : OAI22_X1 port map( A1 => n553, A2 => n1996, B1 => n1990, B2 => n761, 
                           ZN => n1610);
   U106 : OAI22_X1 port map( A1 => n556, A2 => n1996, B1 => n1990, B2 => n763, 
                           ZN => n1608);
   U107 : OAI22_X1 port map( A1 => n559, A2 => n1996, B1 => n1990, B2 => n765, 
                           ZN => n1606);
   U108 : OAI22_X1 port map( A1 => n562, A2 => n1996, B1 => n1990, B2 => n767, 
                           ZN => n1604);
   U109 : OAI22_X1 port map( A1 => n565, A2 => n1996, B1 => n1990, B2 => n769, 
                           ZN => n1602);
   U110 : OAI22_X1 port map( A1 => n568, A2 => n1996, B1 => n1990, B2 => n771, 
                           ZN => n1600);
   U111 : OAI22_X1 port map( A1 => n571, A2 => n1996, B1 => n1990, B2 => n773, 
                           ZN => n1598);
   U112 : OAI22_X1 port map( A1 => n574, A2 => n1996, B1 => n1989, B2 => n775, 
                           ZN => n1596);
   U113 : OAI22_X1 port map( A1 => n577, A2 => n1995, B1 => n1989, B2 => n777, 
                           ZN => n1594);
   U114 : OAI22_X1 port map( A1 => n580, A2 => n1995, B1 => n1989, B2 => n779, 
                           ZN => n1592);
   U115 : OAI22_X1 port map( A1 => n583, A2 => n1995, B1 => n1989, B2 => n781, 
                           ZN => n1590);
   U116 : OAI22_X1 port map( A1 => n587, A2 => n1995, B1 => n1989, B2 => n783, 
                           ZN => n1588);
   U117 : OAI22_X1 port map( A1 => n591, A2 => n1995, B1 => n1989, B2 => n785, 
                           ZN => n1586);
   U118 : OAI22_X1 port map( A1 => n595, A2 => n1995, B1 => n1989, B2 => n787, 
                           ZN => n1584);
   U119 : OAI22_X1 port map( A1 => n599, A2 => n1995, B1 => n1989, B2 => n789, 
                           ZN => n1582);
   U120 : OAI22_X1 port map( A1 => n603, A2 => n1995, B1 => n1989, B2 => n791, 
                           ZN => n1580);
   U121 : OAI22_X1 port map( A1 => n607, A2 => n1995, B1 => n1989, B2 => n793, 
                           ZN => n1578);
   U122 : OAI22_X1 port map( A1 => n611, A2 => n1995, B1 => n1989, B2 => n795, 
                           ZN => n1576);
   U123 : OAI22_X1 port map( A1 => n615, A2 => n1995, B1 => n1989, B2 => n797, 
                           ZN => n1574);
   U124 : OAI22_X1 port map( A1 => n619, A2 => n1995, B1 => n1988, B2 => n799, 
                           ZN => n1572);
   U125 : OAI22_X1 port map( A1 => n623, A2 => n1994, B1 => n1988, B2 => n801, 
                           ZN => n1570);
   U126 : OAI22_X1 port map( A1 => n626, A2 => n1994, B1 => n1988, B2 => n803, 
                           ZN => n1568);
   U127 : OAI22_X1 port map( A1 => n629, A2 => n1994, B1 => n1988, B2 => n805, 
                           ZN => n1566);
   U128 : OAI22_X1 port map( A1 => n632, A2 => n1994, B1 => n1988, B2 => n807, 
                           ZN => n1564);
   U129 : OAI22_X1 port map( A1 => n635, A2 => n1994, B1 => n1988, B2 => n809, 
                           ZN => n1562);
   U130 : OAI22_X1 port map( A1 => n638, A2 => n1994, B1 => n1988, B2 => n811, 
                           ZN => n1560);
   U131 : OAI22_X1 port map( A1 => n641, A2 => n1994, B1 => n1988, B2 => n813, 
                           ZN => n1558);
   U132 : OAI22_X1 port map( A1 => n644, A2 => n1994, B1 => n1988, B2 => n815, 
                           ZN => n1556);
   U133 : OAI22_X1 port map( A1 => n647, A2 => n1994, B1 => n1988, B2 => n817, 
                           ZN => n1554);
   U134 : OAI22_X1 port map( A1 => n650, A2 => n1994, B1 => n1988, B2 => n819, 
                           ZN => n1552);
   U135 : OAI22_X1 port map( A1 => n653, A2 => n1994, B1 => n1988, B2 => n821, 
                           ZN => n1550);
   U136 : OAI22_X1 port map( A1 => n656, A2 => n1994, B1 => n1987, B2 => n823, 
                           ZN => n1548);
   U137 : OAI22_X1 port map( A1 => n659, A2 => n1993, B1 => n1987, B2 => n825, 
                           ZN => n1546);
   U138 : OAI22_X1 port map( A1 => n662, A2 => n1993, B1 => n1987, B2 => n827, 
                           ZN => n1544);
   U139 : OAI22_X1 port map( A1 => n665, A2 => n1993, B1 => n1987, B2 => n829, 
                           ZN => n1542);
   U140 : OAI22_X1 port map( A1 => n668, A2 => n1993, B1 => n1987, B2 => n831, 
                           ZN => n1540);
   U141 : OAI22_X1 port map( A1 => n671, A2 => n1993, B1 => n1987, B2 => n833, 
                           ZN => n1538);
   U142 : OAI22_X1 port map( A1 => n674, A2 => n1993, B1 => n1987, B2 => n835, 
                           ZN => n1536);
   U143 : OAI22_X1 port map( A1 => n677, A2 => n1993, B1 => n1987, B2 => n837, 
                           ZN => n1534);
   U144 : OAI22_X1 port map( A1 => n680, A2 => n1993, B1 => n1987, B2 => n839, 
                           ZN => n1532);
   U145 : OAI22_X1 port map( A1 => n683, A2 => n1993, B1 => n1987, B2 => n841, 
                           ZN => n1530);
   U146 : OAI22_X1 port map( A1 => n686, A2 => n1993, B1 => n1987, B2 => n843, 
                           ZN => n1528);
   U147 : OAI22_X1 port map( A1 => n689, A2 => n1993, B1 => n1987, B2 => n845, 
                           ZN => n1526);
   U148 : OAI22_X1 port map( A1 => n522, A2 => n1997, B1 => n1991, B2 => n743, 
                           ZN => n1628);
   U149 : OAI22_X1 port map( A1 => n529, A2 => n1997, B1 => n1991, B2 => n745, 
                           ZN => n1626);
   U150 : OAI22_X1 port map( A1 => n532, A2 => n1997, B1 => n1991, B2 => n747, 
                           ZN => n1624);
   U151 : OAI22_X1 port map( A1 => n535, A2 => n1997, B1 => n1991, B2 => n749, 
                           ZN => n1622);
   U152 : OAI22_X1 port map( A1 => n692, A2 => n1993, B1 => n1986, B2 => n847, 
                           ZN => n1524);
   U153 : OAI22_X1 port map( A1 => n696, A2 => n1992, B1 => n1986, B2 => n849, 
                           ZN => n1522);
   U154 : OAI22_X1 port map( A1 => n700, A2 => n1992, B1 => n1986, B2 => n851, 
                           ZN => n1520);
   U155 : OAI22_X1 port map( A1 => n704, A2 => n1992, B1 => n1986, B2 => n853, 
                           ZN => n1518);
   U156 : OAI22_X1 port map( A1 => n707, A2 => n1992, B1 => n1986, B2 => n855, 
                           ZN => n1516);
   U157 : OAI22_X1 port map( A1 => n710, A2 => n1992, B1 => n1986, B2 => n857, 
                           ZN => n1514);
   U158 : OAI22_X1 port map( A1 => n713, A2 => n1992, B1 => n1986, B2 => n859, 
                           ZN => n1512);
   U159 : OAI22_X1 port map( A1 => n716, A2 => n1992, B1 => n1986, B2 => n861, 
                           ZN => n1510);
   U160 : OAI22_X1 port map( A1 => n719, A2 => n1992, B1 => n1986, B2 => n863, 
                           ZN => n1508);
   U161 : OAI22_X1 port map( A1 => n722, A2 => n1992, B1 => n1986, B2 => n865, 
                           ZN => n1506);
   U162 : OAI22_X1 port map( A1 => n725, A2 => n1992, B1 => n1986, B2 => n867, 
                           ZN => n1504);
   U163 : OAI22_X1 port map( A1 => n728, A2 => n1992, B1 => n1986, B2 => n871, 
                           ZN => n1502);
   U164 : NAND2_X1 port map( A1 => n734, A2 => n1992, ZN => n742);
   U165 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n873);
   U166 : AND3_X1 port map( A1 => n2059, A2 => n2060, A3 => n2050, ZN => n526);
   U167 : AND3_X1 port map( A1 => n2050, A2 => n2060, A3 => ADD_RD1(0), ZN => 
                           n527);
   U168 : AND3_X1 port map( A1 => n2050, A2 => n2059, A3 => ADD_RD1(1), ZN => 
                           n525);
   U169 : AND3_X1 port map( A1 => n2021, A2 => n2058, A3 => ADD_RD2(0), ZN => 
                           n740);
   U170 : AND3_X1 port map( A1 => n2021, A2 => n2057, A3 => ADD_RD2(1), ZN => 
                           n738);
   U171 : AND3_X1 port map( A1 => n2057, A2 => n2058, A3 => n2021, ZN => n739);
   U172 : AND2_X1 port map( A1 => RD2, A2 => n734, ZN => n736);
   U173 : AND2_X1 port map( A1 => RD1, A2 => n734, ZN => n523);
   U174 : OAI22_X1 port map( A1 => n874, A2 => n1985, B1 => n743, B2 => n1979, 
                           ZN => n1501);
   U175 : OAI22_X1 port map( A1 => n877, A2 => n1985, B1 => n745, B2 => n1979, 
                           ZN => n1500);
   U176 : OAI22_X1 port map( A1 => n878, A2 => n1985, B1 => n747, B2 => n1979, 
                           ZN => n1499);
   U177 : OAI22_X1 port map( A1 => n879, A2 => n1985, B1 => n749, B2 => n1979, 
                           ZN => n1498);
   U178 : OAI22_X1 port map( A1 => n1821, A2 => n1973, B1 => n743, B2 => n1967,
                           ZN => n1437);
   U179 : OAI22_X1 port map( A1 => n1820, A2 => n1973, B1 => n745, B2 => n1967,
                           ZN => n1436);
   U180 : OAI22_X1 port map( A1 => n1819, A2 => n1973, B1 => n747, B2 => n1967,
                           ZN => n1435);
   U181 : OAI22_X1 port map( A1 => n1818, A2 => n1973, B1 => n749, B2 => n1967,
                           ZN => n1434);
   U182 : OAI22_X1 port map( A1 => n977, A2 => n1961, B1 => n743, B2 => n1955, 
                           ZN => n1373);
   U183 : OAI22_X1 port map( A1 => n980, A2 => n1961, B1 => n745, B2 => n1955, 
                           ZN => n1372);
   U184 : OAI22_X1 port map( A1 => n981, A2 => n1961, B1 => n747, B2 => n1955, 
                           ZN => n1371);
   U185 : OAI22_X1 port map( A1 => n982, A2 => n1961, B1 => n749, B2 => n1955, 
                           ZN => n1370);
   U186 : OAI22_X1 port map( A1 => n880, A2 => n1985, B1 => n751, B2 => n1978, 
                           ZN => n1497);
   U187 : OAI22_X1 port map( A1 => n881, A2 => n1984, B1 => n753, B2 => n1978, 
                           ZN => n1496);
   U188 : OAI22_X1 port map( A1 => n882, A2 => n1984, B1 => n755, B2 => n1978, 
                           ZN => n1495);
   U189 : OAI22_X1 port map( A1 => n883, A2 => n1984, B1 => n757, B2 => n1978, 
                           ZN => n1494);
   U190 : OAI22_X1 port map( A1 => n884, A2 => n1984, B1 => n759, B2 => n1978, 
                           ZN => n1493);
   U191 : OAI22_X1 port map( A1 => n885, A2 => n1984, B1 => n761, B2 => n1978, 
                           ZN => n1492);
   U192 : OAI22_X1 port map( A1 => n886, A2 => n1984, B1 => n763, B2 => n1978, 
                           ZN => n1491);
   U193 : OAI22_X1 port map( A1 => n887, A2 => n1984, B1 => n765, B2 => n1978, 
                           ZN => n1490);
   U194 : OAI22_X1 port map( A1 => n888, A2 => n1984, B1 => n767, B2 => n1978, 
                           ZN => n1489);
   U195 : OAI22_X1 port map( A1 => n889, A2 => n1984, B1 => n769, B2 => n1978, 
                           ZN => n1488);
   U196 : OAI22_X1 port map( A1 => n890, A2 => n1984, B1 => n771, B2 => n1978, 
                           ZN => n1487);
   U197 : OAI22_X1 port map( A1 => n891, A2 => n1984, B1 => n773, B2 => n1978, 
                           ZN => n1486);
   U198 : OAI22_X1 port map( A1 => n892, A2 => n1984, B1 => n775, B2 => n1977, 
                           ZN => n1485);
   U199 : OAI22_X1 port map( A1 => n893, A2 => n1983, B1 => n777, B2 => n1977, 
                           ZN => n1484);
   U200 : OAI22_X1 port map( A1 => n894, A2 => n1983, B1 => n779, B2 => n1977, 
                           ZN => n1483);
   U201 : OAI22_X1 port map( A1 => n895, A2 => n1983, B1 => n781, B2 => n1977, 
                           ZN => n1482);
   U202 : OAI22_X1 port map( A1 => n896, A2 => n1983, B1 => n783, B2 => n1977, 
                           ZN => n1481);
   U203 : OAI22_X1 port map( A1 => n897, A2 => n1983, B1 => n785, B2 => n1977, 
                           ZN => n1480);
   U204 : OAI22_X1 port map( A1 => n898, A2 => n1983, B1 => n787, B2 => n1977, 
                           ZN => n1479);
   U205 : OAI22_X1 port map( A1 => n899, A2 => n1983, B1 => n789, B2 => n1977, 
                           ZN => n1478);
   U206 : OAI22_X1 port map( A1 => n900, A2 => n1983, B1 => n791, B2 => n1977, 
                           ZN => n1477);
   U207 : OAI22_X1 port map( A1 => n901, A2 => n1983, B1 => n793, B2 => n1977, 
                           ZN => n1476);
   U208 : OAI22_X1 port map( A1 => n902, A2 => n1983, B1 => n795, B2 => n1977, 
                           ZN => n1475);
   U209 : OAI22_X1 port map( A1 => n903, A2 => n1983, B1 => n797, B2 => n1977, 
                           ZN => n1474);
   U210 : OAI22_X1 port map( A1 => n904, A2 => n1983, B1 => n799, B2 => n1976, 
                           ZN => n1473);
   U211 : OAI22_X1 port map( A1 => n905, A2 => n1982, B1 => n801, B2 => n1976, 
                           ZN => n1472);
   U212 : OAI22_X1 port map( A1 => n906, A2 => n1982, B1 => n803, B2 => n1976, 
                           ZN => n1471);
   U213 : OAI22_X1 port map( A1 => n907, A2 => n1982, B1 => n805, B2 => n1976, 
                           ZN => n1470);
   U214 : OAI22_X1 port map( A1 => n908, A2 => n1982, B1 => n807, B2 => n1976, 
                           ZN => n1469);
   U215 : OAI22_X1 port map( A1 => n909, A2 => n1982, B1 => n809, B2 => n1976, 
                           ZN => n1468);
   U216 : OAI22_X1 port map( A1 => n910, A2 => n1982, B1 => n811, B2 => n1976, 
                           ZN => n1467);
   U217 : OAI22_X1 port map( A1 => n911, A2 => n1982, B1 => n813, B2 => n1976, 
                           ZN => n1466);
   U218 : OAI22_X1 port map( A1 => n912, A2 => n1982, B1 => n815, B2 => n1976, 
                           ZN => n1465);
   U219 : OAI22_X1 port map( A1 => n913, A2 => n1982, B1 => n817, B2 => n1976, 
                           ZN => n1464);
   U220 : OAI22_X1 port map( A1 => n914, A2 => n1982, B1 => n819, B2 => n1976, 
                           ZN => n1463);
   U221 : OAI22_X1 port map( A1 => n915, A2 => n1982, B1 => n821, B2 => n1976, 
                           ZN => n1462);
   U222 : OAI22_X1 port map( A1 => n916, A2 => n1982, B1 => n823, B2 => n1975, 
                           ZN => n1461);
   U223 : OAI22_X1 port map( A1 => n917, A2 => n1981, B1 => n825, B2 => n1975, 
                           ZN => n1460);
   U224 : OAI22_X1 port map( A1 => n918, A2 => n1981, B1 => n827, B2 => n1975, 
                           ZN => n1459);
   U225 : OAI22_X1 port map( A1 => n919, A2 => n1981, B1 => n829, B2 => n1975, 
                           ZN => n1458);
   U226 : OAI22_X1 port map( A1 => n920, A2 => n1981, B1 => n831, B2 => n1975, 
                           ZN => n1457);
   U227 : OAI22_X1 port map( A1 => n921, A2 => n1981, B1 => n833, B2 => n1975, 
                           ZN => n1456);
   U228 : OAI22_X1 port map( A1 => n922, A2 => n1981, B1 => n835, B2 => n1975, 
                           ZN => n1455);
   U229 : OAI22_X1 port map( A1 => n923, A2 => n1981, B1 => n837, B2 => n1975, 
                           ZN => n1454);
   U230 : OAI22_X1 port map( A1 => n924, A2 => n1981, B1 => n839, B2 => n1975, 
                           ZN => n1453);
   U231 : OAI22_X1 port map( A1 => n925, A2 => n1981, B1 => n841, B2 => n1975, 
                           ZN => n1452);
   U232 : OAI22_X1 port map( A1 => n926, A2 => n1981, B1 => n843, B2 => n1975, 
                           ZN => n1451);
   U233 : OAI22_X1 port map( A1 => n927, A2 => n1981, B1 => n845, B2 => n1975, 
                           ZN => n1450);
   U234 : OAI22_X1 port map( A1 => n1204, A2 => n1981, B1 => n847, B2 => n1974,
                           ZN => n1449);
   U235 : OAI22_X1 port map( A1 => n1202, A2 => n1980, B1 => n849, B2 => n1974,
                           ZN => n1448);
   U236 : OAI22_X1 port map( A1 => n1200, A2 => n1980, B1 => n851, B2 => n1974,
                           ZN => n1447);
   U237 : OAI22_X1 port map( A1 => n928, A2 => n1980, B1 => n853, B2 => n1974, 
                           ZN => n1446);
   U238 : OAI22_X1 port map( A1 => n929, A2 => n1980, B1 => n855, B2 => n1974, 
                           ZN => n1445);
   U239 : OAI22_X1 port map( A1 => n930, A2 => n1980, B1 => n857, B2 => n1974, 
                           ZN => n1444);
   U240 : OAI22_X1 port map( A1 => n931, A2 => n1980, B1 => n859, B2 => n1974, 
                           ZN => n1443);
   U241 : OAI22_X1 port map( A1 => n932, A2 => n1980, B1 => n861, B2 => n1974, 
                           ZN => n1442);
   U242 : OAI22_X1 port map( A1 => n933, A2 => n1980, B1 => n863, B2 => n1974, 
                           ZN => n1441);
   U243 : OAI22_X1 port map( A1 => n934, A2 => n1980, B1 => n865, B2 => n1974, 
                           ZN => n1440);
   U244 : OAI22_X1 port map( A1 => n935, A2 => n1980, B1 => n867, B2 => n1974, 
                           ZN => n1439);
   U245 : OAI22_X1 port map( A1 => n415, A2 => n1980, B1 => n871, B2 => n1974, 
                           ZN => n1438);
   U246 : OAI22_X1 port map( A1 => n1817, A2 => n1973, B1 => n751, B2 => n1966,
                           ZN => n1433);
   U247 : OAI22_X1 port map( A1 => n1816, A2 => n1972, B1 => n753, B2 => n1966,
                           ZN => n1432);
   U248 : OAI22_X1 port map( A1 => n1815, A2 => n1972, B1 => n755, B2 => n1966,
                           ZN => n1431);
   U249 : OAI22_X1 port map( A1 => n1814, A2 => n1972, B1 => n757, B2 => n1966,
                           ZN => n1430);
   U250 : OAI22_X1 port map( A1 => n1813, A2 => n1972, B1 => n759, B2 => n1966,
                           ZN => n1429);
   U251 : OAI22_X1 port map( A1 => n1812, A2 => n1972, B1 => n761, B2 => n1966,
                           ZN => n1428);
   U252 : OAI22_X1 port map( A1 => n1811, A2 => n1972, B1 => n763, B2 => n1966,
                           ZN => n1427);
   U253 : OAI22_X1 port map( A1 => n1810, A2 => n1972, B1 => n765, B2 => n1966,
                           ZN => n1426);
   U254 : OAI22_X1 port map( A1 => n1809, A2 => n1972, B1 => n767, B2 => n1966,
                           ZN => n1425);
   U255 : OAI22_X1 port map( A1 => n1808, A2 => n1972, B1 => n769, B2 => n1966,
                           ZN => n1424);
   U256 : OAI22_X1 port map( A1 => n1807, A2 => n1972, B1 => n771, B2 => n1966,
                           ZN => n1423);
   U257 : OAI22_X1 port map( A1 => n1806, A2 => n1972, B1 => n773, B2 => n1966,
                           ZN => n1422);
   U258 : OAI22_X1 port map( A1 => n1805, A2 => n1972, B1 => n775, B2 => n1965,
                           ZN => n1421);
   U259 : OAI22_X1 port map( A1 => n1804, A2 => n1971, B1 => n777, B2 => n1965,
                           ZN => n1420);
   U260 : OAI22_X1 port map( A1 => n1803, A2 => n1971, B1 => n779, B2 => n1965,
                           ZN => n1419);
   U261 : OAI22_X1 port map( A1 => n1802, A2 => n1971, B1 => n781, B2 => n1965,
                           ZN => n1418);
   U262 : OAI22_X1 port map( A1 => n1801, A2 => n1971, B1 => n783, B2 => n1965,
                           ZN => n1417);
   U263 : OAI22_X1 port map( A1 => n1800, A2 => n1971, B1 => n785, B2 => n1965,
                           ZN => n1416);
   U264 : OAI22_X1 port map( A1 => n1799, A2 => n1971, B1 => n787, B2 => n1965,
                           ZN => n1415);
   U265 : OAI22_X1 port map( A1 => n1798, A2 => n1971, B1 => n789, B2 => n1965,
                           ZN => n1414);
   U266 : OAI22_X1 port map( A1 => n1797, A2 => n1971, B1 => n791, B2 => n1965,
                           ZN => n1413);
   U267 : OAI22_X1 port map( A1 => n1796, A2 => n1971, B1 => n793, B2 => n1965,
                           ZN => n1412);
   U268 : OAI22_X1 port map( A1 => n1795, A2 => n1971, B1 => n795, B2 => n1965,
                           ZN => n1411);
   U269 : OAI22_X1 port map( A1 => n1794, A2 => n1971, B1 => n797, B2 => n1965,
                           ZN => n1410);
   U270 : OAI22_X1 port map( A1 => n1793, A2 => n1971, B1 => n799, B2 => n1964,
                           ZN => n1409);
   U271 : OAI22_X1 port map( A1 => n940, A2 => n1970, B1 => n801, B2 => n1964, 
                           ZN => n1408);
   U272 : OAI22_X1 port map( A1 => n941, A2 => n1970, B1 => n803, B2 => n1964, 
                           ZN => n1407);
   U273 : OAI22_X1 port map( A1 => n942, A2 => n1970, B1 => n805, B2 => n1964, 
                           ZN => n1406);
   U274 : OAI22_X1 port map( A1 => n943, A2 => n1970, B1 => n807, B2 => n1964, 
                           ZN => n1405);
   U275 : OAI22_X1 port map( A1 => n944, A2 => n1970, B1 => n809, B2 => n1964, 
                           ZN => n1404);
   U276 : OAI22_X1 port map( A1 => n945, A2 => n1970, B1 => n811, B2 => n1964, 
                           ZN => n1403);
   U277 : OAI22_X1 port map( A1 => n946, A2 => n1970, B1 => n813, B2 => n1964, 
                           ZN => n1402);
   U278 : OAI22_X1 port map( A1 => n947, A2 => n1970, B1 => n815, B2 => n1964, 
                           ZN => n1401);
   U279 : OAI22_X1 port map( A1 => n948, A2 => n1970, B1 => n817, B2 => n1964, 
                           ZN => n1400);
   U280 : OAI22_X1 port map( A1 => n949, A2 => n1970, B1 => n819, B2 => n1964, 
                           ZN => n1399);
   U281 : OAI22_X1 port map( A1 => n950, A2 => n1970, B1 => n821, B2 => n1964, 
                           ZN => n1398);
   U282 : OAI22_X1 port map( A1 => n951, A2 => n1970, B1 => n823, B2 => n1963, 
                           ZN => n1397);
   U283 : OAI22_X1 port map( A1 => n952, A2 => n1969, B1 => n825, B2 => n1963, 
                           ZN => n1396);
   U284 : OAI22_X1 port map( A1 => n953, A2 => n1969, B1 => n827, B2 => n1963, 
                           ZN => n1395);
   U285 : OAI22_X1 port map( A1 => n954, A2 => n1969, B1 => n829, B2 => n1963, 
                           ZN => n1394);
   U286 : OAI22_X1 port map( A1 => n955, A2 => n1969, B1 => n831, B2 => n1963, 
                           ZN => n1393);
   U287 : OAI22_X1 port map( A1 => n956, A2 => n1969, B1 => n833, B2 => n1963, 
                           ZN => n1392);
   U288 : OAI22_X1 port map( A1 => n957, A2 => n1969, B1 => n835, B2 => n1963, 
                           ZN => n1391);
   U289 : OAI22_X1 port map( A1 => n958, A2 => n1969, B1 => n837, B2 => n1963, 
                           ZN => n1390);
   U290 : OAI22_X1 port map( A1 => n959, A2 => n1969, B1 => n839, B2 => n1963, 
                           ZN => n1389);
   U291 : OAI22_X1 port map( A1 => n960, A2 => n1969, B1 => n841, B2 => n1963, 
                           ZN => n1388);
   U292 : OAI22_X1 port map( A1 => n961, A2 => n1969, B1 => n843, B2 => n1963, 
                           ZN => n1387);
   U293 : OAI22_X1 port map( A1 => n962, A2 => n1969, B1 => n845, B2 => n1963, 
                           ZN => n1386);
   U294 : OAI22_X1 port map( A1 => n963, A2 => n1969, B1 => n847, B2 => n1962, 
                           ZN => n1385);
   U295 : OAI22_X1 port map( A1 => n964, A2 => n1968, B1 => n849, B2 => n1962, 
                           ZN => n1384);
   U296 : OAI22_X1 port map( A1 => n965, A2 => n1968, B1 => n851, B2 => n1962, 
                           ZN => n1383);
   U297 : OAI22_X1 port map( A1 => n966, A2 => n1968, B1 => n853, B2 => n1962, 
                           ZN => n1382);
   U298 : OAI22_X1 port map( A1 => n967, A2 => n1968, B1 => n855, B2 => n1962, 
                           ZN => n1381);
   U299 : OAI22_X1 port map( A1 => n968, A2 => n1968, B1 => n857, B2 => n1962, 
                           ZN => n1380);
   U300 : OAI22_X1 port map( A1 => n969, A2 => n1968, B1 => n859, B2 => n1962, 
                           ZN => n1379);
   U301 : OAI22_X1 port map( A1 => n970, A2 => n1968, B1 => n861, B2 => n1962, 
                           ZN => n1378);
   U302 : OAI22_X1 port map( A1 => n971, A2 => n1968, B1 => n863, B2 => n1962, 
                           ZN => n1377);
   U303 : OAI22_X1 port map( A1 => n972, A2 => n1968, B1 => n865, B2 => n1962, 
                           ZN => n1376);
   U304 : OAI22_X1 port map( A1 => n973, A2 => n1968, B1 => n867, B2 => n1962, 
                           ZN => n1375);
   U305 : OAI22_X1 port map( A1 => n974, A2 => n1968, B1 => n871, B2 => n1962, 
                           ZN => n1374);
   U306 : OAI22_X1 port map( A1 => n983, A2 => n1961, B1 => n751, B2 => n1954, 
                           ZN => n1369);
   U307 : OAI22_X1 port map( A1 => n984, A2 => n1960, B1 => n753, B2 => n1954, 
                           ZN => n1368);
   U308 : OAI22_X1 port map( A1 => n985, A2 => n1960, B1 => n755, B2 => n1954, 
                           ZN => n1367);
   U309 : OAI22_X1 port map( A1 => n986, A2 => n1960, B1 => n757, B2 => n1954, 
                           ZN => n1366);
   U310 : OAI22_X1 port map( A1 => n987, A2 => n1960, B1 => n759, B2 => n1954, 
                           ZN => n1365);
   U311 : OAI22_X1 port map( A1 => n988, A2 => n1960, B1 => n761, B2 => n1954, 
                           ZN => n1364);
   U312 : OAI22_X1 port map( A1 => n989, A2 => n1960, B1 => n763, B2 => n1954, 
                           ZN => n1363);
   U313 : OAI22_X1 port map( A1 => n990, A2 => n1960, B1 => n765, B2 => n1954, 
                           ZN => n1362);
   U314 : OAI22_X1 port map( A1 => n991, A2 => n1960, B1 => n767, B2 => n1954, 
                           ZN => n1361);
   U315 : OAI22_X1 port map( A1 => n992, A2 => n1960, B1 => n769, B2 => n1954, 
                           ZN => n1360);
   U316 : OAI22_X1 port map( A1 => n993, A2 => n1960, B1 => n771, B2 => n1954, 
                           ZN => n1359);
   U317 : OAI22_X1 port map( A1 => n994, A2 => n1960, B1 => n773, B2 => n1954, 
                           ZN => n1358);
   U318 : OAI22_X1 port map( A1 => n995, A2 => n1960, B1 => n775, B2 => n1953, 
                           ZN => n1357);
   U319 : OAI22_X1 port map( A1 => n996, A2 => n1959, B1 => n777, B2 => n1953, 
                           ZN => n1356);
   U320 : OAI22_X1 port map( A1 => n997, A2 => n1959, B1 => n779, B2 => n1953, 
                           ZN => n1355);
   U321 : OAI22_X1 port map( A1 => n1738, A2 => n1959, B1 => n781, B2 => n1953,
                           ZN => n1354);
   U322 : OAI22_X1 port map( A1 => n1737, A2 => n1959, B1 => n783, B2 => n1953,
                           ZN => n1353);
   U323 : OAI22_X1 port map( A1 => n1736, A2 => n1959, B1 => n785, B2 => n1953,
                           ZN => n1352);
   U324 : OAI22_X1 port map( A1 => n1735, A2 => n1959, B1 => n787, B2 => n1953,
                           ZN => n1351);
   U325 : OAI22_X1 port map( A1 => n1734, A2 => n1959, B1 => n789, B2 => n1953,
                           ZN => n1350);
   U326 : OAI22_X1 port map( A1 => n1733, A2 => n1959, B1 => n791, B2 => n1953,
                           ZN => n1349);
   U327 : OAI22_X1 port map( A1 => n1732, A2 => n1959, B1 => n793, B2 => n1953,
                           ZN => n1348);
   U328 : OAI22_X1 port map( A1 => n1731, A2 => n1959, B1 => n795, B2 => n1953,
                           ZN => n1347);
   U329 : OAI22_X1 port map( A1 => n1730, A2 => n1959, B1 => n797, B2 => n1953,
                           ZN => n1346);
   U330 : OAI22_X1 port map( A1 => n1729, A2 => n1959, B1 => n799, B2 => n1952,
                           ZN => n1345);
   U331 : OAI22_X1 port map( A1 => n1728, A2 => n1958, B1 => n801, B2 => n1952,
                           ZN => n1344);
   U332 : OAI22_X1 port map( A1 => n1727, A2 => n1958, B1 => n803, B2 => n1952,
                           ZN => n1343);
   U333 : OAI22_X1 port map( A1 => n1726, A2 => n1958, B1 => n805, B2 => n1952,
                           ZN => n1342);
   U334 : OAI22_X1 port map( A1 => n1725, A2 => n1958, B1 => n807, B2 => n1952,
                           ZN => n1341);
   U335 : OAI22_X1 port map( A1 => n1724, A2 => n1958, B1 => n809, B2 => n1952,
                           ZN => n1340);
   U336 : OAI22_X1 port map( A1 => n1723, A2 => n1958, B1 => n811, B2 => n1952,
                           ZN => n1339);
   U337 : OAI22_X1 port map( A1 => n1722, A2 => n1958, B1 => n813, B2 => n1952,
                           ZN => n1338);
   U338 : OAI22_X1 port map( A1 => n1721, A2 => n1958, B1 => n815, B2 => n1952,
                           ZN => n1337);
   U339 : OAI22_X1 port map( A1 => n1720, A2 => n1958, B1 => n817, B2 => n1952,
                           ZN => n1336);
   U340 : OAI22_X1 port map( A1 => n1719, A2 => n1958, B1 => n819, B2 => n1952,
                           ZN => n1335);
   U341 : OAI22_X1 port map( A1 => n1718, A2 => n1958, B1 => n821, B2 => n1952,
                           ZN => n1334);
   U342 : OAI22_X1 port map( A1 => n1717, A2 => n1958, B1 => n823, B2 => n1951,
                           ZN => n1333);
   U343 : OAI22_X1 port map( A1 => n1716, A2 => n1957, B1 => n825, B2 => n1951,
                           ZN => n1332);
   U344 : OAI22_X1 port map( A1 => n1715, A2 => n1957, B1 => n827, B2 => n1951,
                           ZN => n1331);
   U345 : OAI22_X1 port map( A1 => n1714, A2 => n1957, B1 => n829, B2 => n1951,
                           ZN => n1330);
   U346 : OAI22_X1 port map( A1 => n1713, A2 => n1957, B1 => n831, B2 => n1951,
                           ZN => n1329);
   U347 : OAI22_X1 port map( A1 => n1712, A2 => n1957, B1 => n833, B2 => n1951,
                           ZN => n1328);
   U348 : OAI22_X1 port map( A1 => n1711, A2 => n1957, B1 => n835, B2 => n1951,
                           ZN => n1327);
   U349 : OAI22_X1 port map( A1 => n1710, A2 => n1957, B1 => n837, B2 => n1951,
                           ZN => n1326);
   U350 : OAI22_X1 port map( A1 => n1709, A2 => n1957, B1 => n839, B2 => n1951,
                           ZN => n1325);
   U351 : OAI22_X1 port map( A1 => n1708, A2 => n1957, B1 => n841, B2 => n1951,
                           ZN => n1324);
   U352 : OAI22_X1 port map( A1 => n1707, A2 => n1957, B1 => n843, B2 => n1951,
                           ZN => n1323);
   U353 : OAI22_X1 port map( A1 => n1706, A2 => n1957, B1 => n845, B2 => n1951,
                           ZN => n1322);
   U354 : OAI22_X1 port map( A1 => n1705, A2 => n1957, B1 => n847, B2 => n1950,
                           ZN => n1321);
   U355 : OAI22_X1 port map( A1 => n1704, A2 => n1956, B1 => n849, B2 => n1950,
                           ZN => n1320);
   U356 : OAI22_X1 port map( A1 => n1703, A2 => n1956, B1 => n851, B2 => n1950,
                           ZN => n1319);
   U357 : OAI22_X1 port map( A1 => n1702, A2 => n1956, B1 => n853, B2 => n1950,
                           ZN => n1318);
   U358 : OAI22_X1 port map( A1 => n1701, A2 => n1956, B1 => n855, B2 => n1950,
                           ZN => n1317);
   U359 : OAI22_X1 port map( A1 => n1700, A2 => n1956, B1 => n857, B2 => n1950,
                           ZN => n1316);
   U360 : OAI22_X1 port map( A1 => n1699, A2 => n1956, B1 => n859, B2 => n1950,
                           ZN => n1315);
   U361 : OAI22_X1 port map( A1 => n1698, A2 => n1956, B1 => n861, B2 => n1950,
                           ZN => n1314);
   U362 : OAI22_X1 port map( A1 => n1697, A2 => n1956, B1 => n863, B2 => n1950,
                           ZN => n1313);
   U363 : OAI22_X1 port map( A1 => n1696, A2 => n1956, B1 => n865, B2 => n1950,
                           ZN => n1312);
   U364 : OAI22_X1 port map( A1 => n1695, A2 => n1956, B1 => n867, B2 => n1950,
                           ZN => n1311);
   U365 : OAI22_X1 port map( A1 => n1694, A2 => n1956, B1 => n871, B2 => n1950,
                           ZN => n1310);
   U366 : OAI221_X1 port map( B1 => n2055, B2 => n562, C1 => n1937, C2 => n2046
                           , A => n563, ZN => n1681);
   U367 : AOI222_X1 port map( A1 => n52, A2 => n2039, B1 => n180, B2 => n2035, 
                           C1 => n2032, C2 => n564, ZN => n563);
   U368 : OAI221_X1 port map( B1 => n2055, B2 => n565, C1 => n1936, C2 => n2046
                           , A => n566, ZN => n1680);
   U369 : AOI222_X1 port map( A1 => n51, A2 => n2040, B1 => n179, B2 => n2035, 
                           C1 => n2032, C2 => n567, ZN => n566);
   U370 : OAI221_X1 port map( B1 => n2055, B2 => n568, C1 => n1935, C2 => n2046
                           , A => n569, ZN => n1679);
   U371 : AOI222_X1 port map( A1 => n50, A2 => n2040, B1 => n178, B2 => n2035, 
                           C1 => n2032, C2 => n570, ZN => n569);
   U372 : OAI221_X1 port map( B1 => n2055, B2 => n571, C1 => n1934, C2 => n2047
                           , A => n572, ZN => n1678);
   U373 : AOI222_X1 port map( A1 => n49, A2 => n2040, B1 => n177, B2 => n2035, 
                           C1 => n2031, C2 => n573, ZN => n572);
   U374 : OAI221_X1 port map( B1 => n2054, B2 => n574, C1 => n1933, C2 => n2046
                           , A => n575, ZN => n1677);
   U375 : AOI222_X1 port map( A1 => n48, A2 => n2040, B1 => n176, B2 => n2035, 
                           C1 => n2031, C2 => n576, ZN => n575);
   U376 : OAI221_X1 port map( B1 => n2054, B2 => n577, C1 => n1932, C2 => n2046
                           , A => n578, ZN => n1676);
   U377 : AOI222_X1 port map( A1 => n47, A2 => n2040, B1 => n175, B2 => n2035, 
                           C1 => n2031, C2 => n579, ZN => n578);
   U378 : OAI221_X1 port map( B1 => n2054, B2 => n580, C1 => n1931, C2 => n2046
                           , A => n581, ZN => n1675);
   U379 : AOI222_X1 port map( A1 => n46, A2 => n2040, B1 => n174, B2 => n2035, 
                           C1 => n2031, C2 => n582, ZN => n581);
   U380 : OAI221_X1 port map( B1 => n538, B2 => n2026, C1 => n1881, C2 => n2016
                           , A => n750, ZN => n1621);
   U381 : AOI222_X1 port map( A1 => n2014, A2 => n60, B1 => n2008, B2 => n188, 
                           C1 => n2002, C2 => n540, ZN => n750);
   U382 : OAI221_X1 port map( B1 => n541, B2 => n2026, C1 => n1880, C2 => n2016
                           , A => n752, ZN => n1619);
   U383 : AOI222_X1 port map( A1 => n2014, A2 => n59, B1 => n2008, B2 => n187, 
                           C1 => n2002, C2 => n543, ZN => n752);
   U384 : OAI221_X1 port map( B1 => n544, B2 => n2026, C1 => n1879, C2 => n2016
                           , A => n754, ZN => n1617);
   U385 : AOI222_X1 port map( A1 => n2014, A2 => n58, B1 => n2008, B2 => n186, 
                           C1 => n2002, C2 => n546, ZN => n754);
   U386 : OAI221_X1 port map( B1 => n547, B2 => n2026, C1 => n1878, C2 => n2016
                           , A => n756, ZN => n1615);
   U387 : AOI222_X1 port map( A1 => n2014, A2 => n57, B1 => n2008, B2 => n185, 
                           C1 => n2002, C2 => n549, ZN => n756);
   U388 : OAI221_X1 port map( B1 => n550, B2 => n2026, C1 => n1877, C2 => n2016
                           , A => n758, ZN => n1613);
   U389 : AOI222_X1 port map( A1 => n2014, A2 => n56, B1 => n2008, B2 => n184, 
                           C1 => n2002, C2 => n552, ZN => n758);
   U390 : OAI221_X1 port map( B1 => n553, B2 => n2026, C1 => n1876, C2 => n2016
                           , A => n760, ZN => n1611);
   U391 : AOI222_X1 port map( A1 => n2014, A2 => n55, B1 => n2008, B2 => n183, 
                           C1 => n2002, C2 => n555, ZN => n760);
   U392 : OAI221_X1 port map( B1 => n556, B2 => n2026, C1 => n1875, C2 => n2016
                           , A => n762, ZN => n1609);
   U393 : AOI222_X1 port map( A1 => n2014, A2 => n54, B1 => n2008, B2 => n182, 
                           C1 => n2002, C2 => n558, ZN => n762);
   U394 : OAI221_X1 port map( B1 => n559, B2 => n2026, C1 => n1874, C2 => n2016
                           , A => n764, ZN => n1607);
   U395 : AOI222_X1 port map( A1 => n2014, A2 => n53, B1 => n2008, B2 => n181, 
                           C1 => n2002, C2 => n561, ZN => n764);
   U396 : OAI221_X1 port map( B1 => n562, B2 => n2026, C1 => n1873, C2 => n2017
                           , A => n766, ZN => n1605);
   U397 : AOI222_X1 port map( A1 => n2014, A2 => n52, B1 => n2008, B2 => n180, 
                           C1 => n2002, C2 => n564, ZN => n766);
   U398 : OAI221_X1 port map( B1 => n565, B2 => n2026, C1 => n1872, C2 => n2017
                           , A => n768, ZN => n1603);
   U399 : AOI222_X1 port map( A1 => n2014, A2 => n51, B1 => n2008, B2 => n179, 
                           C1 => n2002, C2 => n567, ZN => n768);
   U400 : OAI221_X1 port map( B1 => n568, B2 => n2026, C1 => n1871, C2 => n2017
                           , A => n770, ZN => n1601);
   U401 : AOI222_X1 port map( A1 => n2014, A2 => n50, B1 => n2008, B2 => n178, 
                           C1 => n2002, C2 => n570, ZN => n770);
   U402 : OAI221_X1 port map( B1 => n571, B2 => n2026, C1 => n1870, C2 => n2018
                           , A => n772, ZN => n1599);
   U403 : AOI222_X1 port map( A1 => n2014, A2 => n49, B1 => n2008, B2 => n177, 
                           C1 => n2002, C2 => n573, ZN => n772);
   U404 : OAI221_X1 port map( B1 => n574, B2 => n2025, C1 => n1869, C2 => n2017
                           , A => n774, ZN => n1597);
   U405 : AOI222_X1 port map( A1 => n2013, A2 => n48, B1 => n2007, B2 => n176, 
                           C1 => n2001, C2 => n576, ZN => n774);
   U406 : OAI221_X1 port map( B1 => n577, B2 => n2025, C1 => n1868, C2 => n2017
                           , A => n776, ZN => n1595);
   U407 : AOI222_X1 port map( A1 => n2013, A2 => n47, B1 => n2007, B2 => n175, 
                           C1 => n2001, C2 => n579, ZN => n776);
   U408 : OAI221_X1 port map( B1 => n580, B2 => n2025, C1 => n1867, C2 => n2017
                           , A => n778, ZN => n1593);
   U409 : AOI222_X1 port map( A1 => n2013, A2 => n46, B1 => n2007, B2 => n174, 
                           C1 => n2001, C2 => n582, ZN => n778);
   U410 : OAI221_X1 port map( B1 => n2051, B2 => n716, C1 => n1890, C2 => n2050
                           , A => n717, ZN => n1634);
   U411 : AOI222_X1 port map( A1 => n5, A2 => n2043, B1 => n2038, B2 => n718, 
                           C1 => n69, C2 => n2028, ZN => n717);
   U412 : OAI221_X1 port map( B1 => n2051, B2 => n722, C1 => n1888, C2 => n2050
                           , A => n723, ZN => n1632);
   U413 : AOI222_X1 port map( A1 => n3, A2 => n2043, B1 => n2038, B2 => n724, 
                           C1 => n67, C2 => n2028, ZN => n723);
   U414 : OAI221_X1 port map( B1 => n2051, B2 => n725, C1 => n1887, C2 => n2050
                           , A => n726, ZN => n1631);
   U415 : AOI222_X1 port map( A1 => n2, A2 => n2043, B1 => n2038, B2 => n727, 
                           C1 => n66, C2 => n2028, ZN => n726);
   U416 : OAI221_X1 port map( B1 => n2051, B2 => n728, C1 => n1886, C2 => n2050
                           , A => n729, ZN => n1630);
   U417 : AOI222_X1 port map( A1 => n2044, A2 => n730, B1 => n2036, B2 => n731,
                           C1 => n65, C2 => n2028, ZN => n729);
   U418 : OAI221_X1 port map( B1 => n623, B2 => n2024, C1 => n1856, C2 => n2018
                           , A => n800, ZN => n1571);
   U419 : AOI222_X1 port map( A1 => n2012, A2 => n35, B1 => n2006, B2 => n625, 
                           C1 => n2000, C2 => n99, ZN => n800);
   U420 : OAI221_X1 port map( B1 => n626, B2 => n2024, C1 => n1855, C2 => n2018
                           , A => n802, ZN => n1569);
   U421 : AOI222_X1 port map( A1 => n2012, A2 => n34, B1 => n2006, B2 => n628, 
                           C1 => n2000, C2 => n98, ZN => n802);
   U422 : OAI221_X1 port map( B1 => n629, B2 => n2024, C1 => n1854, C2 => n2018
                           , A => n804, ZN => n1567);
   U423 : AOI222_X1 port map( A1 => n2012, A2 => n33, B1 => n2006, B2 => n631, 
                           C1 => n2000, C2 => n97, ZN => n804);
   U424 : OAI221_X1 port map( B1 => n632, B2 => n2024, C1 => n1853, C2 => n2018
                           , A => n806, ZN => n1565);
   U425 : AOI222_X1 port map( A1 => n2012, A2 => n32, B1 => n2006, B2 => n634, 
                           C1 => n2000, C2 => n96, ZN => n806);
   U426 : OAI221_X1 port map( B1 => n635, B2 => n2024, C1 => n1852, C2 => n2018
                           , A => n808, ZN => n1563);
   U427 : AOI222_X1 port map( A1 => n2012, A2 => n31, B1 => n2006, B2 => n637, 
                           C1 => n2000, C2 => n95, ZN => n808);
   U428 : OAI221_X1 port map( B1 => n638, B2 => n2024, C1 => n1851, C2 => n2018
                           , A => n810, ZN => n1561);
   U429 : AOI222_X1 port map( A1 => n2012, A2 => n30, B1 => n2006, B2 => n640, 
                           C1 => n2000, C2 => n94, ZN => n810);
   U430 : OAI221_X1 port map( B1 => n641, B2 => n2024, C1 => n1850, C2 => n2018
                           , A => n812, ZN => n1559);
   U431 : AOI222_X1 port map( A1 => n2012, A2 => n29, B1 => n2006, B2 => n643, 
                           C1 => n2000, C2 => n93, ZN => n812);
   U432 : OAI221_X1 port map( B1 => n644, B2 => n2024, C1 => n1849, C2 => n2019
                           , A => n814, ZN => n1557);
   U433 : AOI222_X1 port map( A1 => n2012, A2 => n28, B1 => n2006, B2 => n646, 
                           C1 => n2000, C2 => n92, ZN => n814);
   U434 : OAI221_X1 port map( B1 => n647, B2 => n2024, C1 => n1848, C2 => n2019
                           , A => n816, ZN => n1555);
   U435 : AOI222_X1 port map( A1 => n2012, A2 => n27, B1 => n2006, B2 => n649, 
                           C1 => n2000, C2 => n91, ZN => n816);
   U436 : OAI221_X1 port map( B1 => n650, B2 => n2024, C1 => n1847, C2 => n2019
                           , A => n818, ZN => n1553);
   U437 : AOI222_X1 port map( A1 => n2012, A2 => n26, B1 => n2006, B2 => n652, 
                           C1 => n2000, C2 => n90, ZN => n818);
   U438 : OAI221_X1 port map( B1 => n653, B2 => n2024, C1 => n1846, C2 => n2019
                           , A => n820, ZN => n1551);
   U439 : AOI222_X1 port map( A1 => n2012, A2 => n25, B1 => n2006, B2 => n655, 
                           C1 => n2000, C2 => n89, ZN => n820);
   U440 : OAI221_X1 port map( B1 => n656, B2 => n2023, C1 => n1845, C2 => n2019
                           , A => n822, ZN => n1549);
   U441 : AOI222_X1 port map( A1 => n2011, A2 => n24, B1 => n2005, B2 => n658, 
                           C1 => n1999, C2 => n88, ZN => n822);
   U442 : OAI221_X1 port map( B1 => n659, B2 => n2023, C1 => n1844, C2 => n2019
                           , A => n824, ZN => n1547);
   U443 : AOI222_X1 port map( A1 => n2011, A2 => n23, B1 => n2005, B2 => n661, 
                           C1 => n1999, C2 => n87, ZN => n824);
   U444 : OAI221_X1 port map( B1 => n662, B2 => n2023, C1 => n1843, C2 => n2019
                           , A => n826, ZN => n1545);
   U445 : AOI222_X1 port map( A1 => n2011, A2 => n22, B1 => n2005, B2 => n664, 
                           C1 => n1999, C2 => n86, ZN => n826);
   U446 : OAI221_X1 port map( B1 => n665, B2 => n2023, C1 => n1842, C2 => n2019
                           , A => n828, ZN => n1543);
   U447 : AOI222_X1 port map( A1 => n2011, A2 => n21, B1 => n2005, B2 => n667, 
                           C1 => n1999, C2 => n85, ZN => n828);
   U448 : OAI221_X1 port map( B1 => n668, B2 => n2023, C1 => n1841, C2 => n2019
                           , A => n830, ZN => n1541);
   U449 : AOI222_X1 port map( A1 => n2011, A2 => n20, B1 => n2005, B2 => n670, 
                           C1 => n1999, C2 => n84, ZN => n830);
   U450 : OAI221_X1 port map( B1 => n671, B2 => n2023, C1 => n1840, C2 => n2019
                           , A => n832, ZN => n1539);
   U451 : AOI222_X1 port map( A1 => n2011, A2 => n19, B1 => n2005, B2 => n673, 
                           C1 => n1999, C2 => n83, ZN => n832);
   U452 : OAI221_X1 port map( B1 => n674, B2 => n2023, C1 => n1839, C2 => n2019
                           , A => n834, ZN => n1537);
   U453 : AOI222_X1 port map( A1 => n2011, A2 => n18, B1 => n2005, B2 => n676, 
                           C1 => n1999, C2 => n82, ZN => n834);
   U454 : OAI221_X1 port map( B1 => n677, B2 => n2023, C1 => n1838, C2 => n2019
                           , A => n836, ZN => n1535);
   U455 : AOI222_X1 port map( A1 => n2011, A2 => n17, B1 => n2005, B2 => n679, 
                           C1 => n1999, C2 => n81, ZN => n836);
   U456 : OAI221_X1 port map( B1 => n680, B2 => n2023, C1 => n1837, C2 => n2020
                           , A => n838, ZN => n1533);
   U457 : AOI222_X1 port map( A1 => n2011, A2 => n16, B1 => n2005, B2 => n682, 
                           C1 => n1999, C2 => n80, ZN => n838);
   U458 : OAI221_X1 port map( B1 => n683, B2 => n2023, C1 => n1836, C2 => n2020
                           , A => n840, ZN => n1531);
   U459 : AOI222_X1 port map( A1 => n2011, A2 => n15, B1 => n2005, B2 => n685, 
                           C1 => n1999, C2 => n79, ZN => n840);
   U460 : OAI221_X1 port map( B1 => n686, B2 => n2023, C1 => n1835, C2 => n2020
                           , A => n842, ZN => n1529);
   U461 : AOI222_X1 port map( A1 => n2011, A2 => n14, B1 => n2005, B2 => n688, 
                           C1 => n1999, C2 => n78, ZN => n842);
   U462 : OAI221_X1 port map( B1 => n689, B2 => n2023, C1 => n1834, C2 => n2020
                           , A => n844, ZN => n1527);
   U463 : AOI222_X1 port map( A1 => n2011, A2 => n13, B1 => n2005, B2 => n691, 
                           C1 => n1999, C2 => n77, ZN => n844);
   U464 : OAI221_X1 port map( B1 => n692, B2 => n2022, C1 => n1833, C2 => n2020
                           , A => n846, ZN => n1525);
   U465 : AOI222_X1 port map( A1 => n2010, A2 => n694, B1 => n2004, B2 => n695,
                           C1 => n1998, C2 => n76, ZN => n846);
   U466 : OAI221_X1 port map( B1 => n696, B2 => n2022, C1 => n1832, C2 => n2020
                           , A => n848, ZN => n1523);
   U467 : AOI222_X1 port map( A1 => n2010, A2 => n698, B1 => n2004, B2 => n699,
                           C1 => n1998, C2 => n75, ZN => n848);
   U468 : OAI221_X1 port map( B1 => n700, B2 => n2022, C1 => n1831, C2 => n2020
                           , A => n850, ZN => n1521);
   U469 : AOI222_X1 port map( A1 => n2010, A2 => n702, B1 => n2004, B2 => n703,
                           C1 => n1998, C2 => n74, ZN => n850);
   U470 : OAI221_X1 port map( B1 => n704, B2 => n2022, C1 => n1830, C2 => n2020
                           , A => n852, ZN => n1519);
   U471 : AOI222_X1 port map( A1 => n2010, A2 => n9, B1 => n2004, B2 => n706, 
                           C1 => n1998, C2 => n73, ZN => n852);
   U472 : OAI221_X1 port map( B1 => n707, B2 => n2022, C1 => n1829, C2 => n2020
                           , A => n854, ZN => n1517);
   U473 : AOI222_X1 port map( A1 => n2010, A2 => n8, B1 => n2004, B2 => n709, 
                           C1 => n1998, C2 => n72, ZN => n854);
   U474 : OAI221_X1 port map( B1 => n710, B2 => n2022, C1 => n1828, C2 => n2020
                           , A => n856, ZN => n1515);
   U475 : AOI222_X1 port map( A1 => n2010, A2 => n7, B1 => n2004, B2 => n712, 
                           C1 => n1998, C2 => n71, ZN => n856);
   U476 : OAI221_X1 port map( B1 => n713, B2 => n2022, C1 => n1827, C2 => n2020
                           , A => n858, ZN => n1513);
   U477 : AOI222_X1 port map( A1 => n2010, A2 => n6, B1 => n2004, B2 => n715, 
                           C1 => n1998, C2 => n70, ZN => n858);
   U478 : OAI221_X1 port map( B1 => n716, B2 => n2022, C1 => n1826, C2 => n2021
                           , A => n860, ZN => n1511);
   U479 : AOI222_X1 port map( A1 => n2010, A2 => n5, B1 => n2004, B2 => n718, 
                           C1 => n1998, C2 => n69, ZN => n860);
   U480 : OAI221_X1 port map( B1 => n719, B2 => n2022, C1 => n1825, C2 => n2020
                           , A => n862, ZN => n1509);
   U481 : AOI222_X1 port map( A1 => n2010, A2 => n4, B1 => n2004, B2 => n721, 
                           C1 => n1998, C2 => n68, ZN => n862);
   U482 : OAI221_X1 port map( B1 => n722, B2 => n2022, C1 => n1824, C2 => n2021
                           , A => n864, ZN => n1507);
   U483 : AOI222_X1 port map( A1 => n2010, A2 => n3, B1 => n2004, B2 => n724, 
                           C1 => n1998, C2 => n67, ZN => n864);
   U484 : OAI221_X1 port map( B1 => n725, B2 => n2022, C1 => n1823, C2 => n2021
                           , A => n866, ZN => n1505);
   U485 : AOI222_X1 port map( A1 => n2010, A2 => n2, B1 => n2004, B2 => n727, 
                           C1 => n1998, C2 => n66, ZN => n866);
   U486 : OAI221_X1 port map( B1 => n728, B2 => n2022, C1 => n1822, C2 => n2021
                           , A => n868, ZN => n1503);
   U487 : AOI222_X1 port map( A1 => n2010, A2 => n730, B1 => n2004, B2 => n731,
                           C1 => n1998, C2 => n65, ZN => n868);
   U488 : INV_X1 port map( A => RESET, ZN => n734);
   U489 : OAI221_X1 port map( B1 => n2056, B2 => n522, C1 => n1949, C2 => n2045
                           , A => n524, ZN => n1693);
   U490 : AOI222_X1 port map( A1 => n64, A2 => n2041, B1 => n192, B2 => n2034, 
                           C1 => n2033, C2 => n528, ZN => n524);
   U491 : OAI221_X1 port map( B1 => n2056, B2 => n529, C1 => n1948, C2 => n2045
                           , A => n530, ZN => n1692);
   U492 : AOI222_X1 port map( A1 => n63, A2 => n2039, B1 => n191, B2 => n2034, 
                           C1 => n2033, C2 => n531, ZN => n530);
   U493 : OAI221_X1 port map( B1 => n2056, B2 => n532, C1 => n1947, C2 => n2045
                           , A => n533, ZN => n1691);
   U494 : AOI222_X1 port map( A1 => n62, A2 => n2039, B1 => n190, B2 => n2034, 
                           C1 => n2032, C2 => n534, ZN => n533);
   U495 : OAI221_X1 port map( B1 => n2056, B2 => n535, C1 => n1946, C2 => n2045
                           , A => n536, ZN => n1690);
   U496 : AOI222_X1 port map( A1 => n61, A2 => n2039, B1 => n189, B2 => n2034, 
                           C1 => n2032, C2 => n537, ZN => n536);
   U497 : OAI221_X1 port map( B1 => n2053, B2 => n619, C1 => n1921, C2 => n2047
                           , A => n620, ZN => n1665);
   U498 : AOI222_X1 port map( A1 => n36, A2 => n2041, B1 => n2036, B2 => n621, 
                           C1 => n2030, C2 => n622, ZN => n620);
   U499 : OAI221_X1 port map( B1 => n2053, B2 => n623, C1 => n1920, C2 => n2047
                           , A => n624, ZN => n1664);
   U500 : AOI222_X1 port map( A1 => n35, A2 => n2041, B1 => n2036, B2 => n625, 
                           C1 => n99, C2 => n2030, ZN => n624);
   U501 : OAI221_X1 port map( B1 => n2053, B2 => n626, C1 => n1919, C2 => n2047
                           , A => n627, ZN => n1663);
   U502 : AOI222_X1 port map( A1 => n34, A2 => n2041, B1 => n2036, B2 => n628, 
                           C1 => n98, C2 => n2030, ZN => n627);
   U503 : OAI221_X1 port map( B1 => n2053, B2 => n629, C1 => n1918, C2 => n2047
                           , A => n630, ZN => n1662);
   U504 : AOI222_X1 port map( A1 => n33, A2 => n2041, B1 => n2036, B2 => n631, 
                           C1 => n97, C2 => n2030, ZN => n630);
   U505 : OAI221_X1 port map( B1 => n2053, B2 => n632, C1 => n1917, C2 => n2047
                           , A => n633, ZN => n1661);
   U506 : AOI222_X1 port map( A1 => n32, A2 => n2041, B1 => n2036, B2 => n634, 
                           C1 => n96, C2 => n2030, ZN => n633);
   U507 : OAI221_X1 port map( B1 => n2053, B2 => n635, C1 => n1916, C2 => n2047
                           , A => n636, ZN => n1660);
   U508 : AOI222_X1 port map( A1 => n31, A2 => n2041, B1 => n2036, B2 => n637, 
                           C1 => n95, C2 => n2030, ZN => n636);
   U509 : OAI221_X1 port map( B1 => n2053, B2 => n638, C1 => n1915, C2 => n2047
                           , A => n639, ZN => n1659);
   U510 : AOI222_X1 port map( A1 => n30, A2 => n2041, B1 => n2036, B2 => n640, 
                           C1 => n94, C2 => n2030, ZN => n639);
   U511 : OAI221_X1 port map( B1 => n2053, B2 => n641, C1 => n1914, C2 => n2047
                           , A => n642, ZN => n1658);
   U512 : AOI222_X1 port map( A1 => n29, A2 => n2041, B1 => n2036, B2 => n643, 
                           C1 => n93, C2 => n2030, ZN => n642);
   U513 : OAI221_X1 port map( B1 => n2053, B2 => n644, C1 => n1913, C2 => n2048
                           , A => n645, ZN => n1657);
   U514 : AOI222_X1 port map( A1 => n28, A2 => n2042, B1 => n2036, B2 => n646, 
                           C1 => n92, C2 => n2030, ZN => n645);
   U515 : OAI221_X1 port map( B1 => n2053, B2 => n647, C1 => n1912, C2 => n2048
                           , A => n648, ZN => n1656);
   U516 : AOI222_X1 port map( A1 => n27, A2 => n2042, B1 => n2037, B2 => n649, 
                           C1 => n91, C2 => n2030, ZN => n648);
   U517 : OAI221_X1 port map( B1 => n2053, B2 => n650, C1 => n1911, C2 => n2048
                           , A => n651, ZN => n1655);
   U518 : AOI222_X1 port map( A1 => n26, A2 => n2042, B1 => n2037, B2 => n652, 
                           C1 => n90, C2 => n2030, ZN => n651);
   U519 : OAI221_X1 port map( B1 => n2053, B2 => n653, C1 => n1910, C2 => n2048
                           , A => n654, ZN => n1654);
   U520 : AOI222_X1 port map( A1 => n25, A2 => n2042, B1 => n2037, B2 => n655, 
                           C1 => n89, C2 => n2030, ZN => n654);
   U521 : OAI221_X1 port map( B1 => n2052, B2 => n656, C1 => n1909, C2 => n2048
                           , A => n657, ZN => n1653);
   U522 : AOI222_X1 port map( A1 => n24, A2 => n2042, B1 => n2037, B2 => n658, 
                           C1 => n88, C2 => n2029, ZN => n657);
   U523 : OAI221_X1 port map( B1 => n2052, B2 => n659, C1 => n1908, C2 => n2048
                           , A => n660, ZN => n1652);
   U524 : AOI222_X1 port map( A1 => n23, A2 => n2042, B1 => n2037, B2 => n661, 
                           C1 => n87, C2 => n2029, ZN => n660);
   U525 : OAI221_X1 port map( B1 => n2052, B2 => n662, C1 => n1907, C2 => n2048
                           , A => n663, ZN => n1651);
   U526 : AOI222_X1 port map( A1 => n22, A2 => n2042, B1 => n2037, B2 => n664, 
                           C1 => n86, C2 => n2029, ZN => n663);
   U527 : OAI221_X1 port map( B1 => n2052, B2 => n665, C1 => n1906, C2 => n2048
                           , A => n666, ZN => n1650);
   U528 : AOI222_X1 port map( A1 => n21, A2 => n2042, B1 => n2037, B2 => n667, 
                           C1 => n85, C2 => n2029, ZN => n666);
   U529 : OAI221_X1 port map( B1 => n2052, B2 => n668, C1 => n1905, C2 => n2048
                           , A => n669, ZN => n1649);
   U530 : AOI222_X1 port map( A1 => n20, A2 => n2042, B1 => n2037, B2 => n670, 
                           C1 => n84, C2 => n2029, ZN => n669);
   U531 : OAI221_X1 port map( B1 => n2052, B2 => n671, C1 => n1904, C2 => n2048
                           , A => n672, ZN => n1648);
   U532 : AOI222_X1 port map( A1 => n19, A2 => n2042, B1 => n2037, B2 => n673, 
                           C1 => n83, C2 => n2029, ZN => n672);
   U533 : OAI221_X1 port map( B1 => n2052, B2 => n674, C1 => n1903, C2 => n2048
                           , A => n675, ZN => n1647);
   U534 : AOI222_X1 port map( A1 => n18, A2 => n2042, B1 => n2037, B2 => n676, 
                           C1 => n82, C2 => n2029, ZN => n675);
   U535 : OAI221_X1 port map( B1 => n2052, B2 => n677, C1 => n1902, C2 => n2048
                           , A => n678, ZN => n1646);
   U536 : AOI222_X1 port map( A1 => n17, A2 => n2042, B1 => n2037, B2 => n679, 
                           C1 => n81, C2 => n2029, ZN => n678);
   U537 : OAI221_X1 port map( B1 => n2052, B2 => n680, C1 => n1901, C2 => n2049
                           , A => n681, ZN => n1645);
   U538 : AOI222_X1 port map( A1 => n16, A2 => n2043, B1 => n2037, B2 => n682, 
                           C1 => n80, C2 => n2029, ZN => n681);
   U539 : OAI221_X1 port map( B1 => n2052, B2 => n683, C1 => n1900, C2 => n2049
                           , A => n684, ZN => n1644);
   U540 : AOI222_X1 port map( A1 => n15, A2 => n2043, B1 => n2037, B2 => n685, 
                           C1 => n79, C2 => n2029, ZN => n684);
   U541 : OAI221_X1 port map( B1 => n2052, B2 => n686, C1 => n1899, C2 => n2049
                           , A => n687, ZN => n1643);
   U542 : AOI222_X1 port map( A1 => n14, A2 => n2043, B1 => n2038, B2 => n688, 
                           C1 => n78, C2 => n2029, ZN => n687);
   U543 : OAI221_X1 port map( B1 => n2052, B2 => n689, C1 => n1898, C2 => n2049
                           , A => n690, ZN => n1642);
   U544 : AOI222_X1 port map( A1 => n13, A2 => n2043, B1 => n2038, B2 => n691, 
                           C1 => n77, C2 => n2029, ZN => n690);
   U545 : OAI221_X1 port map( B1 => n2051, B2 => n692, C1 => n1897, C2 => n2049
                           , A => n693, ZN => n1641);
   U546 : AOI222_X1 port map( A1 => n2044, A2 => n694, B1 => n2038, B2 => n695,
                           C1 => n76, C2 => n2028, ZN => n693);
   U547 : OAI221_X1 port map( B1 => n2051, B2 => n696, C1 => n1896, C2 => n2049
                           , A => n697, ZN => n1640);
   U548 : AOI222_X1 port map( A1 => n2044, A2 => n698, B1 => n2038, B2 => n699,
                           C1 => n75, C2 => n2028, ZN => n697);
   U549 : OAI221_X1 port map( B1 => n2051, B2 => n700, C1 => n1895, C2 => n2049
                           , A => n701, ZN => n1639);
   U550 : AOI222_X1 port map( A1 => n2044, A2 => n702, B1 => n2038, B2 => n703,
                           C1 => n74, C2 => n2028, ZN => n701);
   U551 : OAI221_X1 port map( B1 => n2051, B2 => n704, C1 => n1894, C2 => n2049
                           , A => n705, ZN => n1638);
   U552 : AOI222_X1 port map( A1 => n9, A2 => n2043, B1 => n2038, B2 => n706, 
                           C1 => n73, C2 => n2028, ZN => n705);
   U553 : OAI221_X1 port map( B1 => n2051, B2 => n707, C1 => n1893, C2 => n2049
                           , A => n708, ZN => n1637);
   U554 : AOI222_X1 port map( A1 => n8, A2 => n2043, B1 => n2038, B2 => n709, 
                           C1 => n72, C2 => n2028, ZN => n708);
   U555 : OAI221_X1 port map( B1 => n2051, B2 => n710, C1 => n1892, C2 => n2049
                           , A => n711, ZN => n1636);
   U556 : AOI222_X1 port map( A1 => n7, A2 => n2043, B1 => n2038, B2 => n712, 
                           C1 => n71, C2 => n2028, ZN => n711);
   U557 : OAI221_X1 port map( B1 => n2051, B2 => n713, C1 => n1891, C2 => n2049
                           , A => n714, ZN => n1635);
   U558 : AOI222_X1 port map( A1 => n6, A2 => n2043, B1 => n2038, B2 => n715, 
                           C1 => n70, C2 => n2028, ZN => n714);
   U559 : OAI221_X1 port map( B1 => n2051, B2 => n719, C1 => n1889, C2 => n2049
                           , A => n720, ZN => n1633);
   U560 : AOI222_X1 port map( A1 => n4, A2 => n2043, B1 => n2038, B2 => n721, 
                           C1 => n68, C2 => n2028, ZN => n720);
   U561 : OAI221_X1 port map( B1 => n522, B2 => n2027, C1 => n1885, C2 => n2016
                           , A => n737, ZN => n1629);
   U562 : AOI222_X1 port map( A1 => n2015, A2 => n64, B1 => n2009, B2 => n192, 
                           C1 => n2003, C2 => n528, ZN => n737);
   U563 : OAI221_X1 port map( B1 => n529, B2 => n2027, C1 => n1884, C2 => n2016
                           , A => n744, ZN => n1627);
   U564 : AOI222_X1 port map( A1 => n2015, A2 => n63, B1 => n2009, B2 => n191, 
                           C1 => n2003, C2 => n531, ZN => n744);
   U565 : OAI221_X1 port map( B1 => n532, B2 => n2027, C1 => n1883, C2 => n2016
                           , A => n746, ZN => n1625);
   U566 : AOI222_X1 port map( A1 => n2015, A2 => n62, B1 => n2009, B2 => n190, 
                           C1 => n2003, C2 => n534, ZN => n746);
   U567 : OAI221_X1 port map( B1 => n535, B2 => n2027, C1 => n1882, C2 => n2016
                           , A => n748, ZN => n1623);
   U568 : AOI222_X1 port map( A1 => n2015, A2 => n61, B1 => n2009, B2 => n189, 
                           C1 => n2003, C2 => n537, ZN => n748);
   U569 : OAI221_X1 port map( B1 => n583, B2 => n2025, C1 => n1866, C2 => n2017
                           , A => n780, ZN => n1591);
   U570 : AOI222_X1 port map( A1 => n2013, A2 => n45, B1 => n2007, B2 => n585, 
                           C1 => n2001, C2 => n586, ZN => n780);
   U571 : OAI221_X1 port map( B1 => n587, B2 => n2025, C1 => n1865, C2 => n2017
                           , A => n782, ZN => n1589);
   U572 : AOI222_X1 port map( A1 => n2013, A2 => n44, B1 => n2007, B2 => n589, 
                           C1 => n2001, C2 => n590, ZN => n782);
   U573 : OAI221_X1 port map( B1 => n591, B2 => n2025, C1 => n1864, C2 => n2017
                           , A => n784, ZN => n1587);
   U574 : AOI222_X1 port map( A1 => n2013, A2 => n43, B1 => n2007, B2 => n593, 
                           C1 => n2001, C2 => n594, ZN => n784);
   U575 : OAI221_X1 port map( B1 => n595, B2 => n2025, C1 => n1863, C2 => n2017
                           , A => n786, ZN => n1585);
   U576 : AOI222_X1 port map( A1 => n2013, A2 => n42, B1 => n2007, B2 => n597, 
                           C1 => n2001, C2 => n598, ZN => n786);
   U577 : OAI221_X1 port map( B1 => n599, B2 => n2025, C1 => n1862, C2 => n2017
                           , A => n788, ZN => n1583);
   U578 : AOI222_X1 port map( A1 => n2013, A2 => n41, B1 => n2007, B2 => n601, 
                           C1 => n2001, C2 => n602, ZN => n788);
   U579 : OAI221_X1 port map( B1 => n603, B2 => n2025, C1 => n1861, C2 => n2017
                           , A => n790, ZN => n1581);
   U580 : AOI222_X1 port map( A1 => n2013, A2 => n40, B1 => n2007, B2 => n605, 
                           C1 => n2001, C2 => n606, ZN => n790);
   U581 : OAI221_X1 port map( B1 => n607, B2 => n2025, C1 => n1860, C2 => n2018
                           , A => n792, ZN => n1579);
   U582 : AOI222_X1 port map( A1 => n2013, A2 => n39, B1 => n2007, B2 => n609, 
                           C1 => n2001, C2 => n610, ZN => n792);
   U583 : OAI221_X1 port map( B1 => n611, B2 => n2025, C1 => n1859, C2 => n2018
                           , A => n794, ZN => n1577);
   U584 : AOI222_X1 port map( A1 => n2013, A2 => n38, B1 => n2007, B2 => n613, 
                           C1 => n2001, C2 => n614, ZN => n794);
   U585 : OAI221_X1 port map( B1 => n615, B2 => n2025, C1 => n1858, C2 => n2018
                           , A => n796, ZN => n1575);
   U586 : AOI222_X1 port map( A1 => n2013, A2 => n37, B1 => n2007, B2 => n617, 
                           C1 => n2001, C2 => n618, ZN => n796);
   U587 : OAI221_X1 port map( B1 => n619, B2 => n2024, C1 => n1857, C2 => n2018
                           , A => n798, ZN => n1573);
   U588 : AOI222_X1 port map( A1 => n2012, A2 => n36, B1 => n2006, B2 => n621, 
                           C1 => n2000, C2 => n622, ZN => n798);
   U589 : OAI221_X1 port map( B1 => n2055, B2 => n538, C1 => n1945, C2 => n2045
                           , A => n539, ZN => n1689);
   U590 : AOI222_X1 port map( A1 => n60, A2 => n2039, B1 => n188, B2 => n2034, 
                           C1 => n2032, C2 => n540, ZN => n539);
   U591 : OAI221_X1 port map( B1 => n2055, B2 => n541, C1 => n1944, C2 => n2045
                           , A => n542, ZN => n1688);
   U592 : AOI222_X1 port map( A1 => n59, A2 => n2039, B1 => n187, B2 => n2034, 
                           C1 => n2032, C2 => n543, ZN => n542);
   U593 : OAI221_X1 port map( B1 => n2055, B2 => n544, C1 => n1943, C2 => n2045
                           , A => n545, ZN => n1687);
   U594 : AOI222_X1 port map( A1 => n58, A2 => n2039, B1 => n186, B2 => n2034, 
                           C1 => n2032, C2 => n546, ZN => n545);
   U595 : OAI221_X1 port map( B1 => n2055, B2 => n547, C1 => n1942, C2 => n2045
                           , A => n548, ZN => n1686);
   U596 : AOI222_X1 port map( A1 => n57, A2 => n2039, B1 => n185, B2 => n2034, 
                           C1 => n2032, C2 => n549, ZN => n548);
   U597 : OAI221_X1 port map( B1 => n2055, B2 => n550, C1 => n1941, C2 => n2045
                           , A => n551, ZN => n1685);
   U598 : AOI222_X1 port map( A1 => n56, A2 => n2039, B1 => n184, B2 => n2034, 
                           C1 => n2032, C2 => n552, ZN => n551);
   U599 : OAI221_X1 port map( B1 => n2055, B2 => n553, C1 => n1940, C2 => n2045
                           , A => n554, ZN => n1684);
   U600 : AOI222_X1 port map( A1 => n55, A2 => n2039, B1 => n183, B2 => n2034, 
                           C1 => n2032, C2 => n555, ZN => n554);
   U601 : OAI221_X1 port map( B1 => n2055, B2 => n556, C1 => n1939, C2 => n2045
                           , A => n557, ZN => n1683);
   U602 : AOI222_X1 port map( A1 => n54, A2 => n2039, B1 => n182, B2 => n2034, 
                           C1 => n2032, C2 => n558, ZN => n557);
   U603 : OAI221_X1 port map( B1 => n2055, B2 => n559, C1 => n1938, C2 => n2045
                           , A => n560, ZN => n1682);
   U604 : AOI222_X1 port map( A1 => n53, A2 => n2039, B1 => n181, B2 => n2034, 
                           C1 => n2032, C2 => n561, ZN => n560);
   U605 : OAI221_X1 port map( B1 => n2054, B2 => n583, C1 => n1930, C2 => n2046
                           , A => n584, ZN => n1674);
   U606 : AOI222_X1 port map( A1 => n45, A2 => n2040, B1 => n2035, B2 => n585, 
                           C1 => n2031, C2 => n586, ZN => n584);
   U607 : OAI221_X1 port map( B1 => n2054, B2 => n587, C1 => n1929, C2 => n2046
                           , A => n588, ZN => n1673);
   U608 : AOI222_X1 port map( A1 => n44, A2 => n2040, B1 => n2035, B2 => n589, 
                           C1 => n2031, C2 => n590, ZN => n588);
   U609 : OAI221_X1 port map( B1 => n2054, B2 => n591, C1 => n1928, C2 => n2046
                           , A => n592, ZN => n1672);
   U610 : AOI222_X1 port map( A1 => n43, A2 => n2040, B1 => n2035, B2 => n593, 
                           C1 => n2031, C2 => n594, ZN => n592);
   U611 : OAI221_X1 port map( B1 => n2054, B2 => n595, C1 => n1927, C2 => n2046
                           , A => n596, ZN => n1671);
   U612 : AOI222_X1 port map( A1 => n42, A2 => n2040, B1 => n2035, B2 => n597, 
                           C1 => n2031, C2 => n598, ZN => n596);
   U613 : OAI221_X1 port map( B1 => n2054, B2 => n599, C1 => n1926, C2 => n2046
                           , A => n600, ZN => n1670);
   U614 : AOI222_X1 port map( A1 => n41, A2 => n2040, B1 => n2035, B2 => n601, 
                           C1 => n2031, C2 => n602, ZN => n600);
   U615 : OAI221_X1 port map( B1 => n2054, B2 => n603, C1 => n1925, C2 => n2046
                           , A => n604, ZN => n1669);
   U616 : AOI222_X1 port map( A1 => n40, A2 => n2040, B1 => n2036, B2 => n605, 
                           C1 => n2031, C2 => n606, ZN => n604);
   U617 : OAI221_X1 port map( B1 => n2054, B2 => n607, C1 => n1924, C2 => n2047
                           , A => n608, ZN => n1668);
   U618 : AOI222_X1 port map( A1 => n39, A2 => n2041, B1 => n2036, B2 => n609, 
                           C1 => n2031, C2 => n610, ZN => n608);
   U619 : OAI221_X1 port map( B1 => n2054, B2 => n611, C1 => n1923, C2 => n2047
                           , A => n612, ZN => n1667);
   U620 : AOI222_X1 port map( A1 => n38, A2 => n2041, B1 => n2036, B2 => n613, 
                           C1 => n2031, C2 => n614, ZN => n612);
   U621 : OAI221_X1 port map( B1 => n2054, B2 => n615, C1 => n1922, C2 => n2047
                           , A => n616, ZN => n1666);
   U622 : AOI222_X1 port map( A1 => n37, A2 => n2041, B1 => n2036, B2 => n617, 
                           C1 => n2031, C2 => n618, ZN => n616);
   U623 : INV_X1 port map( A => DATAIN(0), ZN => n743);
   U624 : INV_X1 port map( A => DATAIN(1), ZN => n745);
   U625 : INV_X1 port map( A => DATAIN(2), ZN => n747);
   U626 : INV_X1 port map( A => DATAIN(3), ZN => n749);
   U627 : INV_X1 port map( A => DATAIN(4), ZN => n751);
   U628 : INV_X1 port map( A => DATAIN(5), ZN => n753);
   U629 : INV_X1 port map( A => DATAIN(6), ZN => n755);
   U630 : INV_X1 port map( A => DATAIN(7), ZN => n757);
   U631 : INV_X1 port map( A => DATAIN(8), ZN => n759);
   U632 : INV_X1 port map( A => DATAIN(9), ZN => n761);
   U633 : INV_X1 port map( A => DATAIN(10), ZN => n763);
   U634 : INV_X1 port map( A => DATAIN(11), ZN => n765);
   U635 : INV_X1 port map( A => DATAIN(12), ZN => n767);
   U636 : INV_X1 port map( A => DATAIN(13), ZN => n769);
   U637 : INV_X1 port map( A => DATAIN(14), ZN => n771);
   U638 : INV_X1 port map( A => DATAIN(15), ZN => n773);
   U639 : INV_X1 port map( A => DATAIN(16), ZN => n775);
   U640 : INV_X1 port map( A => DATAIN(17), ZN => n777);
   U641 : INV_X1 port map( A => DATAIN(18), ZN => n779);
   U642 : INV_X1 port map( A => DATAIN(19), ZN => n781);
   U643 : INV_X1 port map( A => DATAIN(20), ZN => n783);
   U644 : INV_X1 port map( A => DATAIN(21), ZN => n785);
   U645 : INV_X1 port map( A => DATAIN(22), ZN => n787);
   U646 : INV_X1 port map( A => DATAIN(23), ZN => n789);
   U647 : INV_X1 port map( A => DATAIN(24), ZN => n791);
   U648 : INV_X1 port map( A => DATAIN(25), ZN => n793);
   U649 : INV_X1 port map( A => DATAIN(26), ZN => n795);
   U650 : INV_X1 port map( A => DATAIN(27), ZN => n797);
   U651 : INV_X1 port map( A => DATAIN(28), ZN => n799);
   U652 : INV_X1 port map( A => DATAIN(29), ZN => n801);
   U653 : INV_X1 port map( A => DATAIN(30), ZN => n803);
   U654 : INV_X1 port map( A => DATAIN(31), ZN => n805);
   U655 : INV_X1 port map( A => DATAIN(32), ZN => n807);
   U656 : INV_X1 port map( A => DATAIN(33), ZN => n809);
   U657 : INV_X1 port map( A => DATAIN(34), ZN => n811);
   U658 : INV_X1 port map( A => DATAIN(35), ZN => n813);
   U659 : INV_X1 port map( A => DATAIN(36), ZN => n815);
   U660 : INV_X1 port map( A => DATAIN(37), ZN => n817);
   U661 : INV_X1 port map( A => DATAIN(38), ZN => n819);
   U662 : INV_X1 port map( A => DATAIN(39), ZN => n821);
   U663 : INV_X1 port map( A => DATAIN(40), ZN => n823);
   U664 : INV_X1 port map( A => DATAIN(41), ZN => n825);
   U665 : INV_X1 port map( A => DATAIN(42), ZN => n827);
   U666 : INV_X1 port map( A => DATAIN(43), ZN => n829);
   U667 : INV_X1 port map( A => DATAIN(44), ZN => n831);
   U668 : INV_X1 port map( A => DATAIN(45), ZN => n833);
   U669 : INV_X1 port map( A => DATAIN(46), ZN => n835);
   U670 : INV_X1 port map( A => DATAIN(47), ZN => n837);
   U671 : INV_X1 port map( A => DATAIN(48), ZN => n839);
   U672 : INV_X1 port map( A => DATAIN(49), ZN => n841);
   U673 : INV_X1 port map( A => DATAIN(50), ZN => n843);
   U674 : INV_X1 port map( A => DATAIN(51), ZN => n845);
   U675 : INV_X1 port map( A => DATAIN(52), ZN => n847);
   U676 : INV_X1 port map( A => DATAIN(53), ZN => n849);
   U677 : INV_X1 port map( A => DATAIN(54), ZN => n851);
   U678 : INV_X1 port map( A => DATAIN(55), ZN => n853);
   U679 : INV_X1 port map( A => DATAIN(56), ZN => n855);
   U680 : INV_X1 port map( A => DATAIN(57), ZN => n857);
   U681 : INV_X1 port map( A => DATAIN(58), ZN => n859);
   U682 : INV_X1 port map( A => DATAIN(59), ZN => n861);
   U683 : INV_X1 port map( A => DATAIN(60), ZN => n863);
   U684 : INV_X1 port map( A => DATAIN(61), ZN => n865);
   U685 : INV_X1 port map( A => DATAIN(62), ZN => n867);
   U686 : INV_X1 port map( A => DATAIN(63), ZN => n871);
   U687 : CLKBUF_X1 port map( A => n979, Z => n1955);
   U688 : CLKBUF_X1 port map( A => n978, Z => n1961);
   U689 : CLKBUF_X1 port map( A => n939, Z => n1967);
   U690 : CLKBUF_X1 port map( A => n938, Z => n1973);
   U691 : CLKBUF_X1 port map( A => n876, Z => n1979);
   U692 : CLKBUF_X1 port map( A => n875, Z => n1985);
   U693 : CLKBUF_X1 port map( A => n742, Z => n1991);
   U694 : CLKBUF_X1 port map( A => n741, Z => n1997);
   U695 : CLKBUF_X1 port map( A => n740, Z => n2003);
   U696 : CLKBUF_X1 port map( A => n739, Z => n2009);
   U697 : CLKBUF_X1 port map( A => n738, Z => n2015);
   U698 : CLKBUF_X1 port map( A => n736, Z => n2021);
   U699 : CLKBUF_X1 port map( A => n735, Z => n2027);
   U700 : CLKBUF_X1 port map( A => n527, Z => n2033);
   U701 : CLKBUF_X1 port map( A => n525, Z => n2044);
   U702 : CLKBUF_X1 port map( A => n523, Z => n2050);
   U703 : CLKBUF_X1 port map( A => n521, Z => n2056);
   U704 : INV_X1 port map( A => ADD_RD2(0), ZN => n2057);
   U705 : INV_X1 port map( A => ADD_RD2(1), ZN => n2058);
   U706 : INV_X1 port map( A => ADD_RD1(0), ZN => n2059);
   U707 : INV_X1 port map( A => ADD_RD1(1), ZN => n2060);
   U708 : INV_X1 port map( A => ADD_WR(0), ZN => n2061);
   U709 : INV_X1 port map( A => ADD_WR(1), ZN => n2062);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4.all;

entity register_file_reg_size64_file_size4_7 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_reg_size64_file_size4_7;

architecture SYN_BEHAVIORAL of register_file_reg_size64_file_size4_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n415, n1200, n1202, n1204, n1310, n1311, n1312, n1313, n1314, n1315
      , n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n871, n872, 
      n873, n875, n876, n936, n938, n939, n975, n978, n979, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176 : std_logic
      ;

begin
   
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => n174,
                           QN => n2028);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => n175,
                           QN => n2027);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => n176,
                           QN => n2026);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => n177,
                           QN => n2025);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => n178,
                           QN => n2024);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => n179,
                           QN => n2023);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => n180,
                           QN => n2022);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => n181,
                           QN => n2021);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => n182,
                           QN => n2020);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => n183, 
                           QN => n2019);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => n184, 
                           QN => n2018);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => n185, 
                           QN => n2017);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => n186, 
                           QN => n2016);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => n187, 
                           QN => n2015);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => n188, 
                           QN => n2014);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => n189, 
                           QN => n2013);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => n190, 
                           QN => n2012);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => n191, 
                           QN => n2011);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => n192, 
                           QN => n2010);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => n65, 
                           QN => n2063);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => n66, 
                           QN => n2062);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n67, 
                           QN => n2061);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => n68, 
                           QN => n2060);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => n69, 
                           QN => n2059);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => n70, 
                           QN => n2058);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => n71, 
                           QN => n2057);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => n72, 
                           QN => n2056);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => n73, 
                           QN => n2055);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => n74, 
                           QN => n2054);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => n75, 
                           QN => n2053);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => n76, 
                           QN => n2052);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => n77, 
                           QN => n2051);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => n78, 
                           QN => n2050);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => n79, 
                           QN => n2049);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => n80, 
                           QN => n2048);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => n81, 
                           QN => n2047);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => n82, 
                           QN => n2046);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => n83, 
                           QN => n2045);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => n84, 
                           QN => n2044);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => n85, 
                           QN => n2043);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => n86, 
                           QN => n2042);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => n87, 
                           QN => n2041);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => n88, 
                           QN => n2040);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => n89, 
                           QN => n2039);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => n90, 
                           QN => n2038);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => n91, 
                           QN => n2037);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => n92, 
                           QN => n2036);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => n93, 
                           QN => n2035);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => n94, 
                           QN => n2034);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => n95, 
                           QN => n2033);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => n96, 
                           QN => n2032);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => n97, 
                           QN => n2031);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => n98, 
                           QN => n2030);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => n99, 
                           QN => n2029);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => n2, 
                           QN => n2009);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => n3, 
                           QN => n2008);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => n4, 
                           QN => n2007);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => n5, 
                           QN => n2006);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => n6, 
                           QN => n2005);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => n7, 
                           QN => n2004);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => n8, 
                           QN => n2003);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => n9, 
                           QN => n2002);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => n13, 
                           QN => n2001);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => n14, 
                           QN => n2000);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => n15, 
                           QN => n1999);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => n16, 
                           QN => n1998);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => n17, 
                           QN => n1997);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => n18, 
                           QN => n1996);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => n19, 
                           QN => n1995);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => n20, 
                           QN => n1994);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => n21, 
                           QN => n1993);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => n22, 
                           QN => n1992);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => n23, 
                           QN => n1991);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => n24, 
                           QN => n1990);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => n25, 
                           QN => n1989);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => n26, 
                           QN => n1988);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n27, 
                           QN => n1987);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => n28, 
                           QN => n1986);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n29, 
                           QN => n1985);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => n30, 
                           QN => n1984);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n31, 
                           QN => n1983);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => n32, 
                           QN => n1982);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n33, 
                           QN => n1981);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => n34, 
                           QN => n1980);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n35, 
                           QN => n1979);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => n36, 
                           QN => n1978);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => n37, 
                           QN => n1977);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => n38, 
                           QN => n1976);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => n39, 
                           QN => n1975);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => n40, 
                           QN => n1974);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => n41, 
                           QN => n1973);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => n42, 
                           QN => n1972);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => n43, 
                           QN => n1971);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => n44, 
                           QN => n1970);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => n45, 
                           QN => n1969);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => n46, 
                           QN => n1968);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => n47, 
                           QN => n1967);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => n48, 
                           QN => n1966);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => n49, 
                           QN => n1965);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => n50, 
                           QN => n1964);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => n51, 
                           QN => n1963);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => n52, 
                           QN => n1962);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => n53, 
                           QN => n1961);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => n54, 
                           QN => n1960);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n55, 
                           QN => n1959);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => n56, 
                           QN => n1958);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n57, 
                           QN => n1957);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => n58, 
                           QN => n1956);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n59, 
                           QN => n1955);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => n60, 
                           QN => n1954);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n61, 
                           QN => n1953);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => n62, 
                           QN => n1952);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n63, 
                           QN => n1951);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => n64, 
                           QN => n1950);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n999,
                           QN => n728);
   OUT2_reg_63_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => OUT2(63), QN
                           => n1822);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n1000
                           , QN => n725);
   OUT2_reg_62_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => OUT2(62), QN
                           => n1823);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n1001
                           , QN => n722);
   OUT2_reg_61_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => OUT2(61), QN
                           => n1824);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n1002
                           , QN => n719);
   OUT2_reg_60_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => OUT2(60), QN
                           => n1825);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n1003
                           , QN => n716);
   OUT2_reg_59_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => OUT2(59), QN
                           => n1826);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n1004
                           , QN => n713);
   OUT2_reg_58_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => OUT2(58), QN
                           => n1827);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n1005
                           , QN => n710);
   OUT2_reg_57_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => OUT2(57), QN
                           => n1828);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n1006
                           , QN => n707);
   OUT2_reg_56_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => OUT2(56), QN
                           => n1829);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n1007
                           , QN => n704);
   OUT2_reg_55_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => OUT2(55), QN
                           => n1830);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n1008
                           , QN => n700);
   OUT2_reg_54_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => OUT2(54), QN
                           => n1831);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n1009
                           , QN => n696);
   OUT2_reg_53_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => OUT2(53), QN
                           => n1832);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n1010
                           , QN => n692);
   OUT2_reg_52_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => OUT2(52), QN
                           => n1833);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n1011
                           , QN => n689);
   OUT2_reg_51_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => OUT2(51), QN
                           => n1834);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n1012
                           , QN => n686);
   OUT2_reg_50_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => OUT2(50), QN
                           => n1835);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n1013
                           , QN => n683);
   OUT2_reg_49_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => OUT2(49), QN
                           => n1836);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n1014
                           , QN => n680);
   OUT2_reg_48_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => OUT2(48), QN
                           => n1837);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n1015
                           , QN => n677);
   OUT2_reg_47_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => OUT2(47), QN
                           => n1838);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n1016
                           , QN => n674);
   OUT2_reg_46_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => OUT2(46), QN
                           => n1839);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n1017
                           , QN => n671);
   OUT2_reg_45_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => OUT2(45), QN
                           => n1840);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n1018
                           , QN => n668);
   OUT2_reg_44_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => OUT2(44), QN
                           => n1841);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n1019
                           , QN => n665);
   OUT2_reg_43_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => OUT2(43), QN
                           => n1842);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n1020
                           , QN => n662);
   OUT2_reg_42_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => OUT2(42), QN
                           => n1843);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n1021
                           , QN => n659);
   OUT2_reg_41_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => OUT2(41), QN
                           => n1844);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n1022
                           , QN => n656);
   OUT2_reg_40_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => OUT2(40), QN
                           => n1845);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n1023
                           , QN => n653);
   OUT2_reg_39_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => OUT2(39), QN
                           => n1846);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n1024
                           , QN => n650);
   OUT2_reg_38_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => OUT2(38), QN
                           => n1847);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n1025
                           , QN => n647);
   OUT2_reg_37_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => OUT2(37), QN
                           => n1848);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n1026
                           , QN => n644);
   OUT2_reg_36_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => OUT2(36), QN
                           => n1849);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n1027
                           , QN => n641);
   OUT2_reg_35_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => OUT2(35), QN
                           => n1850);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n1028
                           , QN => n638);
   OUT2_reg_34_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => OUT2(34), QN
                           => n1851);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n1029
                           , QN => n635);
   OUT2_reg_33_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => OUT2(33), QN
                           => n1852);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n1030
                           , QN => n632);
   OUT2_reg_32_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => OUT2(32), QN
                           => n1853);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n1031
                           , QN => n629);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => OUT2(31), QN
                           => n1854);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n1032
                           , QN => n626);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => OUT2(30), QN
                           => n1855);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n1033
                           , QN => n623);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => OUT2(29), QN
                           => n1856);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n1034
                           , QN => n619);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => OUT2(28), QN
                           => n1857);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n1035
                           , QN => n615);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => OUT2(27), QN
                           => n1858);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n1036
                           , QN => n611);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => OUT2(26), QN
                           => n1859);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n1037
                           , QN => n607);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => OUT2(25), QN
                           => n1860);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n1038
                           , QN => n603);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => OUT2(24), QN
                           => n1861);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n1039
                           , QN => n599);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => OUT2(23), QN
                           => n1862);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n1040
                           , QN => n595);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => OUT2(22), QN
                           => n1863);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n1041
                           , QN => n591);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => OUT2(21), QN
                           => n1864);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n1042
                           , QN => n587);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => OUT2(20), QN
                           => n1865);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n1043
                           , QN => n583);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => OUT2(19), QN
                           => n1866);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n1044
                           , QN => n580);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => OUT2(18), QN
                           => n1867);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n1045
                           , QN => n577);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => OUT2(17), QN
                           => n1868);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n1046
                           , QN => n574);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => OUT2(16), QN
                           => n1869);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n1047
                           , QN => n571);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => OUT2(15), QN
                           => n1870);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n1048
                           , QN => n568);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => OUT2(14), QN
                           => n1871);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n1049
                           , QN => n565);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => OUT2(13), QN
                           => n1872);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n1050
                           , QN => n562);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => OUT2(12), QN
                           => n1873);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n1051
                           , QN => n559);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => OUT2(11), QN
                           => n1874);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n1052
                           , QN => n556);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => OUT2(10), QN
                           => n1875);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n1053,
                           QN => n553);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => OUT2(9), QN 
                           => n1876);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => n1054,
                           QN => n550);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => OUT2(8), QN 
                           => n1877);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => n1055,
                           QN => n547);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => OUT2(7), QN 
                           => n1878);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => n1056,
                           QN => n544);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => OUT2(6), QN 
                           => n1879);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => n1057,
                           QN => n541);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => OUT2(5), QN 
                           => n1880);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => n1058,
                           QN => n538);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => OUT2(4), QN 
                           => n1881);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => n1059,
                           QN => n535);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => OUT2(3), QN 
                           => n1882);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n1060,
                           QN => n532);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => OUT2(2), QN 
                           => n1883);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n1061,
                           QN => n529);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => OUT2(1), QN 
                           => n1884);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n1062,
                           QN => n522);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => OUT2(0), QN 
                           => n1885);
   OUT1_reg_63_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => OUT1(63), QN
                           => n1886);
   OUT1_reg_62_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => OUT1(62), QN
                           => n1887);
   OUT1_reg_61_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => OUT1(61), QN
                           => n1888);
   OUT1_reg_60_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => OUT1(60), QN
                           => n1889);
   OUT1_reg_59_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => OUT1(59), QN
                           => n1890);
   OUT1_reg_58_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => OUT1(58), QN
                           => n1891);
   OUT1_reg_57_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => OUT1(57), QN
                           => n1892);
   OUT1_reg_56_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => OUT1(56), QN
                           => n1893);
   OUT1_reg_55_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => OUT1(55), QN
                           => n1894);
   OUT1_reg_54_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => OUT1(54), QN
                           => n1895);
   OUT1_reg_53_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => OUT1(53), QN
                           => n1896);
   OUT1_reg_52_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => OUT1(52), QN
                           => n1897);
   OUT1_reg_51_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => OUT1(51), QN
                           => n1898);
   OUT1_reg_50_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => OUT1(50), QN
                           => n1899);
   OUT1_reg_49_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => OUT1(49), QN
                           => n1900);
   OUT1_reg_48_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => OUT1(48), QN
                           => n1901);
   OUT1_reg_47_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => OUT1(47), QN
                           => n1902);
   OUT1_reg_46_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => OUT1(46), QN
                           => n1903);
   OUT1_reg_45_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => OUT1(45), QN
                           => n1904);
   OUT1_reg_44_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => OUT1(44), QN
                           => n1905);
   OUT1_reg_43_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => OUT1(43), QN
                           => n1906);
   OUT1_reg_42_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => OUT1(42), QN
                           => n1907);
   OUT1_reg_41_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => OUT1(41), QN
                           => n1908);
   OUT1_reg_40_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => OUT1(40), QN
                           => n1909);
   OUT1_reg_39_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => OUT1(39), QN
                           => n1910);
   OUT1_reg_38_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => OUT1(38), QN
                           => n1911);
   OUT1_reg_37_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => OUT1(37), QN
                           => n1912);
   OUT1_reg_36_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => OUT1(36), QN
                           => n1913);
   OUT1_reg_35_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => OUT1(35), QN
                           => n1914);
   OUT1_reg_34_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => OUT1(34), QN
                           => n1915);
   OUT1_reg_33_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => OUT1(33), QN
                           => n1916);
   OUT1_reg_32_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => OUT1(32), QN
                           => n1917);
   OUT1_reg_31_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => OUT1(31), QN
                           => n1918);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => OUT1(30), QN
                           => n1919);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => OUT1(29), QN
                           => n1920);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => OUT1(28), QN
                           => n1921);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => OUT1(27), QN
                           => n1922);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => OUT1(26), QN
                           => n1923);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => OUT1(25), QN
                           => n1924);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => OUT1(24), QN
                           => n1925);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => OUT1(23), QN
                           => n1926);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => OUT1(22), QN
                           => n1927);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => OUT1(21), QN
                           => n1928);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => OUT1(20), QN
                           => n1929);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => OUT1(19), QN
                           => n1930);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => OUT1(18), QN
                           => n1931);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => OUT1(17), QN
                           => n1932);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => OUT1(16), QN
                           => n1933);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => OUT1(15), QN
                           => n1934);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => OUT1(14), QN
                           => n1935);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => OUT1(13), QN
                           => n1936);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => OUT1(12), QN
                           => n1937);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => OUT1(11), QN
                           => n1938);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => OUT1(10), QN
                           => n1939);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => OUT1(9), QN 
                           => n1940);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => OUT1(8), QN 
                           => n1941);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => OUT1(7), QN 
                           => n1942);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => OUT1(6), QN 
                           => n1943);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => OUT1(5), QN 
                           => n1944);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => OUT1(4), QN 
                           => n1945);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => OUT1(3), QN 
                           => n1946);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => OUT1(2), QN 
                           => n1947);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => OUT1(1), QN 
                           => n1948);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => OUT1(0), QN 
                           => n1949);
   U859 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n2164, A3 => ADD_RD1(1), 
                           ZN => n521);
   U860 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n2135, A3 => ADD_RD2(1), 
                           ZN => n735);
   U861 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n873, A3 => ADD_WR(1), ZN 
                           => n872);
   U862 : NAND3_X1 port map( A1 => n873, A2 => n2175, A3 => ADD_WR(1), ZN => 
                           n936);
   U863 : NAND3_X1 port map( A1 => n873, A2 => n2176, A3 => ADD_WR(0), ZN => 
                           n975);
   U864 : NAND3_X1 port map( A1 => n2175, A2 => n2176, A3 => n873, ZN => n998);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => n537, 
                           QN => n1818);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => n534, 
                           QN => n1819);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => n531, 
                           QN => n1820);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => n528, 
                           QN => n1821);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => n730,
                           QN => n415);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => n702,
                           QN => n1200);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => n698,
                           QN => n1202);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => n694,
                           QN => n1204);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => n622,
                           QN => n1793);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => n618,
                           QN => n1794);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => n614,
                           QN => n1795);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => n610,
                           QN => n1796);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => n606,
                           QN => n1797);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => n602,
                           QN => n1798);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => n598,
                           QN => n1799);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => n594,
                           QN => n1800);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => n590,
                           QN => n1801);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => n586,
                           QN => n1802);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => n582,
                           QN => n1803);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => n579,
                           QN => n1804);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => n576,
                           QN => n1805);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => n573,
                           QN => n1806);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => n570,
                           QN => n1807);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => n567,
                           QN => n1808);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => n564,
                           QN => n1809);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => n561,
                           QN => n1810);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => n558,
                           QN => n1811);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => n555, 
                           QN => n1812);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => n552, 
                           QN => n1813);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => n549, 
                           QN => n1814);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => n546, 
                           QN => n1815);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => n543, 
                           QN => n1816);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => n540, 
                           QN => n1817);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => n731,
                           QN => n1694);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => n727,
                           QN => n1695);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => n724,
                           QN => n1696);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => n721,
                           QN => n1697);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => n718,
                           QN => n1698);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => n715,
                           QN => n1699);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => n712,
                           QN => n1700);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => n709,
                           QN => n1701);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => n706,
                           QN => n1702);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => n703,
                           QN => n1703);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => n699,
                           QN => n1704);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => n695,
                           QN => n1705);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => n691,
                           QN => n1706);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => n688,
                           QN => n1707);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => n685,
                           QN => n1708);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => n682,
                           QN => n1709);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => n679,
                           QN => n1710);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => n676,
                           QN => n1711);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => n673,
                           QN => n1712);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => n670,
                           QN => n1713);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => n667,
                           QN => n1714);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => n664,
                           QN => n1715);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => n661,
                           QN => n1716);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => n658,
                           QN => n1717);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => n655,
                           QN => n1718);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => n652,
                           QN => n1719);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => n649,
                           QN => n1720);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => n646,
                           QN => n1721);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => n643,
                           QN => n1722);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => n640,
                           QN => n1723);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => n637,
                           QN => n1724);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => n634,
                           QN => n1725);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => n631,
                           QN => n1726);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => n628,
                           QN => n1727);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n625,
                           QN => n1728);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => n621,
                           QN => n1729);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => n617,
                           QN => n1730);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => n613,
                           QN => n1731);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => n609,
                           QN => n1732);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => n605,
                           QN => n1733);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => n601,
                           QN => n1734);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => n597,
                           QN => n1735);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => n593,
                           QN => n1736);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => n589,
                           QN => n1737);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => n585,
                           QN => n1738);
   U3 : BUF_X1 port map( A => n521, Z => n2167);
   U4 : BUF_X1 port map( A => n521, Z => n2166);
   U5 : BUF_X1 port map( A => n521, Z => n2165);
   U6 : BUF_X1 port map( A => n735, Z => n2139);
   U7 : BUF_X1 port map( A => n735, Z => n2138);
   U8 : BUF_X1 port map( A => n735, Z => n2137);
   U9 : BUF_X1 port map( A => n735, Z => n2136);
   U10 : BUF_X1 port map( A => n521, Z => n2169);
   U11 : BUF_X1 port map( A => n521, Z => n2168);
   U12 : BUF_X1 port map( A => n735, Z => n2140);
   U13 : BUF_X1 port map( A => n526, Z => n2151);
   U14 : BUF_X1 port map( A => n526, Z => n2152);
   U15 : BUF_X1 port map( A => n527, Z => n2144);
   U16 : BUF_X1 port map( A => n527, Z => n2146);
   U17 : BUF_X1 port map( A => n527, Z => n2145);
   U18 : BUF_X1 port map( A => n523, Z => n2159);
   U19 : BUF_X1 port map( A => n523, Z => n2160);
   U20 : BUF_X1 port map( A => n523, Z => n2161);
   U21 : BUF_X1 port map( A => n523, Z => n2162);
   U22 : BUF_X1 port map( A => n523, Z => n2163);
   U23 : BUF_X1 port map( A => n736, Z => n2130);
   U24 : BUF_X1 port map( A => n736, Z => n2131);
   U25 : BUF_X1 port map( A => n736, Z => n2132);
   U26 : BUF_X1 port map( A => n736, Z => n2133);
   U27 : BUF_X1 port map( A => n736, Z => n2134);
   U28 : BUF_X1 port map( A => n525, Z => n2154);
   U29 : BUF_X1 port map( A => n525, Z => n2155);
   U30 : BUF_X1 port map( A => n525, Z => n2156);
   U31 : BUF_X1 port map( A => n525, Z => n2157);
   U32 : BUF_X1 port map( A => n738, Z => n2128);
   U33 : BUF_X1 port map( A => n738, Z => n2127);
   U34 : BUF_X1 port map( A => n738, Z => n2126);
   U35 : BUF_X1 port map( A => n738, Z => n2125);
   U36 : BUF_X1 port map( A => n738, Z => n2124);
   U37 : BUF_X1 port map( A => n742, Z => n2104);
   U38 : BUF_X1 port map( A => n742, Z => n2103);
   U39 : BUF_X1 port map( A => n742, Z => n2102);
   U40 : BUF_X1 port map( A => n742, Z => n2101);
   U41 : BUF_X1 port map( A => n739, Z => n2122);
   U42 : BUF_X1 port map( A => n739, Z => n2121);
   U43 : BUF_X1 port map( A => n739, Z => n2120);
   U44 : BUF_X1 port map( A => n739, Z => n2119);
   U45 : BUF_X1 port map( A => n739, Z => n2118);
   U46 : BUF_X1 port map( A => n740, Z => n2116);
   U47 : BUF_X1 port map( A => n740, Z => n2115);
   U48 : BUF_X1 port map( A => n740, Z => n2114);
   U49 : BUF_X1 port map( A => n740, Z => n2113);
   U50 : BUF_X1 port map( A => n740, Z => n2112);
   U51 : BUF_X1 port map( A => n741, Z => n2106);
   U52 : BUF_X1 port map( A => n875, Z => n2094);
   U53 : BUF_X1 port map( A => n938, Z => n2082);
   U54 : BUF_X1 port map( A => n978, Z => n2070);
   U55 : BUF_X1 port map( A => n741, Z => n2110);
   U56 : BUF_X1 port map( A => n741, Z => n2109);
   U57 : BUF_X1 port map( A => n741, Z => n2108);
   U58 : BUF_X1 port map( A => n741, Z => n2107);
   U59 : BUF_X1 port map( A => n875, Z => n2098);
   U60 : BUF_X1 port map( A => n875, Z => n2097);
   U61 : BUF_X1 port map( A => n875, Z => n2096);
   U62 : BUF_X1 port map( A => n875, Z => n2095);
   U63 : BUF_X1 port map( A => n938, Z => n2086);
   U64 : BUF_X1 port map( A => n938, Z => n2085);
   U65 : BUF_X1 port map( A => n938, Z => n2084);
   U66 : BUF_X1 port map( A => n938, Z => n2083);
   U67 : BUF_X1 port map( A => n978, Z => n2074);
   U68 : BUF_X1 port map( A => n978, Z => n2073);
   U69 : BUF_X1 port map( A => n978, Z => n2072);
   U70 : BUF_X1 port map( A => n978, Z => n2071);
   U71 : BUF_X1 port map( A => n526, Z => n2148);
   U72 : BUF_X1 port map( A => n526, Z => n2150);
   U73 : BUF_X1 port map( A => n876, Z => n2092);
   U74 : BUF_X1 port map( A => n876, Z => n2091);
   U75 : BUF_X1 port map( A => n876, Z => n2090);
   U76 : BUF_X1 port map( A => n876, Z => n2089);
   U77 : BUF_X1 port map( A => n876, Z => n2088);
   U78 : BUF_X1 port map( A => n939, Z => n2080);
   U79 : BUF_X1 port map( A => n939, Z => n2079);
   U80 : BUF_X1 port map( A => n939, Z => n2078);
   U81 : BUF_X1 port map( A => n939, Z => n2077);
   U82 : BUF_X1 port map( A => n939, Z => n2076);
   U83 : BUF_X1 port map( A => n979, Z => n2068);
   U84 : BUF_X1 port map( A => n979, Z => n2067);
   U85 : BUF_X1 port map( A => n979, Z => n2066);
   U86 : BUF_X1 port map( A => n979, Z => n2065);
   U87 : BUF_X1 port map( A => n979, Z => n2064);
   U88 : BUF_X1 port map( A => n527, Z => n2143);
   U89 : BUF_X1 port map( A => n527, Z => n2142);
   U90 : BUF_X1 port map( A => n526, Z => n2149);
   U91 : BUF_X1 port map( A => n525, Z => n2153);
   U92 : BUF_X1 port map( A => n742, Z => n2100);
   U93 : NAND2_X1 port map( A1 => n734, A2 => n872, ZN => n741);
   U94 : NAND2_X1 port map( A1 => n734, A2 => n936, ZN => n875);
   U95 : NAND2_X1 port map( A1 => n734, A2 => n2094, ZN => n876);
   U96 : NAND2_X1 port map( A1 => n734, A2 => n975, ZN => n938);
   U97 : NAND2_X1 port map( A1 => n734, A2 => n2082, ZN => n939);
   U98 : NAND2_X1 port map( A1 => n734, A2 => n998, ZN => n978);
   U99 : NAND2_X1 port map( A1 => n734, A2 => n2070, ZN => n979);
   U100 : OAI22_X1 port map( A1 => n538, A2 => n2111, B1 => n2104, B2 => n751, 
                           ZN => n1620);
   U101 : OAI22_X1 port map( A1 => n541, A2 => n2110, B1 => n2104, B2 => n753, 
                           ZN => n1618);
   U102 : OAI22_X1 port map( A1 => n544, A2 => n2110, B1 => n2104, B2 => n755, 
                           ZN => n1616);
   U103 : OAI22_X1 port map( A1 => n547, A2 => n2110, B1 => n2104, B2 => n757, 
                           ZN => n1614);
   U104 : OAI22_X1 port map( A1 => n550, A2 => n2110, B1 => n2104, B2 => n759, 
                           ZN => n1612);
   U105 : OAI22_X1 port map( A1 => n553, A2 => n2110, B1 => n2104, B2 => n761, 
                           ZN => n1610);
   U106 : OAI22_X1 port map( A1 => n556, A2 => n2110, B1 => n2104, B2 => n763, 
                           ZN => n1608);
   U107 : OAI22_X1 port map( A1 => n559, A2 => n2110, B1 => n2104, B2 => n765, 
                           ZN => n1606);
   U108 : OAI22_X1 port map( A1 => n562, A2 => n2110, B1 => n2104, B2 => n767, 
                           ZN => n1604);
   U109 : OAI22_X1 port map( A1 => n565, A2 => n2110, B1 => n2104, B2 => n769, 
                           ZN => n1602);
   U110 : OAI22_X1 port map( A1 => n568, A2 => n2110, B1 => n2104, B2 => n771, 
                           ZN => n1600);
   U111 : OAI22_X1 port map( A1 => n571, A2 => n2110, B1 => n2104, B2 => n773, 
                           ZN => n1598);
   U112 : OAI22_X1 port map( A1 => n574, A2 => n2110, B1 => n2103, B2 => n775, 
                           ZN => n1596);
   U113 : OAI22_X1 port map( A1 => n577, A2 => n2109, B1 => n2103, B2 => n777, 
                           ZN => n1594);
   U114 : OAI22_X1 port map( A1 => n580, A2 => n2109, B1 => n2103, B2 => n779, 
                           ZN => n1592);
   U115 : OAI22_X1 port map( A1 => n583, A2 => n2109, B1 => n2103, B2 => n781, 
                           ZN => n1590);
   U116 : OAI22_X1 port map( A1 => n587, A2 => n2109, B1 => n2103, B2 => n783, 
                           ZN => n1588);
   U117 : OAI22_X1 port map( A1 => n591, A2 => n2109, B1 => n2103, B2 => n785, 
                           ZN => n1586);
   U118 : OAI22_X1 port map( A1 => n595, A2 => n2109, B1 => n2103, B2 => n787, 
                           ZN => n1584);
   U119 : OAI22_X1 port map( A1 => n599, A2 => n2109, B1 => n2103, B2 => n789, 
                           ZN => n1582);
   U120 : OAI22_X1 port map( A1 => n603, A2 => n2109, B1 => n2103, B2 => n791, 
                           ZN => n1580);
   U121 : OAI22_X1 port map( A1 => n607, A2 => n2109, B1 => n2103, B2 => n793, 
                           ZN => n1578);
   U122 : OAI22_X1 port map( A1 => n611, A2 => n2109, B1 => n2103, B2 => n795, 
                           ZN => n1576);
   U123 : OAI22_X1 port map( A1 => n615, A2 => n2109, B1 => n2103, B2 => n797, 
                           ZN => n1574);
   U124 : OAI22_X1 port map( A1 => n619, A2 => n2109, B1 => n2102, B2 => n799, 
                           ZN => n1572);
   U125 : OAI22_X1 port map( A1 => n623, A2 => n2108, B1 => n2102, B2 => n801, 
                           ZN => n1570);
   U126 : OAI22_X1 port map( A1 => n626, A2 => n2108, B1 => n2102, B2 => n803, 
                           ZN => n1568);
   U127 : OAI22_X1 port map( A1 => n629, A2 => n2108, B1 => n2102, B2 => n805, 
                           ZN => n1566);
   U128 : OAI22_X1 port map( A1 => n632, A2 => n2108, B1 => n2102, B2 => n807, 
                           ZN => n1564);
   U129 : OAI22_X1 port map( A1 => n635, A2 => n2108, B1 => n2102, B2 => n809, 
                           ZN => n1562);
   U130 : OAI22_X1 port map( A1 => n638, A2 => n2108, B1 => n2102, B2 => n811, 
                           ZN => n1560);
   U131 : OAI22_X1 port map( A1 => n641, A2 => n2108, B1 => n2102, B2 => n813, 
                           ZN => n1558);
   U132 : OAI22_X1 port map( A1 => n644, A2 => n2108, B1 => n2102, B2 => n815, 
                           ZN => n1556);
   U133 : OAI22_X1 port map( A1 => n647, A2 => n2108, B1 => n2102, B2 => n817, 
                           ZN => n1554);
   U134 : OAI22_X1 port map( A1 => n650, A2 => n2108, B1 => n2102, B2 => n819, 
                           ZN => n1552);
   U135 : OAI22_X1 port map( A1 => n653, A2 => n2108, B1 => n2102, B2 => n821, 
                           ZN => n1550);
   U136 : OAI22_X1 port map( A1 => n656, A2 => n2108, B1 => n2101, B2 => n823, 
                           ZN => n1548);
   U137 : OAI22_X1 port map( A1 => n659, A2 => n2107, B1 => n2101, B2 => n825, 
                           ZN => n1546);
   U138 : OAI22_X1 port map( A1 => n662, A2 => n2107, B1 => n2101, B2 => n827, 
                           ZN => n1544);
   U139 : OAI22_X1 port map( A1 => n665, A2 => n2107, B1 => n2101, B2 => n829, 
                           ZN => n1542);
   U140 : OAI22_X1 port map( A1 => n668, A2 => n2107, B1 => n2101, B2 => n831, 
                           ZN => n1540);
   U141 : OAI22_X1 port map( A1 => n671, A2 => n2107, B1 => n2101, B2 => n833, 
                           ZN => n1538);
   U142 : OAI22_X1 port map( A1 => n674, A2 => n2107, B1 => n2101, B2 => n835, 
                           ZN => n1536);
   U143 : OAI22_X1 port map( A1 => n677, A2 => n2107, B1 => n2101, B2 => n837, 
                           ZN => n1534);
   U144 : OAI22_X1 port map( A1 => n680, A2 => n2107, B1 => n2101, B2 => n839, 
                           ZN => n1532);
   U145 : OAI22_X1 port map( A1 => n683, A2 => n2107, B1 => n2101, B2 => n841, 
                           ZN => n1530);
   U146 : OAI22_X1 port map( A1 => n686, A2 => n2107, B1 => n2101, B2 => n843, 
                           ZN => n1528);
   U147 : OAI22_X1 port map( A1 => n689, A2 => n2107, B1 => n2101, B2 => n845, 
                           ZN => n1526);
   U148 : OAI22_X1 port map( A1 => n522, A2 => n2111, B1 => n2105, B2 => n743, 
                           ZN => n1628);
   U149 : OAI22_X1 port map( A1 => n529, A2 => n2111, B1 => n2105, B2 => n745, 
                           ZN => n1626);
   U150 : OAI22_X1 port map( A1 => n532, A2 => n2111, B1 => n2105, B2 => n747, 
                           ZN => n1624);
   U151 : OAI22_X1 port map( A1 => n535, A2 => n2111, B1 => n2105, B2 => n749, 
                           ZN => n1622);
   U152 : OAI22_X1 port map( A1 => n692, A2 => n2107, B1 => n2100, B2 => n847, 
                           ZN => n1524);
   U153 : OAI22_X1 port map( A1 => n696, A2 => n2106, B1 => n2100, B2 => n849, 
                           ZN => n1522);
   U154 : OAI22_X1 port map( A1 => n700, A2 => n2106, B1 => n2100, B2 => n851, 
                           ZN => n1520);
   U155 : OAI22_X1 port map( A1 => n704, A2 => n2106, B1 => n2100, B2 => n853, 
                           ZN => n1518);
   U156 : OAI22_X1 port map( A1 => n707, A2 => n2106, B1 => n2100, B2 => n855, 
                           ZN => n1516);
   U157 : OAI22_X1 port map( A1 => n710, A2 => n2106, B1 => n2100, B2 => n857, 
                           ZN => n1514);
   U158 : OAI22_X1 port map( A1 => n713, A2 => n2106, B1 => n2100, B2 => n859, 
                           ZN => n1512);
   U159 : OAI22_X1 port map( A1 => n716, A2 => n2106, B1 => n2100, B2 => n861, 
                           ZN => n1510);
   U160 : OAI22_X1 port map( A1 => n719, A2 => n2106, B1 => n2100, B2 => n863, 
                           ZN => n1508);
   U161 : OAI22_X1 port map( A1 => n722, A2 => n2106, B1 => n2100, B2 => n865, 
                           ZN => n1506);
   U162 : OAI22_X1 port map( A1 => n725, A2 => n2106, B1 => n2100, B2 => n867, 
                           ZN => n1504);
   U163 : OAI22_X1 port map( A1 => n728, A2 => n2106, B1 => n2100, B2 => n871, 
                           ZN => n1502);
   U164 : AND3_X1 port map( A1 => n2173, A2 => n2174, A3 => n2164, ZN => n526);
   U165 : AND3_X1 port map( A1 => n2164, A2 => n2174, A3 => ADD_RD1(0), ZN => 
                           n527);
   U166 : AND3_X1 port map( A1 => n2164, A2 => n2173, A3 => ADD_RD1(1), ZN => 
                           n525);
   U167 : NAND2_X1 port map( A1 => n734, A2 => n2106, ZN => n742);
   U168 : AND3_X1 port map( A1 => n2135, A2 => n2172, A3 => ADD_RD2(0), ZN => 
                           n740);
   U169 : AND3_X1 port map( A1 => n2135, A2 => n2171, A3 => ADD_RD2(1), ZN => 
                           n738);
   U170 : AND3_X1 port map( A1 => n2171, A2 => n2172, A3 => n2135, ZN => n739);
   U171 : AND2_X1 port map( A1 => RD1, A2 => n734, ZN => n523);
   U172 : AND2_X1 port map( A1 => RD2, A2 => n734, ZN => n736);
   U173 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n873);
   U174 : OAI221_X1 port map( B1 => n2169, B2 => n562, C1 => n1937, C2 => n2160
                           , A => n563, ZN => n1681);
   U175 : AOI222_X1 port map( A1 => n52, A2 => n2153, B1 => n180, B2 => n2149, 
                           C1 => n2146, C2 => n564, ZN => n563);
   U176 : OAI221_X1 port map( B1 => n2169, B2 => n565, C1 => n1936, C2 => n2160
                           , A => n566, ZN => n1680);
   U177 : AOI222_X1 port map( A1 => n51, A2 => n2154, B1 => n179, B2 => n2149, 
                           C1 => n2146, C2 => n567, ZN => n566);
   U178 : OAI221_X1 port map( B1 => n2169, B2 => n568, C1 => n1935, C2 => n2160
                           , A => n569, ZN => n1679);
   U179 : AOI222_X1 port map( A1 => n50, A2 => n2154, B1 => n178, B2 => n2149, 
                           C1 => n2146, C2 => n570, ZN => n569);
   U180 : OAI221_X1 port map( B1 => n2169, B2 => n571, C1 => n1934, C2 => n2161
                           , A => n572, ZN => n1678);
   U181 : AOI222_X1 port map( A1 => n49, A2 => n2154, B1 => n177, B2 => n2149, 
                           C1 => n2145, C2 => n573, ZN => n572);
   U182 : OAI221_X1 port map( B1 => n2168, B2 => n574, C1 => n1933, C2 => n2160
                           , A => n575, ZN => n1677);
   U183 : AOI222_X1 port map( A1 => n48, A2 => n2154, B1 => n176, B2 => n2149, 
                           C1 => n2145, C2 => n576, ZN => n575);
   U184 : OAI221_X1 port map( B1 => n2168, B2 => n577, C1 => n1932, C2 => n2160
                           , A => n578, ZN => n1676);
   U185 : AOI222_X1 port map( A1 => n47, A2 => n2154, B1 => n175, B2 => n2149, 
                           C1 => n2145, C2 => n579, ZN => n578);
   U186 : OAI221_X1 port map( B1 => n2168, B2 => n580, C1 => n1931, C2 => n2160
                           , A => n581, ZN => n1675);
   U187 : AOI222_X1 port map( A1 => n46, A2 => n2154, B1 => n174, B2 => n2149, 
                           C1 => n2145, C2 => n582, ZN => n581);
   U188 : OAI221_X1 port map( B1 => n538, B2 => n2140, C1 => n1881, C2 => n2130
                           , A => n750, ZN => n1621);
   U189 : AOI222_X1 port map( A1 => n2128, A2 => n60, B1 => n2122, B2 => n188, 
                           C1 => n2116, C2 => n540, ZN => n750);
   U190 : OAI221_X1 port map( B1 => n541, B2 => n2140, C1 => n1880, C2 => n2130
                           , A => n752, ZN => n1619);
   U191 : AOI222_X1 port map( A1 => n2128, A2 => n59, B1 => n2122, B2 => n187, 
                           C1 => n2116, C2 => n543, ZN => n752);
   U192 : OAI221_X1 port map( B1 => n544, B2 => n2140, C1 => n1879, C2 => n2130
                           , A => n754, ZN => n1617);
   U193 : AOI222_X1 port map( A1 => n2128, A2 => n58, B1 => n2122, B2 => n186, 
                           C1 => n2116, C2 => n546, ZN => n754);
   U194 : OAI221_X1 port map( B1 => n547, B2 => n2140, C1 => n1878, C2 => n2130
                           , A => n756, ZN => n1615);
   U195 : AOI222_X1 port map( A1 => n2128, A2 => n57, B1 => n2122, B2 => n185, 
                           C1 => n2116, C2 => n549, ZN => n756);
   U196 : OAI221_X1 port map( B1 => n550, B2 => n2140, C1 => n1877, C2 => n2130
                           , A => n758, ZN => n1613);
   U197 : AOI222_X1 port map( A1 => n2128, A2 => n56, B1 => n2122, B2 => n184, 
                           C1 => n2116, C2 => n552, ZN => n758);
   U198 : OAI221_X1 port map( B1 => n553, B2 => n2140, C1 => n1876, C2 => n2130
                           , A => n760, ZN => n1611);
   U199 : AOI222_X1 port map( A1 => n2128, A2 => n55, B1 => n2122, B2 => n183, 
                           C1 => n2116, C2 => n555, ZN => n760);
   U200 : OAI221_X1 port map( B1 => n556, B2 => n2140, C1 => n1875, C2 => n2130
                           , A => n762, ZN => n1609);
   U201 : AOI222_X1 port map( A1 => n2128, A2 => n54, B1 => n2122, B2 => n182, 
                           C1 => n2116, C2 => n558, ZN => n762);
   U202 : OAI221_X1 port map( B1 => n559, B2 => n2140, C1 => n1874, C2 => n2130
                           , A => n764, ZN => n1607);
   U203 : AOI222_X1 port map( A1 => n2128, A2 => n53, B1 => n2122, B2 => n181, 
                           C1 => n2116, C2 => n561, ZN => n764);
   U204 : OAI221_X1 port map( B1 => n562, B2 => n2140, C1 => n1873, C2 => n2131
                           , A => n766, ZN => n1605);
   U205 : AOI222_X1 port map( A1 => n2128, A2 => n52, B1 => n2122, B2 => n180, 
                           C1 => n2116, C2 => n564, ZN => n766);
   U206 : OAI221_X1 port map( B1 => n565, B2 => n2140, C1 => n1872, C2 => n2131
                           , A => n768, ZN => n1603);
   U207 : AOI222_X1 port map( A1 => n2128, A2 => n51, B1 => n2122, B2 => n179, 
                           C1 => n2116, C2 => n567, ZN => n768);
   U208 : OAI221_X1 port map( B1 => n568, B2 => n2140, C1 => n1871, C2 => n2131
                           , A => n770, ZN => n1601);
   U209 : AOI222_X1 port map( A1 => n2128, A2 => n50, B1 => n2122, B2 => n178, 
                           C1 => n2116, C2 => n570, ZN => n770);
   U210 : OAI221_X1 port map( B1 => n571, B2 => n2140, C1 => n1870, C2 => n2132
                           , A => n772, ZN => n1599);
   U211 : AOI222_X1 port map( A1 => n2128, A2 => n49, B1 => n2122, B2 => n177, 
                           C1 => n2116, C2 => n573, ZN => n772);
   U212 : OAI221_X1 port map( B1 => n574, B2 => n2139, C1 => n1869, C2 => n2131
                           , A => n774, ZN => n1597);
   U213 : AOI222_X1 port map( A1 => n2127, A2 => n48, B1 => n2121, B2 => n176, 
                           C1 => n2115, C2 => n576, ZN => n774);
   U214 : OAI221_X1 port map( B1 => n577, B2 => n2139, C1 => n1868, C2 => n2131
                           , A => n776, ZN => n1595);
   U215 : AOI222_X1 port map( A1 => n2127, A2 => n47, B1 => n2121, B2 => n175, 
                           C1 => n2115, C2 => n579, ZN => n776);
   U216 : OAI221_X1 port map( B1 => n580, B2 => n2139, C1 => n1867, C2 => n2131
                           , A => n778, ZN => n1593);
   U217 : AOI222_X1 port map( A1 => n2127, A2 => n46, B1 => n2121, B2 => n174, 
                           C1 => n2115, C2 => n582, ZN => n778);
   U218 : OAI221_X1 port map( B1 => n2166, B2 => n656, C1 => n1909, C2 => n2162
                           , A => n657, ZN => n1653);
   U219 : AOI222_X1 port map( A1 => n24, A2 => n2156, B1 => n2151, B2 => n658, 
                           C1 => n88, C2 => n2143, ZN => n657);
   U220 : OAI221_X1 port map( B1 => n2166, B2 => n659, C1 => n1908, C2 => n2162
                           , A => n660, ZN => n1652);
   U221 : AOI222_X1 port map( A1 => n23, A2 => n2156, B1 => n2151, B2 => n661, 
                           C1 => n87, C2 => n2143, ZN => n660);
   U222 : OAI221_X1 port map( B1 => n2166, B2 => n662, C1 => n1907, C2 => n2162
                           , A => n663, ZN => n1651);
   U223 : AOI222_X1 port map( A1 => n22, A2 => n2156, B1 => n2151, B2 => n664, 
                           C1 => n86, C2 => n2143, ZN => n663);
   U224 : OAI221_X1 port map( B1 => n2166, B2 => n665, C1 => n1906, C2 => n2162
                           , A => n666, ZN => n1650);
   U225 : AOI222_X1 port map( A1 => n21, A2 => n2156, B1 => n2151, B2 => n667, 
                           C1 => n85, C2 => n2143, ZN => n666);
   U226 : OAI221_X1 port map( B1 => n2166, B2 => n668, C1 => n1905, C2 => n2162
                           , A => n669, ZN => n1649);
   U227 : AOI222_X1 port map( A1 => n20, A2 => n2156, B1 => n2151, B2 => n670, 
                           C1 => n84, C2 => n2143, ZN => n669);
   U228 : OAI221_X1 port map( B1 => n2166, B2 => n671, C1 => n1904, C2 => n2162
                           , A => n672, ZN => n1648);
   U229 : AOI222_X1 port map( A1 => n19, A2 => n2156, B1 => n2151, B2 => n673, 
                           C1 => n83, C2 => n2143, ZN => n672);
   U230 : OAI221_X1 port map( B1 => n2166, B2 => n674, C1 => n1903, C2 => n2162
                           , A => n675, ZN => n1647);
   U231 : AOI222_X1 port map( A1 => n18, A2 => n2156, B1 => n2151, B2 => n676, 
                           C1 => n82, C2 => n2143, ZN => n675);
   U232 : OAI221_X1 port map( B1 => n2166, B2 => n677, C1 => n1902, C2 => n2162
                           , A => n678, ZN => n1646);
   U233 : AOI222_X1 port map( A1 => n17, A2 => n2156, B1 => n2151, B2 => n679, 
                           C1 => n81, C2 => n2143, ZN => n678);
   U234 : OAI221_X1 port map( B1 => n2166, B2 => n680, C1 => n1901, C2 => n2163
                           , A => n681, ZN => n1645);
   U235 : AOI222_X1 port map( A1 => n16, A2 => n2157, B1 => n2151, B2 => n682, 
                           C1 => n80, C2 => n2143, ZN => n681);
   U236 : OAI221_X1 port map( B1 => n2166, B2 => n683, C1 => n1900, C2 => n2163
                           , A => n684, ZN => n1644);
   U237 : AOI222_X1 port map( A1 => n15, A2 => n2157, B1 => n2151, B2 => n685, 
                           C1 => n79, C2 => n2143, ZN => n684);
   U238 : OAI221_X1 port map( B1 => n2166, B2 => n686, C1 => n1899, C2 => n2163
                           , A => n687, ZN => n1643);
   U239 : AOI222_X1 port map( A1 => n14, A2 => n2157, B1 => n2152, B2 => n688, 
                           C1 => n78, C2 => n2143, ZN => n687);
   U240 : OAI221_X1 port map( B1 => n2166, B2 => n689, C1 => n1898, C2 => n2163
                           , A => n690, ZN => n1642);
   U241 : AOI222_X1 port map( A1 => n13, A2 => n2157, B1 => n2152, B2 => n691, 
                           C1 => n77, C2 => n2143, ZN => n690);
   U242 : OAI221_X1 port map( B1 => n2165, B2 => n692, C1 => n1897, C2 => n2163
                           , A => n693, ZN => n1641);
   U243 : AOI222_X1 port map( A1 => n2158, A2 => n694, B1 => n2152, B2 => n695,
                           C1 => n76, C2 => n2142, ZN => n693);
   U244 : OAI221_X1 port map( B1 => n2165, B2 => n696, C1 => n1896, C2 => n2163
                           , A => n697, ZN => n1640);
   U245 : AOI222_X1 port map( A1 => n2158, A2 => n698, B1 => n2152, B2 => n699,
                           C1 => n75, C2 => n2142, ZN => n697);
   U246 : OAI221_X1 port map( B1 => n2165, B2 => n700, C1 => n1895, C2 => n2163
                           , A => n701, ZN => n1639);
   U247 : AOI222_X1 port map( A1 => n2158, A2 => n702, B1 => n2152, B2 => n703,
                           C1 => n74, C2 => n2142, ZN => n701);
   U248 : OAI221_X1 port map( B1 => n2165, B2 => n704, C1 => n1894, C2 => n2163
                           , A => n705, ZN => n1638);
   U249 : AOI222_X1 port map( A1 => n9, A2 => n2157, B1 => n2152, B2 => n706, 
                           C1 => n73, C2 => n2142, ZN => n705);
   U250 : OAI221_X1 port map( B1 => n2165, B2 => n707, C1 => n1893, C2 => n2163
                           , A => n708, ZN => n1637);
   U251 : AOI222_X1 port map( A1 => n8, A2 => n2157, B1 => n2152, B2 => n709, 
                           C1 => n72, C2 => n2142, ZN => n708);
   U252 : OAI221_X1 port map( B1 => n2165, B2 => n710, C1 => n1892, C2 => n2163
                           , A => n711, ZN => n1636);
   U253 : AOI222_X1 port map( A1 => n7, A2 => n2157, B1 => n2152, B2 => n712, 
                           C1 => n71, C2 => n2142, ZN => n711);
   U254 : OAI221_X1 port map( B1 => n2165, B2 => n713, C1 => n1891, C2 => n2163
                           , A => n714, ZN => n1635);
   U255 : AOI222_X1 port map( A1 => n6, A2 => n2157, B1 => n2152, B2 => n715, 
                           C1 => n70, C2 => n2142, ZN => n714);
   U256 : OAI221_X1 port map( B1 => n2165, B2 => n719, C1 => n1889, C2 => n2163
                           , A => n720, ZN => n1633);
   U257 : AOI222_X1 port map( A1 => n4, A2 => n2157, B1 => n2152, B2 => n721, 
                           C1 => n68, C2 => n2142, ZN => n720);
   U258 : OAI221_X1 port map( B1 => n2165, B2 => n728, C1 => n1886, C2 => n2164
                           , A => n729, ZN => n1630);
   U259 : AOI222_X1 port map( A1 => n2158, A2 => n730, B1 => n2148, B2 => n731,
                           C1 => n65, C2 => n2142, ZN => n729);
   U260 : OAI221_X1 port map( B1 => n623, B2 => n2138, C1 => n1856, C2 => n2132
                           , A => n800, ZN => n1571);
   U261 : AOI222_X1 port map( A1 => n2126, A2 => n35, B1 => n2120, B2 => n625, 
                           C1 => n2114, C2 => n99, ZN => n800);
   U262 : OAI221_X1 port map( B1 => n626, B2 => n2138, C1 => n1855, C2 => n2132
                           , A => n802, ZN => n1569);
   U263 : AOI222_X1 port map( A1 => n2126, A2 => n34, B1 => n2120, B2 => n628, 
                           C1 => n2114, C2 => n98, ZN => n802);
   U264 : OAI221_X1 port map( B1 => n629, B2 => n2138, C1 => n1854, C2 => n2132
                           , A => n804, ZN => n1567);
   U265 : AOI222_X1 port map( A1 => n2126, A2 => n33, B1 => n2120, B2 => n631, 
                           C1 => n2114, C2 => n97, ZN => n804);
   U266 : OAI221_X1 port map( B1 => n632, B2 => n2138, C1 => n1853, C2 => n2132
                           , A => n806, ZN => n1565);
   U267 : AOI222_X1 port map( A1 => n2126, A2 => n32, B1 => n2120, B2 => n634, 
                           C1 => n2114, C2 => n96, ZN => n806);
   U268 : OAI221_X1 port map( B1 => n635, B2 => n2138, C1 => n1852, C2 => n2132
                           , A => n808, ZN => n1563);
   U269 : AOI222_X1 port map( A1 => n2126, A2 => n31, B1 => n2120, B2 => n637, 
                           C1 => n2114, C2 => n95, ZN => n808);
   U270 : OAI221_X1 port map( B1 => n638, B2 => n2138, C1 => n1851, C2 => n2132
                           , A => n810, ZN => n1561);
   U271 : AOI222_X1 port map( A1 => n2126, A2 => n30, B1 => n2120, B2 => n640, 
                           C1 => n2114, C2 => n94, ZN => n810);
   U272 : OAI221_X1 port map( B1 => n641, B2 => n2138, C1 => n1850, C2 => n2132
                           , A => n812, ZN => n1559);
   U273 : AOI222_X1 port map( A1 => n2126, A2 => n29, B1 => n2120, B2 => n643, 
                           C1 => n2114, C2 => n93, ZN => n812);
   U274 : OAI221_X1 port map( B1 => n644, B2 => n2138, C1 => n1849, C2 => n2133
                           , A => n814, ZN => n1557);
   U275 : AOI222_X1 port map( A1 => n2126, A2 => n28, B1 => n2120, B2 => n646, 
                           C1 => n2114, C2 => n92, ZN => n814);
   U276 : OAI221_X1 port map( B1 => n647, B2 => n2138, C1 => n1848, C2 => n2133
                           , A => n816, ZN => n1555);
   U277 : AOI222_X1 port map( A1 => n2126, A2 => n27, B1 => n2120, B2 => n649, 
                           C1 => n2114, C2 => n91, ZN => n816);
   U278 : OAI221_X1 port map( B1 => n650, B2 => n2138, C1 => n1847, C2 => n2133
                           , A => n818, ZN => n1553);
   U279 : AOI222_X1 port map( A1 => n2126, A2 => n26, B1 => n2120, B2 => n652, 
                           C1 => n2114, C2 => n90, ZN => n818);
   U280 : OAI221_X1 port map( B1 => n653, B2 => n2138, C1 => n1846, C2 => n2133
                           , A => n820, ZN => n1551);
   U281 : AOI222_X1 port map( A1 => n2126, A2 => n25, B1 => n2120, B2 => n655, 
                           C1 => n2114, C2 => n89, ZN => n820);
   U282 : OAI221_X1 port map( B1 => n656, B2 => n2137, C1 => n1845, C2 => n2133
                           , A => n822, ZN => n1549);
   U283 : AOI222_X1 port map( A1 => n2125, A2 => n24, B1 => n2119, B2 => n658, 
                           C1 => n2113, C2 => n88, ZN => n822);
   U284 : OAI221_X1 port map( B1 => n659, B2 => n2137, C1 => n1844, C2 => n2133
                           , A => n824, ZN => n1547);
   U285 : AOI222_X1 port map( A1 => n2125, A2 => n23, B1 => n2119, B2 => n661, 
                           C1 => n2113, C2 => n87, ZN => n824);
   U286 : OAI221_X1 port map( B1 => n662, B2 => n2137, C1 => n1843, C2 => n2133
                           , A => n826, ZN => n1545);
   U287 : AOI222_X1 port map( A1 => n2125, A2 => n22, B1 => n2119, B2 => n664, 
                           C1 => n2113, C2 => n86, ZN => n826);
   U288 : OAI221_X1 port map( B1 => n665, B2 => n2137, C1 => n1842, C2 => n2133
                           , A => n828, ZN => n1543);
   U289 : AOI222_X1 port map( A1 => n2125, A2 => n21, B1 => n2119, B2 => n667, 
                           C1 => n2113, C2 => n85, ZN => n828);
   U290 : OAI221_X1 port map( B1 => n668, B2 => n2137, C1 => n1841, C2 => n2133
                           , A => n830, ZN => n1541);
   U291 : AOI222_X1 port map( A1 => n2125, A2 => n20, B1 => n2119, B2 => n670, 
                           C1 => n2113, C2 => n84, ZN => n830);
   U292 : OAI221_X1 port map( B1 => n671, B2 => n2137, C1 => n1840, C2 => n2133
                           , A => n832, ZN => n1539);
   U293 : AOI222_X1 port map( A1 => n2125, A2 => n19, B1 => n2119, B2 => n673, 
                           C1 => n2113, C2 => n83, ZN => n832);
   U294 : OAI221_X1 port map( B1 => n674, B2 => n2137, C1 => n1839, C2 => n2133
                           , A => n834, ZN => n1537);
   U295 : AOI222_X1 port map( A1 => n2125, A2 => n18, B1 => n2119, B2 => n676, 
                           C1 => n2113, C2 => n82, ZN => n834);
   U296 : OAI221_X1 port map( B1 => n677, B2 => n2137, C1 => n1838, C2 => n2133
                           , A => n836, ZN => n1535);
   U297 : AOI222_X1 port map( A1 => n2125, A2 => n17, B1 => n2119, B2 => n679, 
                           C1 => n2113, C2 => n81, ZN => n836);
   U298 : OAI221_X1 port map( B1 => n680, B2 => n2137, C1 => n1837, C2 => n2134
                           , A => n838, ZN => n1533);
   U299 : AOI222_X1 port map( A1 => n2125, A2 => n16, B1 => n2119, B2 => n682, 
                           C1 => n2113, C2 => n80, ZN => n838);
   U300 : OAI221_X1 port map( B1 => n683, B2 => n2137, C1 => n1836, C2 => n2134
                           , A => n840, ZN => n1531);
   U301 : AOI222_X1 port map( A1 => n2125, A2 => n15, B1 => n2119, B2 => n685, 
                           C1 => n2113, C2 => n79, ZN => n840);
   U302 : OAI221_X1 port map( B1 => n686, B2 => n2137, C1 => n1835, C2 => n2134
                           , A => n842, ZN => n1529);
   U303 : AOI222_X1 port map( A1 => n2125, A2 => n14, B1 => n2119, B2 => n688, 
                           C1 => n2113, C2 => n78, ZN => n842);
   U304 : OAI221_X1 port map( B1 => n689, B2 => n2137, C1 => n1834, C2 => n2134
                           , A => n844, ZN => n1527);
   U305 : AOI222_X1 port map( A1 => n2125, A2 => n13, B1 => n2119, B2 => n691, 
                           C1 => n2113, C2 => n77, ZN => n844);
   U306 : OAI221_X1 port map( B1 => n692, B2 => n2136, C1 => n1833, C2 => n2134
                           , A => n846, ZN => n1525);
   U307 : AOI222_X1 port map( A1 => n2124, A2 => n694, B1 => n2118, B2 => n695,
                           C1 => n2112, C2 => n76, ZN => n846);
   U308 : OAI221_X1 port map( B1 => n696, B2 => n2136, C1 => n1832, C2 => n2134
                           , A => n848, ZN => n1523);
   U309 : AOI222_X1 port map( A1 => n2124, A2 => n698, B1 => n2118, B2 => n699,
                           C1 => n2112, C2 => n75, ZN => n848);
   U310 : OAI221_X1 port map( B1 => n700, B2 => n2136, C1 => n1831, C2 => n2134
                           , A => n850, ZN => n1521);
   U311 : AOI222_X1 port map( A1 => n2124, A2 => n702, B1 => n2118, B2 => n703,
                           C1 => n2112, C2 => n74, ZN => n850);
   U312 : OAI221_X1 port map( B1 => n704, B2 => n2136, C1 => n1830, C2 => n2134
                           , A => n852, ZN => n1519);
   U313 : AOI222_X1 port map( A1 => n2124, A2 => n9, B1 => n2118, B2 => n706, 
                           C1 => n2112, C2 => n73, ZN => n852);
   U314 : OAI221_X1 port map( B1 => n707, B2 => n2136, C1 => n1829, C2 => n2134
                           , A => n854, ZN => n1517);
   U315 : AOI222_X1 port map( A1 => n2124, A2 => n8, B1 => n2118, B2 => n709, 
                           C1 => n2112, C2 => n72, ZN => n854);
   U316 : OAI221_X1 port map( B1 => n710, B2 => n2136, C1 => n1828, C2 => n2134
                           , A => n856, ZN => n1515);
   U317 : AOI222_X1 port map( A1 => n2124, A2 => n7, B1 => n2118, B2 => n712, 
                           C1 => n2112, C2 => n71, ZN => n856);
   U318 : OAI221_X1 port map( B1 => n713, B2 => n2136, C1 => n1827, C2 => n2134
                           , A => n858, ZN => n1513);
   U319 : AOI222_X1 port map( A1 => n2124, A2 => n6, B1 => n2118, B2 => n715, 
                           C1 => n2112, C2 => n70, ZN => n858);
   U320 : OAI221_X1 port map( B1 => n716, B2 => n2136, C1 => n1826, C2 => n2135
                           , A => n860, ZN => n1511);
   U321 : AOI222_X1 port map( A1 => n2124, A2 => n5, B1 => n2118, B2 => n718, 
                           C1 => n2112, C2 => n69, ZN => n860);
   U322 : OAI221_X1 port map( B1 => n719, B2 => n2136, C1 => n1825, C2 => n2134
                           , A => n862, ZN => n1509);
   U323 : AOI222_X1 port map( A1 => n2124, A2 => n4, B1 => n2118, B2 => n721, 
                           C1 => n2112, C2 => n68, ZN => n862);
   U324 : OAI221_X1 port map( B1 => n722, B2 => n2136, C1 => n1824, C2 => n2135
                           , A => n864, ZN => n1507);
   U325 : AOI222_X1 port map( A1 => n2124, A2 => n3, B1 => n2118, B2 => n724, 
                           C1 => n2112, C2 => n67, ZN => n864);
   U326 : OAI221_X1 port map( B1 => n725, B2 => n2136, C1 => n1823, C2 => n2135
                           , A => n866, ZN => n1505);
   U327 : AOI222_X1 port map( A1 => n2124, A2 => n2, B1 => n2118, B2 => n727, 
                           C1 => n2112, C2 => n66, ZN => n866);
   U328 : OAI221_X1 port map( B1 => n728, B2 => n2136, C1 => n1822, C2 => n2135
                           , A => n868, ZN => n1503);
   U329 : AOI222_X1 port map( A1 => n2124, A2 => n730, B1 => n2118, B2 => n731,
                           C1 => n2112, C2 => n65, ZN => n868);
   U330 : INV_X1 port map( A => RESET, ZN => n734);
   U331 : OAI221_X1 port map( B1 => n2170, B2 => n522, C1 => n1949, C2 => n2159
                           , A => n524, ZN => n1693);
   U332 : AOI222_X1 port map( A1 => n64, A2 => n2155, B1 => n192, B2 => n2148, 
                           C1 => n2147, C2 => n528, ZN => n524);
   U333 : OAI221_X1 port map( B1 => n2170, B2 => n529, C1 => n1948, C2 => n2159
                           , A => n530, ZN => n1692);
   U334 : AOI222_X1 port map( A1 => n63, A2 => n2153, B1 => n191, B2 => n2148, 
                           C1 => n2147, C2 => n531, ZN => n530);
   U335 : OAI221_X1 port map( B1 => n2170, B2 => n532, C1 => n1947, C2 => n2159
                           , A => n533, ZN => n1691);
   U336 : AOI222_X1 port map( A1 => n62, A2 => n2153, B1 => n190, B2 => n2148, 
                           C1 => n2146, C2 => n534, ZN => n533);
   U337 : OAI221_X1 port map( B1 => n2170, B2 => n535, C1 => n1946, C2 => n2159
                           , A => n536, ZN => n1690);
   U338 : AOI222_X1 port map( A1 => n61, A2 => n2153, B1 => n189, B2 => n2148, 
                           C1 => n2146, C2 => n537, ZN => n536);
   U339 : OAI221_X1 port map( B1 => n2167, B2 => n619, C1 => n1921, C2 => n2161
                           , A => n620, ZN => n1665);
   U340 : AOI222_X1 port map( A1 => n36, A2 => n2155, B1 => n2150, B2 => n621, 
                           C1 => n2144, C2 => n622, ZN => n620);
   U341 : OAI221_X1 port map( B1 => n2167, B2 => n623, C1 => n1920, C2 => n2161
                           , A => n624, ZN => n1664);
   U342 : AOI222_X1 port map( A1 => n35, A2 => n2155, B1 => n2150, B2 => n625, 
                           C1 => n99, C2 => n2144, ZN => n624);
   U343 : OAI221_X1 port map( B1 => n2167, B2 => n626, C1 => n1919, C2 => n2161
                           , A => n627, ZN => n1663);
   U344 : AOI222_X1 port map( A1 => n34, A2 => n2155, B1 => n2150, B2 => n628, 
                           C1 => n98, C2 => n2144, ZN => n627);
   U345 : OAI221_X1 port map( B1 => n2167, B2 => n629, C1 => n1918, C2 => n2161
                           , A => n630, ZN => n1662);
   U346 : AOI222_X1 port map( A1 => n33, A2 => n2155, B1 => n2150, B2 => n631, 
                           C1 => n97, C2 => n2144, ZN => n630);
   U347 : OAI221_X1 port map( B1 => n2167, B2 => n632, C1 => n1917, C2 => n2161
                           , A => n633, ZN => n1661);
   U348 : AOI222_X1 port map( A1 => n32, A2 => n2155, B1 => n2150, B2 => n634, 
                           C1 => n96, C2 => n2144, ZN => n633);
   U349 : OAI221_X1 port map( B1 => n2167, B2 => n635, C1 => n1916, C2 => n2161
                           , A => n636, ZN => n1660);
   U350 : AOI222_X1 port map( A1 => n31, A2 => n2155, B1 => n2150, B2 => n637, 
                           C1 => n95, C2 => n2144, ZN => n636);
   U351 : OAI221_X1 port map( B1 => n2167, B2 => n638, C1 => n1915, C2 => n2161
                           , A => n639, ZN => n1659);
   U352 : AOI222_X1 port map( A1 => n30, A2 => n2155, B1 => n2150, B2 => n640, 
                           C1 => n94, C2 => n2144, ZN => n639);
   U353 : OAI221_X1 port map( B1 => n2167, B2 => n641, C1 => n1914, C2 => n2161
                           , A => n642, ZN => n1658);
   U354 : AOI222_X1 port map( A1 => n29, A2 => n2155, B1 => n2150, B2 => n643, 
                           C1 => n93, C2 => n2144, ZN => n642);
   U355 : OAI221_X1 port map( B1 => n2167, B2 => n644, C1 => n1913, C2 => n2162
                           , A => n645, ZN => n1657);
   U356 : AOI222_X1 port map( A1 => n28, A2 => n2156, B1 => n2150, B2 => n646, 
                           C1 => n92, C2 => n2144, ZN => n645);
   U357 : OAI221_X1 port map( B1 => n2167, B2 => n647, C1 => n1912, C2 => n2162
                           , A => n648, ZN => n1656);
   U358 : AOI222_X1 port map( A1 => n27, A2 => n2156, B1 => n2151, B2 => n649, 
                           C1 => n91, C2 => n2144, ZN => n648);
   U359 : OAI221_X1 port map( B1 => n2167, B2 => n650, C1 => n1911, C2 => n2162
                           , A => n651, ZN => n1655);
   U360 : AOI222_X1 port map( A1 => n26, A2 => n2156, B1 => n2151, B2 => n652, 
                           C1 => n90, C2 => n2144, ZN => n651);
   U361 : OAI221_X1 port map( B1 => n2167, B2 => n653, C1 => n1910, C2 => n2162
                           , A => n654, ZN => n1654);
   U362 : AOI222_X1 port map( A1 => n25, A2 => n2156, B1 => n2151, B2 => n655, 
                           C1 => n89, C2 => n2144, ZN => n654);
   U363 : OAI221_X1 port map( B1 => n2165, B2 => n716, C1 => n1890, C2 => n2164
                           , A => n717, ZN => n1634);
   U364 : AOI222_X1 port map( A1 => n5, A2 => n2157, B1 => n2152, B2 => n718, 
                           C1 => n69, C2 => n2142, ZN => n717);
   U365 : OAI221_X1 port map( B1 => n2165, B2 => n722, C1 => n1888, C2 => n2164
                           , A => n723, ZN => n1632);
   U366 : AOI222_X1 port map( A1 => n3, A2 => n2157, B1 => n2152, B2 => n724, 
                           C1 => n67, C2 => n2142, ZN => n723);
   U367 : OAI221_X1 port map( B1 => n2165, B2 => n725, C1 => n1887, C2 => n2164
                           , A => n726, ZN => n1631);
   U368 : AOI222_X1 port map( A1 => n2, A2 => n2157, B1 => n2152, B2 => n727, 
                           C1 => n66, C2 => n2142, ZN => n726);
   U369 : OAI221_X1 port map( B1 => n522, B2 => n2141, C1 => n1885, C2 => n2130
                           , A => n737, ZN => n1629);
   U370 : AOI222_X1 port map( A1 => n2129, A2 => n64, B1 => n2123, B2 => n192, 
                           C1 => n2117, C2 => n528, ZN => n737);
   U371 : OAI221_X1 port map( B1 => n529, B2 => n2141, C1 => n1884, C2 => n2130
                           , A => n744, ZN => n1627);
   U372 : AOI222_X1 port map( A1 => n2129, A2 => n63, B1 => n2123, B2 => n191, 
                           C1 => n2117, C2 => n531, ZN => n744);
   U373 : OAI221_X1 port map( B1 => n532, B2 => n2141, C1 => n1883, C2 => n2130
                           , A => n746, ZN => n1625);
   U374 : AOI222_X1 port map( A1 => n2129, A2 => n62, B1 => n2123, B2 => n190, 
                           C1 => n2117, C2 => n534, ZN => n746);
   U375 : OAI221_X1 port map( B1 => n535, B2 => n2141, C1 => n1882, C2 => n2130
                           , A => n748, ZN => n1623);
   U376 : AOI222_X1 port map( A1 => n2129, A2 => n61, B1 => n2123, B2 => n189, 
                           C1 => n2117, C2 => n537, ZN => n748);
   U377 : OAI221_X1 port map( B1 => n583, B2 => n2139, C1 => n1866, C2 => n2131
                           , A => n780, ZN => n1591);
   U378 : AOI222_X1 port map( A1 => n2127, A2 => n45, B1 => n2121, B2 => n585, 
                           C1 => n2115, C2 => n586, ZN => n780);
   U379 : OAI221_X1 port map( B1 => n587, B2 => n2139, C1 => n1865, C2 => n2131
                           , A => n782, ZN => n1589);
   U380 : AOI222_X1 port map( A1 => n2127, A2 => n44, B1 => n2121, B2 => n589, 
                           C1 => n2115, C2 => n590, ZN => n782);
   U381 : OAI221_X1 port map( B1 => n591, B2 => n2139, C1 => n1864, C2 => n2131
                           , A => n784, ZN => n1587);
   U382 : AOI222_X1 port map( A1 => n2127, A2 => n43, B1 => n2121, B2 => n593, 
                           C1 => n2115, C2 => n594, ZN => n784);
   U383 : OAI221_X1 port map( B1 => n595, B2 => n2139, C1 => n1863, C2 => n2131
                           , A => n786, ZN => n1585);
   U384 : AOI222_X1 port map( A1 => n2127, A2 => n42, B1 => n2121, B2 => n597, 
                           C1 => n2115, C2 => n598, ZN => n786);
   U385 : OAI221_X1 port map( B1 => n599, B2 => n2139, C1 => n1862, C2 => n2131
                           , A => n788, ZN => n1583);
   U386 : AOI222_X1 port map( A1 => n2127, A2 => n41, B1 => n2121, B2 => n601, 
                           C1 => n2115, C2 => n602, ZN => n788);
   U387 : OAI221_X1 port map( B1 => n603, B2 => n2139, C1 => n1861, C2 => n2131
                           , A => n790, ZN => n1581);
   U388 : AOI222_X1 port map( A1 => n2127, A2 => n40, B1 => n2121, B2 => n605, 
                           C1 => n2115, C2 => n606, ZN => n790);
   U389 : OAI221_X1 port map( B1 => n607, B2 => n2139, C1 => n1860, C2 => n2132
                           , A => n792, ZN => n1579);
   U390 : AOI222_X1 port map( A1 => n2127, A2 => n39, B1 => n2121, B2 => n609, 
                           C1 => n2115, C2 => n610, ZN => n792);
   U391 : OAI221_X1 port map( B1 => n611, B2 => n2139, C1 => n1859, C2 => n2132
                           , A => n794, ZN => n1577);
   U392 : AOI222_X1 port map( A1 => n2127, A2 => n38, B1 => n2121, B2 => n613, 
                           C1 => n2115, C2 => n614, ZN => n794);
   U393 : OAI221_X1 port map( B1 => n615, B2 => n2139, C1 => n1858, C2 => n2132
                           , A => n796, ZN => n1575);
   U394 : AOI222_X1 port map( A1 => n2127, A2 => n37, B1 => n2121, B2 => n617, 
                           C1 => n2115, C2 => n618, ZN => n796);
   U395 : OAI221_X1 port map( B1 => n619, B2 => n2138, C1 => n1857, C2 => n2132
                           , A => n798, ZN => n1573);
   U396 : AOI222_X1 port map( A1 => n2126, A2 => n36, B1 => n2120, B2 => n621, 
                           C1 => n2114, C2 => n622, ZN => n798);
   U397 : OAI221_X1 port map( B1 => n2169, B2 => n538, C1 => n1945, C2 => n2159
                           , A => n539, ZN => n1689);
   U398 : AOI222_X1 port map( A1 => n60, A2 => n2153, B1 => n188, B2 => n2148, 
                           C1 => n2146, C2 => n540, ZN => n539);
   U399 : OAI221_X1 port map( B1 => n2169, B2 => n541, C1 => n1944, C2 => n2159
                           , A => n542, ZN => n1688);
   U400 : AOI222_X1 port map( A1 => n59, A2 => n2153, B1 => n187, B2 => n2148, 
                           C1 => n2146, C2 => n543, ZN => n542);
   U401 : OAI221_X1 port map( B1 => n2169, B2 => n544, C1 => n1943, C2 => n2159
                           , A => n545, ZN => n1687);
   U402 : AOI222_X1 port map( A1 => n58, A2 => n2153, B1 => n186, B2 => n2148, 
                           C1 => n2146, C2 => n546, ZN => n545);
   U403 : OAI221_X1 port map( B1 => n2169, B2 => n547, C1 => n1942, C2 => n2159
                           , A => n548, ZN => n1686);
   U404 : AOI222_X1 port map( A1 => n57, A2 => n2153, B1 => n185, B2 => n2148, 
                           C1 => n2146, C2 => n549, ZN => n548);
   U405 : OAI221_X1 port map( B1 => n2169, B2 => n550, C1 => n1941, C2 => n2159
                           , A => n551, ZN => n1685);
   U406 : AOI222_X1 port map( A1 => n56, A2 => n2153, B1 => n184, B2 => n2148, 
                           C1 => n2146, C2 => n552, ZN => n551);
   U407 : OAI221_X1 port map( B1 => n2169, B2 => n553, C1 => n1940, C2 => n2159
                           , A => n554, ZN => n1684);
   U408 : AOI222_X1 port map( A1 => n55, A2 => n2153, B1 => n183, B2 => n2148, 
                           C1 => n2146, C2 => n555, ZN => n554);
   U409 : OAI221_X1 port map( B1 => n2169, B2 => n556, C1 => n1939, C2 => n2159
                           , A => n557, ZN => n1683);
   U410 : AOI222_X1 port map( A1 => n54, A2 => n2153, B1 => n182, B2 => n2148, 
                           C1 => n2146, C2 => n558, ZN => n557);
   U411 : OAI221_X1 port map( B1 => n2169, B2 => n559, C1 => n1938, C2 => n2159
                           , A => n560, ZN => n1682);
   U412 : AOI222_X1 port map( A1 => n53, A2 => n2153, B1 => n181, B2 => n2148, 
                           C1 => n2146, C2 => n561, ZN => n560);
   U413 : OAI221_X1 port map( B1 => n2168, B2 => n583, C1 => n1930, C2 => n2160
                           , A => n584, ZN => n1674);
   U414 : AOI222_X1 port map( A1 => n45, A2 => n2154, B1 => n2149, B2 => n585, 
                           C1 => n2145, C2 => n586, ZN => n584);
   U415 : OAI221_X1 port map( B1 => n2168, B2 => n587, C1 => n1929, C2 => n2160
                           , A => n588, ZN => n1673);
   U416 : AOI222_X1 port map( A1 => n44, A2 => n2154, B1 => n2149, B2 => n589, 
                           C1 => n2145, C2 => n590, ZN => n588);
   U417 : OAI221_X1 port map( B1 => n2168, B2 => n591, C1 => n1928, C2 => n2160
                           , A => n592, ZN => n1672);
   U418 : AOI222_X1 port map( A1 => n43, A2 => n2154, B1 => n2149, B2 => n593, 
                           C1 => n2145, C2 => n594, ZN => n592);
   U419 : OAI221_X1 port map( B1 => n2168, B2 => n595, C1 => n1927, C2 => n2160
                           , A => n596, ZN => n1671);
   U420 : AOI222_X1 port map( A1 => n42, A2 => n2154, B1 => n2149, B2 => n597, 
                           C1 => n2145, C2 => n598, ZN => n596);
   U421 : OAI221_X1 port map( B1 => n2168, B2 => n599, C1 => n1926, C2 => n2160
                           , A => n600, ZN => n1670);
   U422 : AOI222_X1 port map( A1 => n41, A2 => n2154, B1 => n2149, B2 => n601, 
                           C1 => n2145, C2 => n602, ZN => n600);
   U423 : OAI221_X1 port map( B1 => n2168, B2 => n603, C1 => n1925, C2 => n2160
                           , A => n604, ZN => n1669);
   U424 : AOI222_X1 port map( A1 => n40, A2 => n2154, B1 => n2150, B2 => n605, 
                           C1 => n2145, C2 => n606, ZN => n604);
   U425 : OAI221_X1 port map( B1 => n2168, B2 => n607, C1 => n1924, C2 => n2161
                           , A => n608, ZN => n1668);
   U426 : AOI222_X1 port map( A1 => n39, A2 => n2155, B1 => n2150, B2 => n609, 
                           C1 => n2145, C2 => n610, ZN => n608);
   U427 : OAI221_X1 port map( B1 => n2168, B2 => n611, C1 => n1923, C2 => n2161
                           , A => n612, ZN => n1667);
   U428 : AOI222_X1 port map( A1 => n38, A2 => n2155, B1 => n2150, B2 => n613, 
                           C1 => n2145, C2 => n614, ZN => n612);
   U429 : OAI221_X1 port map( B1 => n2168, B2 => n615, C1 => n1922, C2 => n2161
                           , A => n616, ZN => n1666);
   U430 : AOI222_X1 port map( A1 => n37, A2 => n2155, B1 => n2150, B2 => n617, 
                           C1 => n2145, C2 => n618, ZN => n616);
   U431 : OAI22_X1 port map( A1 => n1950, A2 => n2099, B1 => n743, B2 => n2093,
                           ZN => n1501);
   U432 : OAI22_X1 port map( A1 => n1951, A2 => n2099, B1 => n745, B2 => n2093,
                           ZN => n1500);
   U433 : OAI22_X1 port map( A1 => n1952, A2 => n2099, B1 => n747, B2 => n2093,
                           ZN => n1499);
   U434 : OAI22_X1 port map( A1 => n1953, A2 => n2099, B1 => n749, B2 => n2093,
                           ZN => n1498);
   U435 : OAI22_X1 port map( A1 => n1821, A2 => n2087, B1 => n743, B2 => n2081,
                           ZN => n1437);
   U436 : OAI22_X1 port map( A1 => n1820, A2 => n2087, B1 => n745, B2 => n2081,
                           ZN => n1436);
   U437 : OAI22_X1 port map( A1 => n1819, A2 => n2087, B1 => n747, B2 => n2081,
                           ZN => n1435);
   U438 : OAI22_X1 port map( A1 => n1818, A2 => n2087, B1 => n749, B2 => n2081,
                           ZN => n1434);
   U439 : OAI22_X1 port map( A1 => n2010, A2 => n2075, B1 => n743, B2 => n2069,
                           ZN => n1373);
   U440 : OAI22_X1 port map( A1 => n2011, A2 => n2075, B1 => n745, B2 => n2069,
                           ZN => n1372);
   U441 : OAI22_X1 port map( A1 => n2012, A2 => n2075, B1 => n747, B2 => n2069,
                           ZN => n1371);
   U442 : OAI22_X1 port map( A1 => n2013, A2 => n2075, B1 => n749, B2 => n2069,
                           ZN => n1370);
   U443 : OAI22_X1 port map( A1 => n1954, A2 => n2099, B1 => n751, B2 => n2092,
                           ZN => n1497);
   U444 : OAI22_X1 port map( A1 => n1955, A2 => n2098, B1 => n753, B2 => n2092,
                           ZN => n1496);
   U445 : OAI22_X1 port map( A1 => n1956, A2 => n2098, B1 => n755, B2 => n2092,
                           ZN => n1495);
   U446 : OAI22_X1 port map( A1 => n1957, A2 => n2098, B1 => n757, B2 => n2092,
                           ZN => n1494);
   U447 : OAI22_X1 port map( A1 => n1958, A2 => n2098, B1 => n759, B2 => n2092,
                           ZN => n1493);
   U448 : OAI22_X1 port map( A1 => n1959, A2 => n2098, B1 => n761, B2 => n2092,
                           ZN => n1492);
   U449 : OAI22_X1 port map( A1 => n1960, A2 => n2098, B1 => n763, B2 => n2092,
                           ZN => n1491);
   U450 : OAI22_X1 port map( A1 => n1961, A2 => n2098, B1 => n765, B2 => n2092,
                           ZN => n1490);
   U451 : OAI22_X1 port map( A1 => n1962, A2 => n2098, B1 => n767, B2 => n2092,
                           ZN => n1489);
   U452 : OAI22_X1 port map( A1 => n1963, A2 => n2098, B1 => n769, B2 => n2092,
                           ZN => n1488);
   U453 : OAI22_X1 port map( A1 => n1964, A2 => n2098, B1 => n771, B2 => n2092,
                           ZN => n1487);
   U454 : OAI22_X1 port map( A1 => n1965, A2 => n2098, B1 => n773, B2 => n2092,
                           ZN => n1486);
   U455 : OAI22_X1 port map( A1 => n1966, A2 => n2098, B1 => n775, B2 => n2091,
                           ZN => n1485);
   U456 : OAI22_X1 port map( A1 => n1967, A2 => n2097, B1 => n777, B2 => n2091,
                           ZN => n1484);
   U457 : OAI22_X1 port map( A1 => n1968, A2 => n2097, B1 => n779, B2 => n2091,
                           ZN => n1483);
   U458 : OAI22_X1 port map( A1 => n1969, A2 => n2097, B1 => n781, B2 => n2091,
                           ZN => n1482);
   U459 : OAI22_X1 port map( A1 => n1970, A2 => n2097, B1 => n783, B2 => n2091,
                           ZN => n1481);
   U460 : OAI22_X1 port map( A1 => n1971, A2 => n2097, B1 => n785, B2 => n2091,
                           ZN => n1480);
   U461 : OAI22_X1 port map( A1 => n1972, A2 => n2097, B1 => n787, B2 => n2091,
                           ZN => n1479);
   U462 : OAI22_X1 port map( A1 => n1973, A2 => n2097, B1 => n789, B2 => n2091,
                           ZN => n1478);
   U463 : OAI22_X1 port map( A1 => n1974, A2 => n2097, B1 => n791, B2 => n2091,
                           ZN => n1477);
   U464 : OAI22_X1 port map( A1 => n1975, A2 => n2097, B1 => n793, B2 => n2091,
                           ZN => n1476);
   U465 : OAI22_X1 port map( A1 => n1976, A2 => n2097, B1 => n795, B2 => n2091,
                           ZN => n1475);
   U466 : OAI22_X1 port map( A1 => n1977, A2 => n2097, B1 => n797, B2 => n2091,
                           ZN => n1474);
   U467 : OAI22_X1 port map( A1 => n1978, A2 => n2097, B1 => n799, B2 => n2090,
                           ZN => n1473);
   U468 : OAI22_X1 port map( A1 => n1979, A2 => n2096, B1 => n801, B2 => n2090,
                           ZN => n1472);
   U469 : OAI22_X1 port map( A1 => n1980, A2 => n2096, B1 => n803, B2 => n2090,
                           ZN => n1471);
   U470 : OAI22_X1 port map( A1 => n1981, A2 => n2096, B1 => n805, B2 => n2090,
                           ZN => n1470);
   U471 : OAI22_X1 port map( A1 => n1982, A2 => n2096, B1 => n807, B2 => n2090,
                           ZN => n1469);
   U472 : OAI22_X1 port map( A1 => n1983, A2 => n2096, B1 => n809, B2 => n2090,
                           ZN => n1468);
   U473 : OAI22_X1 port map( A1 => n1984, A2 => n2096, B1 => n811, B2 => n2090,
                           ZN => n1467);
   U474 : OAI22_X1 port map( A1 => n1985, A2 => n2096, B1 => n813, B2 => n2090,
                           ZN => n1466);
   U475 : OAI22_X1 port map( A1 => n1986, A2 => n2096, B1 => n815, B2 => n2090,
                           ZN => n1465);
   U476 : OAI22_X1 port map( A1 => n1987, A2 => n2096, B1 => n817, B2 => n2090,
                           ZN => n1464);
   U477 : OAI22_X1 port map( A1 => n1988, A2 => n2096, B1 => n819, B2 => n2090,
                           ZN => n1463);
   U478 : OAI22_X1 port map( A1 => n1989, A2 => n2096, B1 => n821, B2 => n2090,
                           ZN => n1462);
   U479 : OAI22_X1 port map( A1 => n1990, A2 => n2096, B1 => n823, B2 => n2089,
                           ZN => n1461);
   U480 : OAI22_X1 port map( A1 => n1991, A2 => n2095, B1 => n825, B2 => n2089,
                           ZN => n1460);
   U481 : OAI22_X1 port map( A1 => n1992, A2 => n2095, B1 => n827, B2 => n2089,
                           ZN => n1459);
   U482 : OAI22_X1 port map( A1 => n1993, A2 => n2095, B1 => n829, B2 => n2089,
                           ZN => n1458);
   U483 : OAI22_X1 port map( A1 => n1994, A2 => n2095, B1 => n831, B2 => n2089,
                           ZN => n1457);
   U484 : OAI22_X1 port map( A1 => n1995, A2 => n2095, B1 => n833, B2 => n2089,
                           ZN => n1456);
   U485 : OAI22_X1 port map( A1 => n1996, A2 => n2095, B1 => n835, B2 => n2089,
                           ZN => n1455);
   U486 : OAI22_X1 port map( A1 => n1997, A2 => n2095, B1 => n837, B2 => n2089,
                           ZN => n1454);
   U487 : OAI22_X1 port map( A1 => n1998, A2 => n2095, B1 => n839, B2 => n2089,
                           ZN => n1453);
   U488 : OAI22_X1 port map( A1 => n1999, A2 => n2095, B1 => n841, B2 => n2089,
                           ZN => n1452);
   U489 : OAI22_X1 port map( A1 => n2000, A2 => n2095, B1 => n843, B2 => n2089,
                           ZN => n1451);
   U490 : OAI22_X1 port map( A1 => n2001, A2 => n2095, B1 => n845, B2 => n2089,
                           ZN => n1450);
   U491 : OAI22_X1 port map( A1 => n1204, A2 => n2095, B1 => n847, B2 => n2088,
                           ZN => n1449);
   U492 : OAI22_X1 port map( A1 => n1202, A2 => n2094, B1 => n849, B2 => n2088,
                           ZN => n1448);
   U493 : OAI22_X1 port map( A1 => n1200, A2 => n2094, B1 => n851, B2 => n2088,
                           ZN => n1447);
   U494 : OAI22_X1 port map( A1 => n2002, A2 => n2094, B1 => n853, B2 => n2088,
                           ZN => n1446);
   U495 : OAI22_X1 port map( A1 => n2003, A2 => n2094, B1 => n855, B2 => n2088,
                           ZN => n1445);
   U496 : OAI22_X1 port map( A1 => n2004, A2 => n2094, B1 => n857, B2 => n2088,
                           ZN => n1444);
   U497 : OAI22_X1 port map( A1 => n2005, A2 => n2094, B1 => n859, B2 => n2088,
                           ZN => n1443);
   U498 : OAI22_X1 port map( A1 => n2006, A2 => n2094, B1 => n861, B2 => n2088,
                           ZN => n1442);
   U499 : OAI22_X1 port map( A1 => n2007, A2 => n2094, B1 => n863, B2 => n2088,
                           ZN => n1441);
   U500 : OAI22_X1 port map( A1 => n2008, A2 => n2094, B1 => n865, B2 => n2088,
                           ZN => n1440);
   U501 : OAI22_X1 port map( A1 => n2009, A2 => n2094, B1 => n867, B2 => n2088,
                           ZN => n1439);
   U502 : OAI22_X1 port map( A1 => n415, A2 => n2094, B1 => n871, B2 => n2088, 
                           ZN => n1438);
   U503 : OAI22_X1 port map( A1 => n1817, A2 => n2087, B1 => n751, B2 => n2080,
                           ZN => n1433);
   U504 : OAI22_X1 port map( A1 => n1816, A2 => n2086, B1 => n753, B2 => n2080,
                           ZN => n1432);
   U505 : OAI22_X1 port map( A1 => n1815, A2 => n2086, B1 => n755, B2 => n2080,
                           ZN => n1431);
   U506 : OAI22_X1 port map( A1 => n1814, A2 => n2086, B1 => n757, B2 => n2080,
                           ZN => n1430);
   U507 : OAI22_X1 port map( A1 => n1813, A2 => n2086, B1 => n759, B2 => n2080,
                           ZN => n1429);
   U508 : OAI22_X1 port map( A1 => n1812, A2 => n2086, B1 => n761, B2 => n2080,
                           ZN => n1428);
   U509 : OAI22_X1 port map( A1 => n1811, A2 => n2086, B1 => n763, B2 => n2080,
                           ZN => n1427);
   U510 : OAI22_X1 port map( A1 => n1810, A2 => n2086, B1 => n765, B2 => n2080,
                           ZN => n1426);
   U511 : OAI22_X1 port map( A1 => n1809, A2 => n2086, B1 => n767, B2 => n2080,
                           ZN => n1425);
   U512 : OAI22_X1 port map( A1 => n1808, A2 => n2086, B1 => n769, B2 => n2080,
                           ZN => n1424);
   U513 : OAI22_X1 port map( A1 => n1807, A2 => n2086, B1 => n771, B2 => n2080,
                           ZN => n1423);
   U514 : OAI22_X1 port map( A1 => n1806, A2 => n2086, B1 => n773, B2 => n2080,
                           ZN => n1422);
   U515 : OAI22_X1 port map( A1 => n1805, A2 => n2086, B1 => n775, B2 => n2079,
                           ZN => n1421);
   U516 : OAI22_X1 port map( A1 => n1804, A2 => n2085, B1 => n777, B2 => n2079,
                           ZN => n1420);
   U517 : OAI22_X1 port map( A1 => n1803, A2 => n2085, B1 => n779, B2 => n2079,
                           ZN => n1419);
   U518 : OAI22_X1 port map( A1 => n1802, A2 => n2085, B1 => n781, B2 => n2079,
                           ZN => n1418);
   U519 : OAI22_X1 port map( A1 => n1801, A2 => n2085, B1 => n783, B2 => n2079,
                           ZN => n1417);
   U520 : OAI22_X1 port map( A1 => n1800, A2 => n2085, B1 => n785, B2 => n2079,
                           ZN => n1416);
   U521 : OAI22_X1 port map( A1 => n1799, A2 => n2085, B1 => n787, B2 => n2079,
                           ZN => n1415);
   U522 : OAI22_X1 port map( A1 => n1798, A2 => n2085, B1 => n789, B2 => n2079,
                           ZN => n1414);
   U523 : OAI22_X1 port map( A1 => n1797, A2 => n2085, B1 => n791, B2 => n2079,
                           ZN => n1413);
   U524 : OAI22_X1 port map( A1 => n1796, A2 => n2085, B1 => n793, B2 => n2079,
                           ZN => n1412);
   U525 : OAI22_X1 port map( A1 => n1795, A2 => n2085, B1 => n795, B2 => n2079,
                           ZN => n1411);
   U526 : OAI22_X1 port map( A1 => n1794, A2 => n2085, B1 => n797, B2 => n2079,
                           ZN => n1410);
   U527 : OAI22_X1 port map( A1 => n1793, A2 => n2085, B1 => n799, B2 => n2078,
                           ZN => n1409);
   U528 : OAI22_X1 port map( A1 => n2029, A2 => n2084, B1 => n801, B2 => n2078,
                           ZN => n1408);
   U529 : OAI22_X1 port map( A1 => n2030, A2 => n2084, B1 => n803, B2 => n2078,
                           ZN => n1407);
   U530 : OAI22_X1 port map( A1 => n2031, A2 => n2084, B1 => n805, B2 => n2078,
                           ZN => n1406);
   U531 : OAI22_X1 port map( A1 => n2032, A2 => n2084, B1 => n807, B2 => n2078,
                           ZN => n1405);
   U532 : OAI22_X1 port map( A1 => n2033, A2 => n2084, B1 => n809, B2 => n2078,
                           ZN => n1404);
   U533 : OAI22_X1 port map( A1 => n2034, A2 => n2084, B1 => n811, B2 => n2078,
                           ZN => n1403);
   U534 : OAI22_X1 port map( A1 => n2035, A2 => n2084, B1 => n813, B2 => n2078,
                           ZN => n1402);
   U535 : OAI22_X1 port map( A1 => n2036, A2 => n2084, B1 => n815, B2 => n2078,
                           ZN => n1401);
   U536 : OAI22_X1 port map( A1 => n2037, A2 => n2084, B1 => n817, B2 => n2078,
                           ZN => n1400);
   U537 : OAI22_X1 port map( A1 => n2038, A2 => n2084, B1 => n819, B2 => n2078,
                           ZN => n1399);
   U538 : OAI22_X1 port map( A1 => n2039, A2 => n2084, B1 => n821, B2 => n2078,
                           ZN => n1398);
   U539 : OAI22_X1 port map( A1 => n2040, A2 => n2084, B1 => n823, B2 => n2077,
                           ZN => n1397);
   U540 : OAI22_X1 port map( A1 => n2041, A2 => n2083, B1 => n825, B2 => n2077,
                           ZN => n1396);
   U541 : OAI22_X1 port map( A1 => n2042, A2 => n2083, B1 => n827, B2 => n2077,
                           ZN => n1395);
   U542 : OAI22_X1 port map( A1 => n2043, A2 => n2083, B1 => n829, B2 => n2077,
                           ZN => n1394);
   U543 : OAI22_X1 port map( A1 => n2044, A2 => n2083, B1 => n831, B2 => n2077,
                           ZN => n1393);
   U544 : OAI22_X1 port map( A1 => n2045, A2 => n2083, B1 => n833, B2 => n2077,
                           ZN => n1392);
   U545 : OAI22_X1 port map( A1 => n2046, A2 => n2083, B1 => n835, B2 => n2077,
                           ZN => n1391);
   U546 : OAI22_X1 port map( A1 => n2047, A2 => n2083, B1 => n837, B2 => n2077,
                           ZN => n1390);
   U547 : OAI22_X1 port map( A1 => n2048, A2 => n2083, B1 => n839, B2 => n2077,
                           ZN => n1389);
   U548 : OAI22_X1 port map( A1 => n2049, A2 => n2083, B1 => n841, B2 => n2077,
                           ZN => n1388);
   U549 : OAI22_X1 port map( A1 => n2050, A2 => n2083, B1 => n843, B2 => n2077,
                           ZN => n1387);
   U550 : OAI22_X1 port map( A1 => n2051, A2 => n2083, B1 => n845, B2 => n2077,
                           ZN => n1386);
   U551 : OAI22_X1 port map( A1 => n2052, A2 => n2083, B1 => n847, B2 => n2076,
                           ZN => n1385);
   U552 : OAI22_X1 port map( A1 => n2053, A2 => n2082, B1 => n849, B2 => n2076,
                           ZN => n1384);
   U553 : OAI22_X1 port map( A1 => n2054, A2 => n2082, B1 => n851, B2 => n2076,
                           ZN => n1383);
   U554 : OAI22_X1 port map( A1 => n2055, A2 => n2082, B1 => n853, B2 => n2076,
                           ZN => n1382);
   U555 : OAI22_X1 port map( A1 => n2056, A2 => n2082, B1 => n855, B2 => n2076,
                           ZN => n1381);
   U556 : OAI22_X1 port map( A1 => n2057, A2 => n2082, B1 => n857, B2 => n2076,
                           ZN => n1380);
   U557 : OAI22_X1 port map( A1 => n2058, A2 => n2082, B1 => n859, B2 => n2076,
                           ZN => n1379);
   U558 : OAI22_X1 port map( A1 => n2059, A2 => n2082, B1 => n861, B2 => n2076,
                           ZN => n1378);
   U559 : OAI22_X1 port map( A1 => n2060, A2 => n2082, B1 => n863, B2 => n2076,
                           ZN => n1377);
   U560 : OAI22_X1 port map( A1 => n2061, A2 => n2082, B1 => n865, B2 => n2076,
                           ZN => n1376);
   U561 : OAI22_X1 port map( A1 => n2062, A2 => n2082, B1 => n867, B2 => n2076,
                           ZN => n1375);
   U562 : OAI22_X1 port map( A1 => n2063, A2 => n2082, B1 => n871, B2 => n2076,
                           ZN => n1374);
   U563 : OAI22_X1 port map( A1 => n2014, A2 => n2075, B1 => n751, B2 => n2068,
                           ZN => n1369);
   U564 : OAI22_X1 port map( A1 => n2015, A2 => n2074, B1 => n753, B2 => n2068,
                           ZN => n1368);
   U565 : OAI22_X1 port map( A1 => n2016, A2 => n2074, B1 => n755, B2 => n2068,
                           ZN => n1367);
   U566 : OAI22_X1 port map( A1 => n2017, A2 => n2074, B1 => n757, B2 => n2068,
                           ZN => n1366);
   U567 : OAI22_X1 port map( A1 => n2018, A2 => n2074, B1 => n759, B2 => n2068,
                           ZN => n1365);
   U568 : OAI22_X1 port map( A1 => n2019, A2 => n2074, B1 => n761, B2 => n2068,
                           ZN => n1364);
   U569 : OAI22_X1 port map( A1 => n2020, A2 => n2074, B1 => n763, B2 => n2068,
                           ZN => n1363);
   U570 : OAI22_X1 port map( A1 => n2021, A2 => n2074, B1 => n765, B2 => n2068,
                           ZN => n1362);
   U571 : OAI22_X1 port map( A1 => n2022, A2 => n2074, B1 => n767, B2 => n2068,
                           ZN => n1361);
   U572 : OAI22_X1 port map( A1 => n2023, A2 => n2074, B1 => n769, B2 => n2068,
                           ZN => n1360);
   U573 : OAI22_X1 port map( A1 => n2024, A2 => n2074, B1 => n771, B2 => n2068,
                           ZN => n1359);
   U574 : OAI22_X1 port map( A1 => n2025, A2 => n2074, B1 => n773, B2 => n2068,
                           ZN => n1358);
   U575 : OAI22_X1 port map( A1 => n2026, A2 => n2074, B1 => n775, B2 => n2067,
                           ZN => n1357);
   U576 : OAI22_X1 port map( A1 => n2027, A2 => n2073, B1 => n777, B2 => n2067,
                           ZN => n1356);
   U577 : OAI22_X1 port map( A1 => n2028, A2 => n2073, B1 => n779, B2 => n2067,
                           ZN => n1355);
   U578 : OAI22_X1 port map( A1 => n1738, A2 => n2073, B1 => n781, B2 => n2067,
                           ZN => n1354);
   U579 : OAI22_X1 port map( A1 => n1737, A2 => n2073, B1 => n783, B2 => n2067,
                           ZN => n1353);
   U580 : OAI22_X1 port map( A1 => n1736, A2 => n2073, B1 => n785, B2 => n2067,
                           ZN => n1352);
   U581 : OAI22_X1 port map( A1 => n1735, A2 => n2073, B1 => n787, B2 => n2067,
                           ZN => n1351);
   U582 : OAI22_X1 port map( A1 => n1734, A2 => n2073, B1 => n789, B2 => n2067,
                           ZN => n1350);
   U583 : OAI22_X1 port map( A1 => n1733, A2 => n2073, B1 => n791, B2 => n2067,
                           ZN => n1349);
   U584 : OAI22_X1 port map( A1 => n1732, A2 => n2073, B1 => n793, B2 => n2067,
                           ZN => n1348);
   U585 : OAI22_X1 port map( A1 => n1731, A2 => n2073, B1 => n795, B2 => n2067,
                           ZN => n1347);
   U586 : OAI22_X1 port map( A1 => n1730, A2 => n2073, B1 => n797, B2 => n2067,
                           ZN => n1346);
   U587 : OAI22_X1 port map( A1 => n1729, A2 => n2073, B1 => n799, B2 => n2066,
                           ZN => n1345);
   U588 : OAI22_X1 port map( A1 => n1728, A2 => n2072, B1 => n801, B2 => n2066,
                           ZN => n1344);
   U589 : OAI22_X1 port map( A1 => n1727, A2 => n2072, B1 => n803, B2 => n2066,
                           ZN => n1343);
   U590 : OAI22_X1 port map( A1 => n1726, A2 => n2072, B1 => n805, B2 => n2066,
                           ZN => n1342);
   U591 : OAI22_X1 port map( A1 => n1725, A2 => n2072, B1 => n807, B2 => n2066,
                           ZN => n1341);
   U592 : OAI22_X1 port map( A1 => n1724, A2 => n2072, B1 => n809, B2 => n2066,
                           ZN => n1340);
   U593 : OAI22_X1 port map( A1 => n1723, A2 => n2072, B1 => n811, B2 => n2066,
                           ZN => n1339);
   U594 : OAI22_X1 port map( A1 => n1722, A2 => n2072, B1 => n813, B2 => n2066,
                           ZN => n1338);
   U595 : OAI22_X1 port map( A1 => n1721, A2 => n2072, B1 => n815, B2 => n2066,
                           ZN => n1337);
   U596 : OAI22_X1 port map( A1 => n1720, A2 => n2072, B1 => n817, B2 => n2066,
                           ZN => n1336);
   U597 : OAI22_X1 port map( A1 => n1719, A2 => n2072, B1 => n819, B2 => n2066,
                           ZN => n1335);
   U598 : OAI22_X1 port map( A1 => n1718, A2 => n2072, B1 => n821, B2 => n2066,
                           ZN => n1334);
   U599 : OAI22_X1 port map( A1 => n1717, A2 => n2072, B1 => n823, B2 => n2065,
                           ZN => n1333);
   U600 : OAI22_X1 port map( A1 => n1716, A2 => n2071, B1 => n825, B2 => n2065,
                           ZN => n1332);
   U601 : OAI22_X1 port map( A1 => n1715, A2 => n2071, B1 => n827, B2 => n2065,
                           ZN => n1331);
   U602 : OAI22_X1 port map( A1 => n1714, A2 => n2071, B1 => n829, B2 => n2065,
                           ZN => n1330);
   U603 : OAI22_X1 port map( A1 => n1713, A2 => n2071, B1 => n831, B2 => n2065,
                           ZN => n1329);
   U604 : OAI22_X1 port map( A1 => n1712, A2 => n2071, B1 => n833, B2 => n2065,
                           ZN => n1328);
   U605 : OAI22_X1 port map( A1 => n1711, A2 => n2071, B1 => n835, B2 => n2065,
                           ZN => n1327);
   U606 : OAI22_X1 port map( A1 => n1710, A2 => n2071, B1 => n837, B2 => n2065,
                           ZN => n1326);
   U607 : OAI22_X1 port map( A1 => n1709, A2 => n2071, B1 => n839, B2 => n2065,
                           ZN => n1325);
   U608 : OAI22_X1 port map( A1 => n1708, A2 => n2071, B1 => n841, B2 => n2065,
                           ZN => n1324);
   U609 : OAI22_X1 port map( A1 => n1707, A2 => n2071, B1 => n843, B2 => n2065,
                           ZN => n1323);
   U610 : OAI22_X1 port map( A1 => n1706, A2 => n2071, B1 => n845, B2 => n2065,
                           ZN => n1322);
   U611 : OAI22_X1 port map( A1 => n1705, A2 => n2071, B1 => n847, B2 => n2064,
                           ZN => n1321);
   U612 : OAI22_X1 port map( A1 => n1704, A2 => n2070, B1 => n849, B2 => n2064,
                           ZN => n1320);
   U613 : OAI22_X1 port map( A1 => n1703, A2 => n2070, B1 => n851, B2 => n2064,
                           ZN => n1319);
   U614 : OAI22_X1 port map( A1 => n1702, A2 => n2070, B1 => n853, B2 => n2064,
                           ZN => n1318);
   U615 : OAI22_X1 port map( A1 => n1701, A2 => n2070, B1 => n855, B2 => n2064,
                           ZN => n1317);
   U616 : OAI22_X1 port map( A1 => n1700, A2 => n2070, B1 => n857, B2 => n2064,
                           ZN => n1316);
   U617 : OAI22_X1 port map( A1 => n1699, A2 => n2070, B1 => n859, B2 => n2064,
                           ZN => n1315);
   U618 : OAI22_X1 port map( A1 => n1698, A2 => n2070, B1 => n861, B2 => n2064,
                           ZN => n1314);
   U619 : OAI22_X1 port map( A1 => n1697, A2 => n2070, B1 => n863, B2 => n2064,
                           ZN => n1313);
   U620 : OAI22_X1 port map( A1 => n1696, A2 => n2070, B1 => n865, B2 => n2064,
                           ZN => n1312);
   U621 : OAI22_X1 port map( A1 => n1695, A2 => n2070, B1 => n867, B2 => n2064,
                           ZN => n1311);
   U622 : OAI22_X1 port map( A1 => n1694, A2 => n2070, B1 => n871, B2 => n2064,
                           ZN => n1310);
   U623 : INV_X1 port map( A => DATAIN(0), ZN => n743);
   U624 : INV_X1 port map( A => DATAIN(1), ZN => n745);
   U625 : INV_X1 port map( A => DATAIN(2), ZN => n747);
   U626 : INV_X1 port map( A => DATAIN(3), ZN => n749);
   U627 : INV_X1 port map( A => DATAIN(4), ZN => n751);
   U628 : INV_X1 port map( A => DATAIN(5), ZN => n753);
   U629 : INV_X1 port map( A => DATAIN(6), ZN => n755);
   U630 : INV_X1 port map( A => DATAIN(7), ZN => n757);
   U631 : INV_X1 port map( A => DATAIN(8), ZN => n759);
   U632 : INV_X1 port map( A => DATAIN(9), ZN => n761);
   U633 : INV_X1 port map( A => DATAIN(10), ZN => n763);
   U634 : INV_X1 port map( A => DATAIN(11), ZN => n765);
   U635 : INV_X1 port map( A => DATAIN(12), ZN => n767);
   U636 : INV_X1 port map( A => DATAIN(13), ZN => n769);
   U637 : INV_X1 port map( A => DATAIN(14), ZN => n771);
   U638 : INV_X1 port map( A => DATAIN(15), ZN => n773);
   U639 : INV_X1 port map( A => DATAIN(16), ZN => n775);
   U640 : INV_X1 port map( A => DATAIN(17), ZN => n777);
   U641 : INV_X1 port map( A => DATAIN(18), ZN => n779);
   U642 : INV_X1 port map( A => DATAIN(19), ZN => n781);
   U643 : INV_X1 port map( A => DATAIN(20), ZN => n783);
   U644 : INV_X1 port map( A => DATAIN(21), ZN => n785);
   U645 : INV_X1 port map( A => DATAIN(22), ZN => n787);
   U646 : INV_X1 port map( A => DATAIN(23), ZN => n789);
   U647 : INV_X1 port map( A => DATAIN(24), ZN => n791);
   U648 : INV_X1 port map( A => DATAIN(25), ZN => n793);
   U649 : INV_X1 port map( A => DATAIN(26), ZN => n795);
   U650 : INV_X1 port map( A => DATAIN(27), ZN => n797);
   U651 : INV_X1 port map( A => DATAIN(28), ZN => n799);
   U652 : INV_X1 port map( A => DATAIN(29), ZN => n801);
   U653 : INV_X1 port map( A => DATAIN(30), ZN => n803);
   U654 : INV_X1 port map( A => DATAIN(31), ZN => n805);
   U655 : INV_X1 port map( A => DATAIN(32), ZN => n807);
   U656 : INV_X1 port map( A => DATAIN(33), ZN => n809);
   U657 : INV_X1 port map( A => DATAIN(34), ZN => n811);
   U658 : INV_X1 port map( A => DATAIN(35), ZN => n813);
   U659 : INV_X1 port map( A => DATAIN(36), ZN => n815);
   U660 : INV_X1 port map( A => DATAIN(37), ZN => n817);
   U661 : INV_X1 port map( A => DATAIN(38), ZN => n819);
   U662 : INV_X1 port map( A => DATAIN(39), ZN => n821);
   U663 : INV_X1 port map( A => DATAIN(40), ZN => n823);
   U664 : INV_X1 port map( A => DATAIN(41), ZN => n825);
   U665 : INV_X1 port map( A => DATAIN(42), ZN => n827);
   U666 : INV_X1 port map( A => DATAIN(43), ZN => n829);
   U667 : INV_X1 port map( A => DATAIN(44), ZN => n831);
   U668 : INV_X1 port map( A => DATAIN(45), ZN => n833);
   U669 : INV_X1 port map( A => DATAIN(46), ZN => n835);
   U670 : INV_X1 port map( A => DATAIN(47), ZN => n837);
   U671 : INV_X1 port map( A => DATAIN(48), ZN => n839);
   U672 : INV_X1 port map( A => DATAIN(49), ZN => n841);
   U673 : INV_X1 port map( A => DATAIN(50), ZN => n843);
   U674 : INV_X1 port map( A => DATAIN(51), ZN => n845);
   U675 : INV_X1 port map( A => DATAIN(52), ZN => n847);
   U676 : INV_X1 port map( A => DATAIN(53), ZN => n849);
   U677 : INV_X1 port map( A => DATAIN(54), ZN => n851);
   U678 : INV_X1 port map( A => DATAIN(55), ZN => n853);
   U679 : INV_X1 port map( A => DATAIN(56), ZN => n855);
   U680 : INV_X1 port map( A => DATAIN(57), ZN => n857);
   U681 : INV_X1 port map( A => DATAIN(58), ZN => n859);
   U682 : INV_X1 port map( A => DATAIN(59), ZN => n861);
   U683 : INV_X1 port map( A => DATAIN(60), ZN => n863);
   U684 : INV_X1 port map( A => DATAIN(61), ZN => n865);
   U685 : INV_X1 port map( A => DATAIN(62), ZN => n867);
   U686 : INV_X1 port map( A => DATAIN(63), ZN => n871);
   U687 : CLKBUF_X1 port map( A => n979, Z => n2069);
   U688 : CLKBUF_X1 port map( A => n978, Z => n2075);
   U689 : CLKBUF_X1 port map( A => n939, Z => n2081);
   U690 : CLKBUF_X1 port map( A => n938, Z => n2087);
   U691 : CLKBUF_X1 port map( A => n876, Z => n2093);
   U692 : CLKBUF_X1 port map( A => n875, Z => n2099);
   U693 : CLKBUF_X1 port map( A => n742, Z => n2105);
   U694 : CLKBUF_X1 port map( A => n741, Z => n2111);
   U695 : CLKBUF_X1 port map( A => n740, Z => n2117);
   U696 : CLKBUF_X1 port map( A => n739, Z => n2123);
   U697 : CLKBUF_X1 port map( A => n738, Z => n2129);
   U698 : CLKBUF_X1 port map( A => n736, Z => n2135);
   U699 : CLKBUF_X1 port map( A => n735, Z => n2141);
   U700 : CLKBUF_X1 port map( A => n527, Z => n2147);
   U701 : CLKBUF_X1 port map( A => n525, Z => n2158);
   U702 : CLKBUF_X1 port map( A => n523, Z => n2164);
   U703 : CLKBUF_X1 port map( A => n521, Z => n2170);
   U704 : INV_X1 port map( A => ADD_RD2(0), ZN => n2171);
   U705 : INV_X1 port map( A => ADD_RD2(1), ZN => n2172);
   U706 : INV_X1 port map( A => ADD_RD1(0), ZN => n2173);
   U707 : INV_X1 port map( A => ADD_RD1(1), ZN => n2174);
   U708 : INV_X1 port map( A => ADD_WR(0), ZN => n2175);
   U709 : INV_X1 port map( A => ADD_WR(1), ZN => n2176);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4.all;

entity register_file_reg_size64_file_size4_8 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_reg_size64_file_size4_8;

architecture SYN_BEHAVIORAL of register_file_reg_size64_file_size4_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n2, n3, n4, n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19, 
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n174, n175, n176, n177, n178, n179, 
      n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, 
      n192, n415, n1200, n1202, n1204, n1310, n1311, n1312, n1313, n1314, n1315
      , n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, 
      n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, 
      n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, 
      n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, 
      n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, 
      n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, 
      n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, 
      n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, 
      n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, 
      n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, 
      n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, 
      n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, 
      n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, 
      n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, 
      n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, 
      n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, 
      n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, 
      n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, 
      n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, 
      n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, 
      n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, 
      n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, 
      n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, 
      n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, 
      n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, 
      n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, 
      n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, 
      n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, 
      n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, 
      n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, 
      n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, 
      n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, 
      n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, 
      n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, 
      n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, 
      n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, 
      n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, 
      n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, 
      n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, 
      n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, 
      n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, 
      n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, 
      n1736, n1737, n1738, n1793, n1794, n1795, n1796, n1797, n1798, n1799, 
      n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, 
      n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, 
      n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, 
      n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, 
      n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, 
      n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, 
      n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, 
      n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, 
      n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, 
      n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, 
      n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, 
      n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, 
      n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, 
      n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, 
      n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, 
      n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, 
      n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, 
      n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, 
      n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, 
      n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580, 
      n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, 
      n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, 
      n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, 
      n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, 
      n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, 
      n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, 
      n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, 
      n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, 
      n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, 
      n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, 
      n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, 
      n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, 
      n725, n726, n727, n728, n729, n730, n731, n734, n735, n736, n737, n738, 
      n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750, 
      n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, 
      n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774, 
      n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, n786, 
      n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, 
      n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, 
      n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822, 
      n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, 
      n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, 
      n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, 
      n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n871, n872, 
      n873, n875, n876, n936, n938, n939, n975, n978, n979, n998, n999, n1000, 
      n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, 
      n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, 
      n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, 
      n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, 
      n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, 
      n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, 
      n1061, n1062, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, 
      n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, 
      n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, 
      n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, 
      n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, 
      n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, 
      n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, 
      n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, 
      n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, 
      n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, 
      n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, 
      n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, 
      n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, 
      n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, 
      n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, 
      n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, 
      n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, 
      n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, 
      n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, 
      n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, 
      n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, 
      n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, 
      n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176 : std_logic
      ;

begin
   
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1355, CK => CLK, Q => n174,
                           QN => n2028);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1356, CK => CLK, Q => n175,
                           QN => n2027);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1357, CK => CLK, Q => n176,
                           QN => n2026);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1358, CK => CLK, Q => n177,
                           QN => n2025);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1359, CK => CLK, Q => n178,
                           QN => n2024);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1360, CK => CLK, Q => n179,
                           QN => n2023);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1361, CK => CLK, Q => n180,
                           QN => n2022);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1362, CK => CLK, Q => n181,
                           QN => n2021);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1363, CK => CLK, Q => n182,
                           QN => n2020);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1364, CK => CLK, Q => n183, 
                           QN => n2019);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1365, CK => CLK, Q => n184, 
                           QN => n2018);
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n1366, CK => CLK, Q => n185, 
                           QN => n2017);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n1367, CK => CLK, Q => n186, 
                           QN => n2016);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n1368, CK => CLK, Q => n187, 
                           QN => n2015);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n1369, CK => CLK, Q => n188, 
                           QN => n2014);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n1370, CK => CLK, Q => n189, 
                           QN => n2013);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n1371, CK => CLK, Q => n190, 
                           QN => n2012);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n1372, CK => CLK, Q => n191, 
                           QN => n2011);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n1373, CK => CLK, Q => n192, 
                           QN => n2010);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n1374, CK => CLK, Q => n65, 
                           QN => n2063);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n1375, CK => CLK, Q => n66, 
                           QN => n2062);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n1376, CK => CLK, Q => n67, 
                           QN => n2061);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n1377, CK => CLK, Q => n68, 
                           QN => n2060);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n1378, CK => CLK, Q => n69, 
                           QN => n2059);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n1379, CK => CLK, Q => n70, 
                           QN => n2058);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n1380, CK => CLK, Q => n71, 
                           QN => n2057);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n1381, CK => CLK, Q => n72, 
                           QN => n2056);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n1382, CK => CLK, Q => n73, 
                           QN => n2055);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n1383, CK => CLK, Q => n74, 
                           QN => n2054);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n1384, CK => CLK, Q => n75, 
                           QN => n2053);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n1385, CK => CLK, Q => n76, 
                           QN => n2052);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n1386, CK => CLK, Q => n77, 
                           QN => n2051);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n1387, CK => CLK, Q => n78, 
                           QN => n2050);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n1388, CK => CLK, Q => n79, 
                           QN => n2049);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n1389, CK => CLK, Q => n80, 
                           QN => n2048);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n1390, CK => CLK, Q => n81, 
                           QN => n2047);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n1391, CK => CLK, Q => n82, 
                           QN => n2046);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n1392, CK => CLK, Q => n83, 
                           QN => n2045);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n1393, CK => CLK, Q => n84, 
                           QN => n2044);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n1394, CK => CLK, Q => n85, 
                           QN => n2043);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n1395, CK => CLK, Q => n86, 
                           QN => n2042);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n1396, CK => CLK, Q => n87, 
                           QN => n2041);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n1397, CK => CLK, Q => n88, 
                           QN => n2040);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n1398, CK => CLK, Q => n89, 
                           QN => n2039);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n1399, CK => CLK, Q => n90, 
                           QN => n2038);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n1400, CK => CLK, Q => n91, 
                           QN => n2037);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n1401, CK => CLK, Q => n92, 
                           QN => n2036);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n1402, CK => CLK, Q => n93, 
                           QN => n2035);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n1403, CK => CLK, Q => n94, 
                           QN => n2034);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n1404, CK => CLK, Q => n95, 
                           QN => n2033);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n1405, CK => CLK, Q => n96, 
                           QN => n2032);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n1406, CK => CLK, Q => n97, 
                           QN => n2031);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n1407, CK => CLK, Q => n98, 
                           QN => n2030);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n1408, CK => CLK, Q => n99, 
                           QN => n2029);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n1439, CK => CLK, Q => n2, 
                           QN => n2009);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n1440, CK => CLK, Q => n3, 
                           QN => n2008);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n1441, CK => CLK, Q => n4, 
                           QN => n2007);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n1442, CK => CLK, Q => n5, 
                           QN => n2006);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n1443, CK => CLK, Q => n6, 
                           QN => n2005);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n1444, CK => CLK, Q => n7, 
                           QN => n2004);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n1445, CK => CLK, Q => n8, 
                           QN => n2003);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n1446, CK => CLK, Q => n9, 
                           QN => n2002);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n1450, CK => CLK, Q => n13, 
                           QN => n2001);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n1451, CK => CLK, Q => n14, 
                           QN => n2000);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n1452, CK => CLK, Q => n15, 
                           QN => n1999);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n1453, CK => CLK, Q => n16, 
                           QN => n1998);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n1454, CK => CLK, Q => n17, 
                           QN => n1997);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n1455, CK => CLK, Q => n18, 
                           QN => n1996);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n1456, CK => CLK, Q => n19, 
                           QN => n1995);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n1457, CK => CLK, Q => n20, 
                           QN => n1994);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n1458, CK => CLK, Q => n21, 
                           QN => n1993);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n1459, CK => CLK, Q => n22, 
                           QN => n1992);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n1460, CK => CLK, Q => n23, 
                           QN => n1991);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n1461, CK => CLK, Q => n24, 
                           QN => n1990);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n1462, CK => CLK, Q => n25, 
                           QN => n1989);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n1463, CK => CLK, Q => n26, 
                           QN => n1988);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n1464, CK => CLK, Q => n27, 
                           QN => n1987);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n1465, CK => CLK, Q => n28, 
                           QN => n1986);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n1466, CK => CLK, Q => n29, 
                           QN => n1985);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n1467, CK => CLK, Q => n30, 
                           QN => n1984);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n1468, CK => CLK, Q => n31, 
                           QN => n1983);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n1469, CK => CLK, Q => n32, 
                           QN => n1982);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n1470, CK => CLK, Q => n33, 
                           QN => n1981);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n1471, CK => CLK, Q => n34, 
                           QN => n1980);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n1472, CK => CLK, Q => n35, 
                           QN => n1979);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n1473, CK => CLK, Q => n36, 
                           QN => n1978);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n1474, CK => CLK, Q => n37, 
                           QN => n1977);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n1475, CK => CLK, Q => n38, 
                           QN => n1976);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n1476, CK => CLK, Q => n39, 
                           QN => n1975);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n1477, CK => CLK, Q => n40, 
                           QN => n1974);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n1478, CK => CLK, Q => n41, 
                           QN => n1973);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n1479, CK => CLK, Q => n42, 
                           QN => n1972);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n1480, CK => CLK, Q => n43, 
                           QN => n1971);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n1481, CK => CLK, Q => n44, 
                           QN => n1970);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n1482, CK => CLK, Q => n45, 
                           QN => n1969);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n1483, CK => CLK, Q => n46, 
                           QN => n1968);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n1484, CK => CLK, Q => n47, 
                           QN => n1967);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n1485, CK => CLK, Q => n48, 
                           QN => n1966);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n1486, CK => CLK, Q => n49, 
                           QN => n1965);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n1487, CK => CLK, Q => n50, 
                           QN => n1964);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n1488, CK => CLK, Q => n51, 
                           QN => n1963);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n1489, CK => CLK, Q => n52, 
                           QN => n1962);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n1490, CK => CLK, Q => n53, 
                           QN => n1961);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n1491, CK => CLK, Q => n54, 
                           QN => n1960);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n1492, CK => CLK, Q => n55, 
                           QN => n1959);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n1493, CK => CLK, Q => n56, 
                           QN => n1958);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n1494, CK => CLK, Q => n57, 
                           QN => n1957);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n1495, CK => CLK, Q => n58, 
                           QN => n1956);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n1496, CK => CLK, Q => n59, 
                           QN => n1955);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n1497, CK => CLK, Q => n60, 
                           QN => n1954);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n1498, CK => CLK, Q => n61, 
                           QN => n1953);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n1499, CK => CLK, Q => n62, 
                           QN => n1952);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n1500, CK => CLK, Q => n63, 
                           QN => n1951);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n1501, CK => CLK, Q => n64, 
                           QN => n1950);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n1502, CK => CLK, Q => n999,
                           QN => n728);
   OUT2_reg_63_inst : DFF_X1 port map( D => n1503, CK => CLK, Q => OUT2(63), QN
                           => n1822);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n1504, CK => CLK, Q => n1000
                           , QN => n725);
   OUT2_reg_62_inst : DFF_X1 port map( D => n1505, CK => CLK, Q => OUT2(62), QN
                           => n1823);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n1506, CK => CLK, Q => n1001
                           , QN => n722);
   OUT2_reg_61_inst : DFF_X1 port map( D => n1507, CK => CLK, Q => OUT2(61), QN
                           => n1824);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n1508, CK => CLK, Q => n1002
                           , QN => n719);
   OUT2_reg_60_inst : DFF_X1 port map( D => n1509, CK => CLK, Q => OUT2(60), QN
                           => n1825);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n1510, CK => CLK, Q => n1003
                           , QN => n716);
   OUT2_reg_59_inst : DFF_X1 port map( D => n1511, CK => CLK, Q => OUT2(59), QN
                           => n1826);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n1512, CK => CLK, Q => n1004
                           , QN => n713);
   OUT2_reg_58_inst : DFF_X1 port map( D => n1513, CK => CLK, Q => OUT2(58), QN
                           => n1827);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n1514, CK => CLK, Q => n1005
                           , QN => n710);
   OUT2_reg_57_inst : DFF_X1 port map( D => n1515, CK => CLK, Q => OUT2(57), QN
                           => n1828);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n1516, CK => CLK, Q => n1006
                           , QN => n707);
   OUT2_reg_56_inst : DFF_X1 port map( D => n1517, CK => CLK, Q => OUT2(56), QN
                           => n1829);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n1518, CK => CLK, Q => n1007
                           , QN => n704);
   OUT2_reg_55_inst : DFF_X1 port map( D => n1519, CK => CLK, Q => OUT2(55), QN
                           => n1830);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n1520, CK => CLK, Q => n1008
                           , QN => n700);
   OUT2_reg_54_inst : DFF_X1 port map( D => n1521, CK => CLK, Q => OUT2(54), QN
                           => n1831);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n1522, CK => CLK, Q => n1009
                           , QN => n696);
   OUT2_reg_53_inst : DFF_X1 port map( D => n1523, CK => CLK, Q => OUT2(53), QN
                           => n1832);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n1524, CK => CLK, Q => n1010
                           , QN => n692);
   OUT2_reg_52_inst : DFF_X1 port map( D => n1525, CK => CLK, Q => OUT2(52), QN
                           => n1833);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n1526, CK => CLK, Q => n1011
                           , QN => n689);
   OUT2_reg_51_inst : DFF_X1 port map( D => n1527, CK => CLK, Q => OUT2(51), QN
                           => n1834);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n1528, CK => CLK, Q => n1012
                           , QN => n686);
   OUT2_reg_50_inst : DFF_X1 port map( D => n1529, CK => CLK, Q => OUT2(50), QN
                           => n1835);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n1530, CK => CLK, Q => n1013
                           , QN => n683);
   OUT2_reg_49_inst : DFF_X1 port map( D => n1531, CK => CLK, Q => OUT2(49), QN
                           => n1836);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n1532, CK => CLK, Q => n1014
                           , QN => n680);
   OUT2_reg_48_inst : DFF_X1 port map( D => n1533, CK => CLK, Q => OUT2(48), QN
                           => n1837);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n1534, CK => CLK, Q => n1015
                           , QN => n677);
   OUT2_reg_47_inst : DFF_X1 port map( D => n1535, CK => CLK, Q => OUT2(47), QN
                           => n1838);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n1536, CK => CLK, Q => n1016
                           , QN => n674);
   OUT2_reg_46_inst : DFF_X1 port map( D => n1537, CK => CLK, Q => OUT2(46), QN
                           => n1839);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n1538, CK => CLK, Q => n1017
                           , QN => n671);
   OUT2_reg_45_inst : DFF_X1 port map( D => n1539, CK => CLK, Q => OUT2(45), QN
                           => n1840);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n1540, CK => CLK, Q => n1018
                           , QN => n668);
   OUT2_reg_44_inst : DFF_X1 port map( D => n1541, CK => CLK, Q => OUT2(44), QN
                           => n1841);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n1542, CK => CLK, Q => n1019
                           , QN => n665);
   OUT2_reg_43_inst : DFF_X1 port map( D => n1543, CK => CLK, Q => OUT2(43), QN
                           => n1842);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n1544, CK => CLK, Q => n1020
                           , QN => n662);
   OUT2_reg_42_inst : DFF_X1 port map( D => n1545, CK => CLK, Q => OUT2(42), QN
                           => n1843);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n1546, CK => CLK, Q => n1021
                           , QN => n659);
   OUT2_reg_41_inst : DFF_X1 port map( D => n1547, CK => CLK, Q => OUT2(41), QN
                           => n1844);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n1548, CK => CLK, Q => n1022
                           , QN => n656);
   OUT2_reg_40_inst : DFF_X1 port map( D => n1549, CK => CLK, Q => OUT2(40), QN
                           => n1845);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n1550, CK => CLK, Q => n1023
                           , QN => n653);
   OUT2_reg_39_inst : DFF_X1 port map( D => n1551, CK => CLK, Q => OUT2(39), QN
                           => n1846);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n1552, CK => CLK, Q => n1024
                           , QN => n650);
   OUT2_reg_38_inst : DFF_X1 port map( D => n1553, CK => CLK, Q => OUT2(38), QN
                           => n1847);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n1554, CK => CLK, Q => n1025
                           , QN => n647);
   OUT2_reg_37_inst : DFF_X1 port map( D => n1555, CK => CLK, Q => OUT2(37), QN
                           => n1848);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n1556, CK => CLK, Q => n1026
                           , QN => n644);
   OUT2_reg_36_inst : DFF_X1 port map( D => n1557, CK => CLK, Q => OUT2(36), QN
                           => n1849);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n1558, CK => CLK, Q => n1027
                           , QN => n641);
   OUT2_reg_35_inst : DFF_X1 port map( D => n1559, CK => CLK, Q => OUT2(35), QN
                           => n1850);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n1560, CK => CLK, Q => n1028
                           , QN => n638);
   OUT2_reg_34_inst : DFF_X1 port map( D => n1561, CK => CLK, Q => OUT2(34), QN
                           => n1851);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n1562, CK => CLK, Q => n1029
                           , QN => n635);
   OUT2_reg_33_inst : DFF_X1 port map( D => n1563, CK => CLK, Q => OUT2(33), QN
                           => n1852);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n1564, CK => CLK, Q => n1030
                           , QN => n632);
   OUT2_reg_32_inst : DFF_X1 port map( D => n1565, CK => CLK, Q => OUT2(32), QN
                           => n1853);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n1566, CK => CLK, Q => n1031
                           , QN => n629);
   OUT2_reg_31_inst : DFF_X1 port map( D => n1567, CK => CLK, Q => OUT2(31), QN
                           => n1854);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n1568, CK => CLK, Q => n1032
                           , QN => n626);
   OUT2_reg_30_inst : DFF_X1 port map( D => n1569, CK => CLK, Q => OUT2(30), QN
                           => n1855);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n1570, CK => CLK, Q => n1033
                           , QN => n623);
   OUT2_reg_29_inst : DFF_X1 port map( D => n1571, CK => CLK, Q => OUT2(29), QN
                           => n1856);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n1572, CK => CLK, Q => n1034
                           , QN => n619);
   OUT2_reg_28_inst : DFF_X1 port map( D => n1573, CK => CLK, Q => OUT2(28), QN
                           => n1857);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n1574, CK => CLK, Q => n1035
                           , QN => n615);
   OUT2_reg_27_inst : DFF_X1 port map( D => n1575, CK => CLK, Q => OUT2(27), QN
                           => n1858);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n1576, CK => CLK, Q => n1036
                           , QN => n611);
   OUT2_reg_26_inst : DFF_X1 port map( D => n1577, CK => CLK, Q => OUT2(26), QN
                           => n1859);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n1578, CK => CLK, Q => n1037
                           , QN => n607);
   OUT2_reg_25_inst : DFF_X1 port map( D => n1579, CK => CLK, Q => OUT2(25), QN
                           => n1860);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n1580, CK => CLK, Q => n1038
                           , QN => n603);
   OUT2_reg_24_inst : DFF_X1 port map( D => n1581, CK => CLK, Q => OUT2(24), QN
                           => n1861);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n1582, CK => CLK, Q => n1039
                           , QN => n599);
   OUT2_reg_23_inst : DFF_X1 port map( D => n1583, CK => CLK, Q => OUT2(23), QN
                           => n1862);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n1584, CK => CLK, Q => n1040
                           , QN => n595);
   OUT2_reg_22_inst : DFF_X1 port map( D => n1585, CK => CLK, Q => OUT2(22), QN
                           => n1863);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n1586, CK => CLK, Q => n1041
                           , QN => n591);
   OUT2_reg_21_inst : DFF_X1 port map( D => n1587, CK => CLK, Q => OUT2(21), QN
                           => n1864);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n1588, CK => CLK, Q => n1042
                           , QN => n587);
   OUT2_reg_20_inst : DFF_X1 port map( D => n1589, CK => CLK, Q => OUT2(20), QN
                           => n1865);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n1590, CK => CLK, Q => n1043
                           , QN => n583);
   OUT2_reg_19_inst : DFF_X1 port map( D => n1591, CK => CLK, Q => OUT2(19), QN
                           => n1866);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n1592, CK => CLK, Q => n1044
                           , QN => n580);
   OUT2_reg_18_inst : DFF_X1 port map( D => n1593, CK => CLK, Q => OUT2(18), QN
                           => n1867);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n1594, CK => CLK, Q => n1045
                           , QN => n577);
   OUT2_reg_17_inst : DFF_X1 port map( D => n1595, CK => CLK, Q => OUT2(17), QN
                           => n1868);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n1596, CK => CLK, Q => n1046
                           , QN => n574);
   OUT2_reg_16_inst : DFF_X1 port map( D => n1597, CK => CLK, Q => OUT2(16), QN
                           => n1869);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n1598, CK => CLK, Q => n1047
                           , QN => n571);
   OUT2_reg_15_inst : DFF_X1 port map( D => n1599, CK => CLK, Q => OUT2(15), QN
                           => n1870);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n1600, CK => CLK, Q => n1048
                           , QN => n568);
   OUT2_reg_14_inst : DFF_X1 port map( D => n1601, CK => CLK, Q => OUT2(14), QN
                           => n1871);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n1602, CK => CLK, Q => n1049
                           , QN => n565);
   OUT2_reg_13_inst : DFF_X1 port map( D => n1603, CK => CLK, Q => OUT2(13), QN
                           => n1872);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n1604, CK => CLK, Q => n1050
                           , QN => n562);
   OUT2_reg_12_inst : DFF_X1 port map( D => n1605, CK => CLK, Q => OUT2(12), QN
                           => n1873);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n1606, CK => CLK, Q => n1051
                           , QN => n559);
   OUT2_reg_11_inst : DFF_X1 port map( D => n1607, CK => CLK, Q => OUT2(11), QN
                           => n1874);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n1608, CK => CLK, Q => n1052
                           , QN => n556);
   OUT2_reg_10_inst : DFF_X1 port map( D => n1609, CK => CLK, Q => OUT2(10), QN
                           => n1875);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n1610, CK => CLK, Q => n1053,
                           QN => n553);
   OUT2_reg_9_inst : DFF_X1 port map( D => n1611, CK => CLK, Q => OUT2(9), QN 
                           => n1876);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n1612, CK => CLK, Q => n1054,
                           QN => n550);
   OUT2_reg_8_inst : DFF_X1 port map( D => n1613, CK => CLK, Q => OUT2(8), QN 
                           => n1877);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n1614, CK => CLK, Q => n1055,
                           QN => n547);
   OUT2_reg_7_inst : DFF_X1 port map( D => n1615, CK => CLK, Q => OUT2(7), QN 
                           => n1878);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n1616, CK => CLK, Q => n1056,
                           QN => n544);
   OUT2_reg_6_inst : DFF_X1 port map( D => n1617, CK => CLK, Q => OUT2(6), QN 
                           => n1879);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n1618, CK => CLK, Q => n1057,
                           QN => n541);
   OUT2_reg_5_inst : DFF_X1 port map( D => n1619, CK => CLK, Q => OUT2(5), QN 
                           => n1880);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n1620, CK => CLK, Q => n1058,
                           QN => n538);
   OUT2_reg_4_inst : DFF_X1 port map( D => n1621, CK => CLK, Q => OUT2(4), QN 
                           => n1881);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n1622, CK => CLK, Q => n1059,
                           QN => n535);
   OUT2_reg_3_inst : DFF_X1 port map( D => n1623, CK => CLK, Q => OUT2(3), QN 
                           => n1882);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n1624, CK => CLK, Q => n1060,
                           QN => n532);
   OUT2_reg_2_inst : DFF_X1 port map( D => n1625, CK => CLK, Q => OUT2(2), QN 
                           => n1883);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n1626, CK => CLK, Q => n1061,
                           QN => n529);
   OUT2_reg_1_inst : DFF_X1 port map( D => n1627, CK => CLK, Q => OUT2(1), QN 
                           => n1884);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n1628, CK => CLK, Q => n1062,
                           QN => n522);
   OUT2_reg_0_inst : DFF_X1 port map( D => n1629, CK => CLK, Q => OUT2(0), QN 
                           => n1885);
   OUT1_reg_63_inst : DFF_X1 port map( D => n1630, CK => CLK, Q => OUT1(63), QN
                           => n1886);
   OUT1_reg_62_inst : DFF_X1 port map( D => n1631, CK => CLK, Q => OUT1(62), QN
                           => n1887);
   OUT1_reg_61_inst : DFF_X1 port map( D => n1632, CK => CLK, Q => OUT1(61), QN
                           => n1888);
   OUT1_reg_60_inst : DFF_X1 port map( D => n1633, CK => CLK, Q => OUT1(60), QN
                           => n1889);
   OUT1_reg_59_inst : DFF_X1 port map( D => n1634, CK => CLK, Q => OUT1(59), QN
                           => n1890);
   OUT1_reg_58_inst : DFF_X1 port map( D => n1635, CK => CLK, Q => OUT1(58), QN
                           => n1891);
   OUT1_reg_57_inst : DFF_X1 port map( D => n1636, CK => CLK, Q => OUT1(57), QN
                           => n1892);
   OUT1_reg_56_inst : DFF_X1 port map( D => n1637, CK => CLK, Q => OUT1(56), QN
                           => n1893);
   OUT1_reg_55_inst : DFF_X1 port map( D => n1638, CK => CLK, Q => OUT1(55), QN
                           => n1894);
   OUT1_reg_54_inst : DFF_X1 port map( D => n1639, CK => CLK, Q => OUT1(54), QN
                           => n1895);
   OUT1_reg_53_inst : DFF_X1 port map( D => n1640, CK => CLK, Q => OUT1(53), QN
                           => n1896);
   OUT1_reg_52_inst : DFF_X1 port map( D => n1641, CK => CLK, Q => OUT1(52), QN
                           => n1897);
   OUT1_reg_51_inst : DFF_X1 port map( D => n1642, CK => CLK, Q => OUT1(51), QN
                           => n1898);
   OUT1_reg_50_inst : DFF_X1 port map( D => n1643, CK => CLK, Q => OUT1(50), QN
                           => n1899);
   OUT1_reg_49_inst : DFF_X1 port map( D => n1644, CK => CLK, Q => OUT1(49), QN
                           => n1900);
   OUT1_reg_48_inst : DFF_X1 port map( D => n1645, CK => CLK, Q => OUT1(48), QN
                           => n1901);
   OUT1_reg_47_inst : DFF_X1 port map( D => n1646, CK => CLK, Q => OUT1(47), QN
                           => n1902);
   OUT1_reg_46_inst : DFF_X1 port map( D => n1647, CK => CLK, Q => OUT1(46), QN
                           => n1903);
   OUT1_reg_45_inst : DFF_X1 port map( D => n1648, CK => CLK, Q => OUT1(45), QN
                           => n1904);
   OUT1_reg_44_inst : DFF_X1 port map( D => n1649, CK => CLK, Q => OUT1(44), QN
                           => n1905);
   OUT1_reg_43_inst : DFF_X1 port map( D => n1650, CK => CLK, Q => OUT1(43), QN
                           => n1906);
   OUT1_reg_42_inst : DFF_X1 port map( D => n1651, CK => CLK, Q => OUT1(42), QN
                           => n1907);
   OUT1_reg_41_inst : DFF_X1 port map( D => n1652, CK => CLK, Q => OUT1(41), QN
                           => n1908);
   OUT1_reg_40_inst : DFF_X1 port map( D => n1653, CK => CLK, Q => OUT1(40), QN
                           => n1909);
   OUT1_reg_39_inst : DFF_X1 port map( D => n1654, CK => CLK, Q => OUT1(39), QN
                           => n1910);
   OUT1_reg_38_inst : DFF_X1 port map( D => n1655, CK => CLK, Q => OUT1(38), QN
                           => n1911);
   OUT1_reg_37_inst : DFF_X1 port map( D => n1656, CK => CLK, Q => OUT1(37), QN
                           => n1912);
   OUT1_reg_36_inst : DFF_X1 port map( D => n1657, CK => CLK, Q => OUT1(36), QN
                           => n1913);
   OUT1_reg_35_inst : DFF_X1 port map( D => n1658, CK => CLK, Q => OUT1(35), QN
                           => n1914);
   OUT1_reg_34_inst : DFF_X1 port map( D => n1659, CK => CLK, Q => OUT1(34), QN
                           => n1915);
   OUT1_reg_33_inst : DFF_X1 port map( D => n1660, CK => CLK, Q => OUT1(33), QN
                           => n1916);
   OUT1_reg_32_inst : DFF_X1 port map( D => n1661, CK => CLK, Q => OUT1(32), QN
                           => n1917);
   OUT1_reg_31_inst : DFF_X1 port map( D => n1662, CK => CLK, Q => OUT1(31), QN
                           => n1918);
   OUT1_reg_30_inst : DFF_X1 port map( D => n1663, CK => CLK, Q => OUT1(30), QN
                           => n1919);
   OUT1_reg_29_inst : DFF_X1 port map( D => n1664, CK => CLK, Q => OUT1(29), QN
                           => n1920);
   OUT1_reg_28_inst : DFF_X1 port map( D => n1665, CK => CLK, Q => OUT1(28), QN
                           => n1921);
   OUT1_reg_27_inst : DFF_X1 port map( D => n1666, CK => CLK, Q => OUT1(27), QN
                           => n1922);
   OUT1_reg_26_inst : DFF_X1 port map( D => n1667, CK => CLK, Q => OUT1(26), QN
                           => n1923);
   OUT1_reg_25_inst : DFF_X1 port map( D => n1668, CK => CLK, Q => OUT1(25), QN
                           => n1924);
   OUT1_reg_24_inst : DFF_X1 port map( D => n1669, CK => CLK, Q => OUT1(24), QN
                           => n1925);
   OUT1_reg_23_inst : DFF_X1 port map( D => n1670, CK => CLK, Q => OUT1(23), QN
                           => n1926);
   OUT1_reg_22_inst : DFF_X1 port map( D => n1671, CK => CLK, Q => OUT1(22), QN
                           => n1927);
   OUT1_reg_21_inst : DFF_X1 port map( D => n1672, CK => CLK, Q => OUT1(21), QN
                           => n1928);
   OUT1_reg_20_inst : DFF_X1 port map( D => n1673, CK => CLK, Q => OUT1(20), QN
                           => n1929);
   OUT1_reg_19_inst : DFF_X1 port map( D => n1674, CK => CLK, Q => OUT1(19), QN
                           => n1930);
   OUT1_reg_18_inst : DFF_X1 port map( D => n1675, CK => CLK, Q => OUT1(18), QN
                           => n1931);
   OUT1_reg_17_inst : DFF_X1 port map( D => n1676, CK => CLK, Q => OUT1(17), QN
                           => n1932);
   OUT1_reg_16_inst : DFF_X1 port map( D => n1677, CK => CLK, Q => OUT1(16), QN
                           => n1933);
   OUT1_reg_15_inst : DFF_X1 port map( D => n1678, CK => CLK, Q => OUT1(15), QN
                           => n1934);
   OUT1_reg_14_inst : DFF_X1 port map( D => n1679, CK => CLK, Q => OUT1(14), QN
                           => n1935);
   OUT1_reg_13_inst : DFF_X1 port map( D => n1680, CK => CLK, Q => OUT1(13), QN
                           => n1936);
   OUT1_reg_12_inst : DFF_X1 port map( D => n1681, CK => CLK, Q => OUT1(12), QN
                           => n1937);
   OUT1_reg_11_inst : DFF_X1 port map( D => n1682, CK => CLK, Q => OUT1(11), QN
                           => n1938);
   OUT1_reg_10_inst : DFF_X1 port map( D => n1683, CK => CLK, Q => OUT1(10), QN
                           => n1939);
   OUT1_reg_9_inst : DFF_X1 port map( D => n1684, CK => CLK, Q => OUT1(9), QN 
                           => n1940);
   OUT1_reg_8_inst : DFF_X1 port map( D => n1685, CK => CLK, Q => OUT1(8), QN 
                           => n1941);
   OUT1_reg_7_inst : DFF_X1 port map( D => n1686, CK => CLK, Q => OUT1(7), QN 
                           => n1942);
   OUT1_reg_6_inst : DFF_X1 port map( D => n1687, CK => CLK, Q => OUT1(6), QN 
                           => n1943);
   OUT1_reg_5_inst : DFF_X1 port map( D => n1688, CK => CLK, Q => OUT1(5), QN 
                           => n1944);
   OUT1_reg_4_inst : DFF_X1 port map( D => n1689, CK => CLK, Q => OUT1(4), QN 
                           => n1945);
   OUT1_reg_3_inst : DFF_X1 port map( D => n1690, CK => CLK, Q => OUT1(3), QN 
                           => n1946);
   OUT1_reg_2_inst : DFF_X1 port map( D => n1691, CK => CLK, Q => OUT1(2), QN 
                           => n1947);
   OUT1_reg_1_inst : DFF_X1 port map( D => n1692, CK => CLK, Q => OUT1(1), QN 
                           => n1948);
   OUT1_reg_0_inst : DFF_X1 port map( D => n1693, CK => CLK, Q => OUT1(0), QN 
                           => n1949);
   U859 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n2164, A3 => ADD_RD1(1), 
                           ZN => n521);
   U860 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n2135, A3 => ADD_RD2(1), 
                           ZN => n735);
   U861 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n873, A3 => ADD_WR(1), ZN 
                           => n872);
   U862 : NAND3_X1 port map( A1 => n873, A2 => n2175, A3 => ADD_WR(1), ZN => 
                           n936);
   U863 : NAND3_X1 port map( A1 => n873, A2 => n2176, A3 => ADD_WR(0), ZN => 
                           n975);
   U864 : NAND3_X1 port map( A1 => n2175, A2 => n2176, A3 => n873, ZN => n998);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n1434, CK => CLK, Q => n537, 
                           QN => n1818);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n1435, CK => CLK, Q => n534, 
                           QN => n1819);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n1436, CK => CLK, Q => n531, 
                           QN => n1820);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n1437, CK => CLK, Q => n528, 
                           QN => n1821);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n1438, CK => CLK, Q => n730,
                           QN => n415);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n1447, CK => CLK, Q => n702,
                           QN => n1200);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n1448, CK => CLK, Q => n698,
                           QN => n1202);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n1449, CK => CLK, Q => n694,
                           QN => n1204);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n1409, CK => CLK, Q => n622,
                           QN => n1793);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n1410, CK => CLK, Q => n618,
                           QN => n1794);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n1411, CK => CLK, Q => n614,
                           QN => n1795);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n1412, CK => CLK, Q => n610,
                           QN => n1796);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n1413, CK => CLK, Q => n606,
                           QN => n1797);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n1414, CK => CLK, Q => n602,
                           QN => n1798);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n1415, CK => CLK, Q => n598,
                           QN => n1799);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n1416, CK => CLK, Q => n594,
                           QN => n1800);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n1417, CK => CLK, Q => n590,
                           QN => n1801);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n1418, CK => CLK, Q => n586,
                           QN => n1802);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n1419, CK => CLK, Q => n582,
                           QN => n1803);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n1420, CK => CLK, Q => n579,
                           QN => n1804);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n1421, CK => CLK, Q => n576,
                           QN => n1805);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n1422, CK => CLK, Q => n573,
                           QN => n1806);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n1423, CK => CLK, Q => n570,
                           QN => n1807);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n1424, CK => CLK, Q => n567,
                           QN => n1808);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n1425, CK => CLK, Q => n564,
                           QN => n1809);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n1426, CK => CLK, Q => n561,
                           QN => n1810);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n1427, CK => CLK, Q => n558,
                           QN => n1811);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n1428, CK => CLK, Q => n555, 
                           QN => n1812);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n1429, CK => CLK, Q => n552, 
                           QN => n1813);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n1430, CK => CLK, Q => n549, 
                           QN => n1814);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n1431, CK => CLK, Q => n546, 
                           QN => n1815);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n1432, CK => CLK, Q => n543, 
                           QN => n1816);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n1433, CK => CLK, Q => n540, 
                           QN => n1817);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n1310, CK => CLK, Q => n731,
                           QN => n1694);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n1311, CK => CLK, Q => n727,
                           QN => n1695);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n1312, CK => CLK, Q => n724,
                           QN => n1696);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n1313, CK => CLK, Q => n721,
                           QN => n1697);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n1314, CK => CLK, Q => n718,
                           QN => n1698);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n1315, CK => CLK, Q => n715,
                           QN => n1699);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n1316, CK => CLK, Q => n712,
                           QN => n1700);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n1317, CK => CLK, Q => n709,
                           QN => n1701);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n1318, CK => CLK, Q => n706,
                           QN => n1702);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n1319, CK => CLK, Q => n703,
                           QN => n1703);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n1320, CK => CLK, Q => n699,
                           QN => n1704);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n1321, CK => CLK, Q => n695,
                           QN => n1705);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n1322, CK => CLK, Q => n691,
                           QN => n1706);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n1323, CK => CLK, Q => n688,
                           QN => n1707);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n1324, CK => CLK, Q => n685,
                           QN => n1708);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n1325, CK => CLK, Q => n682,
                           QN => n1709);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n1326, CK => CLK, Q => n679,
                           QN => n1710);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n1327, CK => CLK, Q => n676,
                           QN => n1711);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n1328, CK => CLK, Q => n673,
                           QN => n1712);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n1329, CK => CLK, Q => n670,
                           QN => n1713);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n1330, CK => CLK, Q => n667,
                           QN => n1714);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n1331, CK => CLK, Q => n664,
                           QN => n1715);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n1332, CK => CLK, Q => n661,
                           QN => n1716);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n1333, CK => CLK, Q => n658,
                           QN => n1717);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n1334, CK => CLK, Q => n655,
                           QN => n1718);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n1335, CK => CLK, Q => n652,
                           QN => n1719);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n1336, CK => CLK, Q => n649,
                           QN => n1720);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n1337, CK => CLK, Q => n646,
                           QN => n1721);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n1338, CK => CLK, Q => n643,
                           QN => n1722);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n1339, CK => CLK, Q => n640,
                           QN => n1723);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n1340, CK => CLK, Q => n637,
                           QN => n1724);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n1341, CK => CLK, Q => n634,
                           QN => n1725);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1342, CK => CLK, Q => n631,
                           QN => n1726);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1343, CK => CLK, Q => n628,
                           QN => n1727);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1344, CK => CLK, Q => n625,
                           QN => n1728);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1345, CK => CLK, Q => n621,
                           QN => n1729);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1346, CK => CLK, Q => n617,
                           QN => n1730);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1347, CK => CLK, Q => n613,
                           QN => n1731);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1348, CK => CLK, Q => n609,
                           QN => n1732);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1349, CK => CLK, Q => n605,
                           QN => n1733);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1350, CK => CLK, Q => n601,
                           QN => n1734);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1351, CK => CLK, Q => n597,
                           QN => n1735);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1352, CK => CLK, Q => n593,
                           QN => n1736);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1353, CK => CLK, Q => n589,
                           QN => n1737);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1354, CK => CLK, Q => n585,
                           QN => n1738);
   U3 : BUF_X1 port map( A => n521, Z => n2167);
   U4 : BUF_X1 port map( A => n521, Z => n2166);
   U5 : BUF_X1 port map( A => n521, Z => n2165);
   U6 : BUF_X1 port map( A => n735, Z => n2139);
   U7 : BUF_X1 port map( A => n735, Z => n2138);
   U8 : BUF_X1 port map( A => n735, Z => n2137);
   U9 : BUF_X1 port map( A => n735, Z => n2136);
   U10 : BUF_X1 port map( A => n521, Z => n2169);
   U11 : BUF_X1 port map( A => n521, Z => n2168);
   U12 : BUF_X1 port map( A => n735, Z => n2140);
   U13 : BUF_X1 port map( A => n526, Z => n2151);
   U14 : BUF_X1 port map( A => n526, Z => n2152);
   U15 : BUF_X1 port map( A => n527, Z => n2144);
   U16 : BUF_X1 port map( A => n527, Z => n2146);
   U17 : BUF_X1 port map( A => n527, Z => n2145);
   U18 : BUF_X1 port map( A => n523, Z => n2159);
   U19 : BUF_X1 port map( A => n523, Z => n2160);
   U20 : BUF_X1 port map( A => n523, Z => n2161);
   U21 : BUF_X1 port map( A => n523, Z => n2162);
   U22 : BUF_X1 port map( A => n523, Z => n2163);
   U23 : BUF_X1 port map( A => n736, Z => n2130);
   U24 : BUF_X1 port map( A => n736, Z => n2131);
   U25 : BUF_X1 port map( A => n736, Z => n2132);
   U26 : BUF_X1 port map( A => n736, Z => n2133);
   U27 : BUF_X1 port map( A => n736, Z => n2134);
   U28 : BUF_X1 port map( A => n525, Z => n2154);
   U29 : BUF_X1 port map( A => n525, Z => n2155);
   U30 : BUF_X1 port map( A => n525, Z => n2156);
   U31 : BUF_X1 port map( A => n525, Z => n2157);
   U32 : BUF_X1 port map( A => n738, Z => n2128);
   U33 : BUF_X1 port map( A => n738, Z => n2127);
   U34 : BUF_X1 port map( A => n738, Z => n2126);
   U35 : BUF_X1 port map( A => n738, Z => n2125);
   U36 : BUF_X1 port map( A => n738, Z => n2124);
   U37 : BUF_X1 port map( A => n742, Z => n2104);
   U38 : BUF_X1 port map( A => n742, Z => n2103);
   U39 : BUF_X1 port map( A => n742, Z => n2102);
   U40 : BUF_X1 port map( A => n742, Z => n2101);
   U41 : BUF_X1 port map( A => n739, Z => n2122);
   U42 : BUF_X1 port map( A => n739, Z => n2121);
   U43 : BUF_X1 port map( A => n739, Z => n2120);
   U44 : BUF_X1 port map( A => n739, Z => n2119);
   U45 : BUF_X1 port map( A => n739, Z => n2118);
   U46 : BUF_X1 port map( A => n740, Z => n2116);
   U47 : BUF_X1 port map( A => n740, Z => n2115);
   U48 : BUF_X1 port map( A => n740, Z => n2114);
   U49 : BUF_X1 port map( A => n740, Z => n2113);
   U50 : BUF_X1 port map( A => n740, Z => n2112);
   U51 : BUF_X1 port map( A => n741, Z => n2106);
   U52 : BUF_X1 port map( A => n875, Z => n2094);
   U53 : BUF_X1 port map( A => n938, Z => n2082);
   U54 : BUF_X1 port map( A => n978, Z => n2070);
   U55 : BUF_X1 port map( A => n741, Z => n2110);
   U56 : BUF_X1 port map( A => n741, Z => n2109);
   U57 : BUF_X1 port map( A => n741, Z => n2108);
   U58 : BUF_X1 port map( A => n741, Z => n2107);
   U59 : BUF_X1 port map( A => n875, Z => n2098);
   U60 : BUF_X1 port map( A => n875, Z => n2097);
   U61 : BUF_X1 port map( A => n875, Z => n2096);
   U62 : BUF_X1 port map( A => n875, Z => n2095);
   U63 : BUF_X1 port map( A => n938, Z => n2086);
   U64 : BUF_X1 port map( A => n938, Z => n2085);
   U65 : BUF_X1 port map( A => n938, Z => n2084);
   U66 : BUF_X1 port map( A => n938, Z => n2083);
   U67 : BUF_X1 port map( A => n978, Z => n2074);
   U68 : BUF_X1 port map( A => n978, Z => n2073);
   U69 : BUF_X1 port map( A => n978, Z => n2072);
   U70 : BUF_X1 port map( A => n978, Z => n2071);
   U71 : BUF_X1 port map( A => n526, Z => n2148);
   U72 : BUF_X1 port map( A => n526, Z => n2150);
   U73 : BUF_X1 port map( A => n876, Z => n2092);
   U74 : BUF_X1 port map( A => n876, Z => n2091);
   U75 : BUF_X1 port map( A => n876, Z => n2090);
   U76 : BUF_X1 port map( A => n876, Z => n2089);
   U77 : BUF_X1 port map( A => n876, Z => n2088);
   U78 : BUF_X1 port map( A => n939, Z => n2080);
   U79 : BUF_X1 port map( A => n939, Z => n2079);
   U80 : BUF_X1 port map( A => n939, Z => n2078);
   U81 : BUF_X1 port map( A => n939, Z => n2077);
   U82 : BUF_X1 port map( A => n939, Z => n2076);
   U83 : BUF_X1 port map( A => n979, Z => n2068);
   U84 : BUF_X1 port map( A => n979, Z => n2067);
   U85 : BUF_X1 port map( A => n979, Z => n2066);
   U86 : BUF_X1 port map( A => n979, Z => n2065);
   U87 : BUF_X1 port map( A => n979, Z => n2064);
   U88 : BUF_X1 port map( A => n527, Z => n2143);
   U89 : BUF_X1 port map( A => n527, Z => n2142);
   U90 : BUF_X1 port map( A => n526, Z => n2149);
   U91 : BUF_X1 port map( A => n525, Z => n2153);
   U92 : BUF_X1 port map( A => n742, Z => n2100);
   U93 : NAND2_X1 port map( A1 => n734, A2 => n872, ZN => n741);
   U94 : NAND2_X1 port map( A1 => n734, A2 => n936, ZN => n875);
   U95 : NAND2_X1 port map( A1 => n734, A2 => n2094, ZN => n876);
   U96 : NAND2_X1 port map( A1 => n734, A2 => n975, ZN => n938);
   U97 : NAND2_X1 port map( A1 => n734, A2 => n2082, ZN => n939);
   U98 : NAND2_X1 port map( A1 => n734, A2 => n998, ZN => n978);
   U99 : NAND2_X1 port map( A1 => n734, A2 => n2070, ZN => n979);
   U100 : OAI22_X1 port map( A1 => n538, A2 => n2111, B1 => n2104, B2 => n751, 
                           ZN => n1620);
   U101 : OAI22_X1 port map( A1 => n541, A2 => n2110, B1 => n2104, B2 => n753, 
                           ZN => n1618);
   U102 : OAI22_X1 port map( A1 => n544, A2 => n2110, B1 => n2104, B2 => n755, 
                           ZN => n1616);
   U103 : OAI22_X1 port map( A1 => n547, A2 => n2110, B1 => n2104, B2 => n757, 
                           ZN => n1614);
   U104 : OAI22_X1 port map( A1 => n550, A2 => n2110, B1 => n2104, B2 => n759, 
                           ZN => n1612);
   U105 : OAI22_X1 port map( A1 => n553, A2 => n2110, B1 => n2104, B2 => n761, 
                           ZN => n1610);
   U106 : OAI22_X1 port map( A1 => n556, A2 => n2110, B1 => n2104, B2 => n763, 
                           ZN => n1608);
   U107 : OAI22_X1 port map( A1 => n559, A2 => n2110, B1 => n2104, B2 => n765, 
                           ZN => n1606);
   U108 : OAI22_X1 port map( A1 => n562, A2 => n2110, B1 => n2104, B2 => n767, 
                           ZN => n1604);
   U109 : OAI22_X1 port map( A1 => n565, A2 => n2110, B1 => n2104, B2 => n769, 
                           ZN => n1602);
   U110 : OAI22_X1 port map( A1 => n568, A2 => n2110, B1 => n2104, B2 => n771, 
                           ZN => n1600);
   U111 : OAI22_X1 port map( A1 => n571, A2 => n2110, B1 => n2104, B2 => n773, 
                           ZN => n1598);
   U112 : OAI22_X1 port map( A1 => n574, A2 => n2110, B1 => n2103, B2 => n775, 
                           ZN => n1596);
   U113 : OAI22_X1 port map( A1 => n577, A2 => n2109, B1 => n2103, B2 => n777, 
                           ZN => n1594);
   U114 : OAI22_X1 port map( A1 => n580, A2 => n2109, B1 => n2103, B2 => n779, 
                           ZN => n1592);
   U115 : OAI22_X1 port map( A1 => n583, A2 => n2109, B1 => n2103, B2 => n781, 
                           ZN => n1590);
   U116 : OAI22_X1 port map( A1 => n587, A2 => n2109, B1 => n2103, B2 => n783, 
                           ZN => n1588);
   U117 : OAI22_X1 port map( A1 => n591, A2 => n2109, B1 => n2103, B2 => n785, 
                           ZN => n1586);
   U118 : OAI22_X1 port map( A1 => n595, A2 => n2109, B1 => n2103, B2 => n787, 
                           ZN => n1584);
   U119 : OAI22_X1 port map( A1 => n599, A2 => n2109, B1 => n2103, B2 => n789, 
                           ZN => n1582);
   U120 : OAI22_X1 port map( A1 => n603, A2 => n2109, B1 => n2103, B2 => n791, 
                           ZN => n1580);
   U121 : OAI22_X1 port map( A1 => n607, A2 => n2109, B1 => n2103, B2 => n793, 
                           ZN => n1578);
   U122 : OAI22_X1 port map( A1 => n611, A2 => n2109, B1 => n2103, B2 => n795, 
                           ZN => n1576);
   U123 : OAI22_X1 port map( A1 => n615, A2 => n2109, B1 => n2103, B2 => n797, 
                           ZN => n1574);
   U124 : OAI22_X1 port map( A1 => n619, A2 => n2109, B1 => n2102, B2 => n799, 
                           ZN => n1572);
   U125 : OAI22_X1 port map( A1 => n623, A2 => n2108, B1 => n2102, B2 => n801, 
                           ZN => n1570);
   U126 : OAI22_X1 port map( A1 => n626, A2 => n2108, B1 => n2102, B2 => n803, 
                           ZN => n1568);
   U127 : OAI22_X1 port map( A1 => n629, A2 => n2108, B1 => n2102, B2 => n805, 
                           ZN => n1566);
   U128 : OAI22_X1 port map( A1 => n632, A2 => n2108, B1 => n2102, B2 => n807, 
                           ZN => n1564);
   U129 : OAI22_X1 port map( A1 => n635, A2 => n2108, B1 => n2102, B2 => n809, 
                           ZN => n1562);
   U130 : OAI22_X1 port map( A1 => n638, A2 => n2108, B1 => n2102, B2 => n811, 
                           ZN => n1560);
   U131 : OAI22_X1 port map( A1 => n641, A2 => n2108, B1 => n2102, B2 => n813, 
                           ZN => n1558);
   U132 : OAI22_X1 port map( A1 => n644, A2 => n2108, B1 => n2102, B2 => n815, 
                           ZN => n1556);
   U133 : OAI22_X1 port map( A1 => n647, A2 => n2108, B1 => n2102, B2 => n817, 
                           ZN => n1554);
   U134 : OAI22_X1 port map( A1 => n650, A2 => n2108, B1 => n2102, B2 => n819, 
                           ZN => n1552);
   U135 : OAI22_X1 port map( A1 => n653, A2 => n2108, B1 => n2102, B2 => n821, 
                           ZN => n1550);
   U136 : OAI22_X1 port map( A1 => n656, A2 => n2108, B1 => n2101, B2 => n823, 
                           ZN => n1548);
   U137 : OAI22_X1 port map( A1 => n659, A2 => n2107, B1 => n2101, B2 => n825, 
                           ZN => n1546);
   U138 : OAI22_X1 port map( A1 => n662, A2 => n2107, B1 => n2101, B2 => n827, 
                           ZN => n1544);
   U139 : OAI22_X1 port map( A1 => n665, A2 => n2107, B1 => n2101, B2 => n829, 
                           ZN => n1542);
   U140 : OAI22_X1 port map( A1 => n668, A2 => n2107, B1 => n2101, B2 => n831, 
                           ZN => n1540);
   U141 : OAI22_X1 port map( A1 => n671, A2 => n2107, B1 => n2101, B2 => n833, 
                           ZN => n1538);
   U142 : OAI22_X1 port map( A1 => n674, A2 => n2107, B1 => n2101, B2 => n835, 
                           ZN => n1536);
   U143 : OAI22_X1 port map( A1 => n677, A2 => n2107, B1 => n2101, B2 => n837, 
                           ZN => n1534);
   U144 : OAI22_X1 port map( A1 => n680, A2 => n2107, B1 => n2101, B2 => n839, 
                           ZN => n1532);
   U145 : OAI22_X1 port map( A1 => n683, A2 => n2107, B1 => n2101, B2 => n841, 
                           ZN => n1530);
   U146 : OAI22_X1 port map( A1 => n686, A2 => n2107, B1 => n2101, B2 => n843, 
                           ZN => n1528);
   U147 : OAI22_X1 port map( A1 => n689, A2 => n2107, B1 => n2101, B2 => n845, 
                           ZN => n1526);
   U148 : OAI22_X1 port map( A1 => n522, A2 => n2111, B1 => n2105, B2 => n743, 
                           ZN => n1628);
   U149 : OAI22_X1 port map( A1 => n529, A2 => n2111, B1 => n2105, B2 => n745, 
                           ZN => n1626);
   U150 : OAI22_X1 port map( A1 => n532, A2 => n2111, B1 => n2105, B2 => n747, 
                           ZN => n1624);
   U151 : OAI22_X1 port map( A1 => n535, A2 => n2111, B1 => n2105, B2 => n749, 
                           ZN => n1622);
   U152 : OAI22_X1 port map( A1 => n692, A2 => n2107, B1 => n2100, B2 => n847, 
                           ZN => n1524);
   U153 : OAI22_X1 port map( A1 => n696, A2 => n2106, B1 => n2100, B2 => n849, 
                           ZN => n1522);
   U154 : OAI22_X1 port map( A1 => n700, A2 => n2106, B1 => n2100, B2 => n851, 
                           ZN => n1520);
   U155 : OAI22_X1 port map( A1 => n704, A2 => n2106, B1 => n2100, B2 => n853, 
                           ZN => n1518);
   U156 : OAI22_X1 port map( A1 => n707, A2 => n2106, B1 => n2100, B2 => n855, 
                           ZN => n1516);
   U157 : OAI22_X1 port map( A1 => n710, A2 => n2106, B1 => n2100, B2 => n857, 
                           ZN => n1514);
   U158 : OAI22_X1 port map( A1 => n713, A2 => n2106, B1 => n2100, B2 => n859, 
                           ZN => n1512);
   U159 : OAI22_X1 port map( A1 => n716, A2 => n2106, B1 => n2100, B2 => n861, 
                           ZN => n1510);
   U160 : OAI22_X1 port map( A1 => n719, A2 => n2106, B1 => n2100, B2 => n863, 
                           ZN => n1508);
   U161 : OAI22_X1 port map( A1 => n722, A2 => n2106, B1 => n2100, B2 => n865, 
                           ZN => n1506);
   U162 : OAI22_X1 port map( A1 => n725, A2 => n2106, B1 => n2100, B2 => n867, 
                           ZN => n1504);
   U163 : OAI22_X1 port map( A1 => n728, A2 => n2106, B1 => n2100, B2 => n871, 
                           ZN => n1502);
   U164 : AND3_X1 port map( A1 => n2173, A2 => n2174, A3 => n2164, ZN => n526);
   U165 : AND3_X1 port map( A1 => n2164, A2 => n2174, A3 => ADD_RD1(0), ZN => 
                           n527);
   U166 : AND3_X1 port map( A1 => n2164, A2 => n2173, A3 => ADD_RD1(1), ZN => 
                           n525);
   U167 : NAND2_X1 port map( A1 => n734, A2 => n2106, ZN => n742);
   U168 : AND3_X1 port map( A1 => n2135, A2 => n2172, A3 => ADD_RD2(0), ZN => 
                           n740);
   U169 : AND3_X1 port map( A1 => n2135, A2 => n2171, A3 => ADD_RD2(1), ZN => 
                           n738);
   U170 : AND3_X1 port map( A1 => n2171, A2 => n2172, A3 => n2135, ZN => n739);
   U171 : AND2_X1 port map( A1 => RD2, A2 => n734, ZN => n736);
   U172 : AND2_X1 port map( A1 => RD1, A2 => n734, ZN => n523);
   U173 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n873);
   U174 : OAI221_X1 port map( B1 => n2169, B2 => n562, C1 => n1937, C2 => n2160
                           , A => n563, ZN => n1681);
   U175 : AOI222_X1 port map( A1 => n52, A2 => n2153, B1 => n180, B2 => n2149, 
                           C1 => n2146, C2 => n564, ZN => n563);
   U176 : OAI221_X1 port map( B1 => n2169, B2 => n565, C1 => n1936, C2 => n2160
                           , A => n566, ZN => n1680);
   U177 : AOI222_X1 port map( A1 => n51, A2 => n2154, B1 => n179, B2 => n2149, 
                           C1 => n2146, C2 => n567, ZN => n566);
   U178 : OAI221_X1 port map( B1 => n2169, B2 => n568, C1 => n1935, C2 => n2160
                           , A => n569, ZN => n1679);
   U179 : AOI222_X1 port map( A1 => n50, A2 => n2154, B1 => n178, B2 => n2149, 
                           C1 => n2146, C2 => n570, ZN => n569);
   U180 : OAI221_X1 port map( B1 => n2169, B2 => n571, C1 => n1934, C2 => n2161
                           , A => n572, ZN => n1678);
   U181 : AOI222_X1 port map( A1 => n49, A2 => n2154, B1 => n177, B2 => n2149, 
                           C1 => n2145, C2 => n573, ZN => n572);
   U182 : OAI221_X1 port map( B1 => n2168, B2 => n574, C1 => n1933, C2 => n2160
                           , A => n575, ZN => n1677);
   U183 : AOI222_X1 port map( A1 => n48, A2 => n2154, B1 => n176, B2 => n2149, 
                           C1 => n2145, C2 => n576, ZN => n575);
   U184 : OAI221_X1 port map( B1 => n2168, B2 => n577, C1 => n1932, C2 => n2160
                           , A => n578, ZN => n1676);
   U185 : AOI222_X1 port map( A1 => n47, A2 => n2154, B1 => n175, B2 => n2149, 
                           C1 => n2145, C2 => n579, ZN => n578);
   U186 : OAI221_X1 port map( B1 => n2168, B2 => n580, C1 => n1931, C2 => n2160
                           , A => n581, ZN => n1675);
   U187 : AOI222_X1 port map( A1 => n46, A2 => n2154, B1 => n174, B2 => n2149, 
                           C1 => n2145, C2 => n582, ZN => n581);
   U188 : OAI221_X1 port map( B1 => n538, B2 => n2140, C1 => n1881, C2 => n2130
                           , A => n750, ZN => n1621);
   U189 : AOI222_X1 port map( A1 => n2128, A2 => n60, B1 => n2122, B2 => n188, 
                           C1 => n2116, C2 => n540, ZN => n750);
   U190 : OAI221_X1 port map( B1 => n541, B2 => n2140, C1 => n1880, C2 => n2130
                           , A => n752, ZN => n1619);
   U191 : AOI222_X1 port map( A1 => n2128, A2 => n59, B1 => n2122, B2 => n187, 
                           C1 => n2116, C2 => n543, ZN => n752);
   U192 : OAI221_X1 port map( B1 => n544, B2 => n2140, C1 => n1879, C2 => n2130
                           , A => n754, ZN => n1617);
   U193 : AOI222_X1 port map( A1 => n2128, A2 => n58, B1 => n2122, B2 => n186, 
                           C1 => n2116, C2 => n546, ZN => n754);
   U194 : OAI221_X1 port map( B1 => n547, B2 => n2140, C1 => n1878, C2 => n2130
                           , A => n756, ZN => n1615);
   U195 : AOI222_X1 port map( A1 => n2128, A2 => n57, B1 => n2122, B2 => n185, 
                           C1 => n2116, C2 => n549, ZN => n756);
   U196 : OAI221_X1 port map( B1 => n550, B2 => n2140, C1 => n1877, C2 => n2130
                           , A => n758, ZN => n1613);
   U197 : AOI222_X1 port map( A1 => n2128, A2 => n56, B1 => n2122, B2 => n184, 
                           C1 => n2116, C2 => n552, ZN => n758);
   U198 : OAI221_X1 port map( B1 => n553, B2 => n2140, C1 => n1876, C2 => n2130
                           , A => n760, ZN => n1611);
   U199 : AOI222_X1 port map( A1 => n2128, A2 => n55, B1 => n2122, B2 => n183, 
                           C1 => n2116, C2 => n555, ZN => n760);
   U200 : OAI221_X1 port map( B1 => n556, B2 => n2140, C1 => n1875, C2 => n2130
                           , A => n762, ZN => n1609);
   U201 : AOI222_X1 port map( A1 => n2128, A2 => n54, B1 => n2122, B2 => n182, 
                           C1 => n2116, C2 => n558, ZN => n762);
   U202 : OAI221_X1 port map( B1 => n559, B2 => n2140, C1 => n1874, C2 => n2130
                           , A => n764, ZN => n1607);
   U203 : AOI222_X1 port map( A1 => n2128, A2 => n53, B1 => n2122, B2 => n181, 
                           C1 => n2116, C2 => n561, ZN => n764);
   U204 : OAI221_X1 port map( B1 => n562, B2 => n2140, C1 => n1873, C2 => n2131
                           , A => n766, ZN => n1605);
   U205 : AOI222_X1 port map( A1 => n2128, A2 => n52, B1 => n2122, B2 => n180, 
                           C1 => n2116, C2 => n564, ZN => n766);
   U206 : OAI221_X1 port map( B1 => n565, B2 => n2140, C1 => n1872, C2 => n2131
                           , A => n768, ZN => n1603);
   U207 : AOI222_X1 port map( A1 => n2128, A2 => n51, B1 => n2122, B2 => n179, 
                           C1 => n2116, C2 => n567, ZN => n768);
   U208 : OAI221_X1 port map( B1 => n568, B2 => n2140, C1 => n1871, C2 => n2131
                           , A => n770, ZN => n1601);
   U209 : AOI222_X1 port map( A1 => n2128, A2 => n50, B1 => n2122, B2 => n178, 
                           C1 => n2116, C2 => n570, ZN => n770);
   U210 : OAI221_X1 port map( B1 => n571, B2 => n2140, C1 => n1870, C2 => n2132
                           , A => n772, ZN => n1599);
   U211 : AOI222_X1 port map( A1 => n2128, A2 => n49, B1 => n2122, B2 => n177, 
                           C1 => n2116, C2 => n573, ZN => n772);
   U212 : OAI221_X1 port map( B1 => n574, B2 => n2139, C1 => n1869, C2 => n2131
                           , A => n774, ZN => n1597);
   U213 : AOI222_X1 port map( A1 => n2127, A2 => n48, B1 => n2121, B2 => n176, 
                           C1 => n2115, C2 => n576, ZN => n774);
   U214 : OAI221_X1 port map( B1 => n577, B2 => n2139, C1 => n1868, C2 => n2131
                           , A => n776, ZN => n1595);
   U215 : AOI222_X1 port map( A1 => n2127, A2 => n47, B1 => n2121, B2 => n175, 
                           C1 => n2115, C2 => n579, ZN => n776);
   U216 : OAI221_X1 port map( B1 => n580, B2 => n2139, C1 => n1867, C2 => n2131
                           , A => n778, ZN => n1593);
   U217 : AOI222_X1 port map( A1 => n2127, A2 => n46, B1 => n2121, B2 => n174, 
                           C1 => n2115, C2 => n582, ZN => n778);
   U218 : OAI221_X1 port map( B1 => n2165, B2 => n716, C1 => n1890, C2 => n2164
                           , A => n717, ZN => n1634);
   U219 : AOI222_X1 port map( A1 => n5, A2 => n2157, B1 => n2152, B2 => n718, 
                           C1 => n69, C2 => n2142, ZN => n717);
   U220 : OAI221_X1 port map( B1 => n2165, B2 => n722, C1 => n1888, C2 => n2164
                           , A => n723, ZN => n1632);
   U221 : AOI222_X1 port map( A1 => n3, A2 => n2157, B1 => n2152, B2 => n724, 
                           C1 => n67, C2 => n2142, ZN => n723);
   U222 : OAI221_X1 port map( B1 => n2165, B2 => n725, C1 => n1887, C2 => n2164
                           , A => n726, ZN => n1631);
   U223 : AOI222_X1 port map( A1 => n2, A2 => n2157, B1 => n2152, B2 => n727, 
                           C1 => n66, C2 => n2142, ZN => n726);
   U224 : OAI221_X1 port map( B1 => n2165, B2 => n728, C1 => n1886, C2 => n2164
                           , A => n729, ZN => n1630);
   U225 : AOI222_X1 port map( A1 => n2158, A2 => n730, B1 => n2150, B2 => n731,
                           C1 => n65, C2 => n2142, ZN => n729);
   U226 : OAI221_X1 port map( B1 => n623, B2 => n2138, C1 => n1856, C2 => n2132
                           , A => n800, ZN => n1571);
   U227 : AOI222_X1 port map( A1 => n2126, A2 => n35, B1 => n2120, B2 => n625, 
                           C1 => n2114, C2 => n99, ZN => n800);
   U228 : OAI221_X1 port map( B1 => n626, B2 => n2138, C1 => n1855, C2 => n2132
                           , A => n802, ZN => n1569);
   U229 : AOI222_X1 port map( A1 => n2126, A2 => n34, B1 => n2120, B2 => n628, 
                           C1 => n2114, C2 => n98, ZN => n802);
   U230 : OAI221_X1 port map( B1 => n629, B2 => n2138, C1 => n1854, C2 => n2132
                           , A => n804, ZN => n1567);
   U231 : AOI222_X1 port map( A1 => n2126, A2 => n33, B1 => n2120, B2 => n631, 
                           C1 => n2114, C2 => n97, ZN => n804);
   U232 : OAI221_X1 port map( B1 => n632, B2 => n2138, C1 => n1853, C2 => n2132
                           , A => n806, ZN => n1565);
   U233 : AOI222_X1 port map( A1 => n2126, A2 => n32, B1 => n2120, B2 => n634, 
                           C1 => n2114, C2 => n96, ZN => n806);
   U234 : OAI221_X1 port map( B1 => n635, B2 => n2138, C1 => n1852, C2 => n2132
                           , A => n808, ZN => n1563);
   U235 : AOI222_X1 port map( A1 => n2126, A2 => n31, B1 => n2120, B2 => n637, 
                           C1 => n2114, C2 => n95, ZN => n808);
   U236 : OAI221_X1 port map( B1 => n638, B2 => n2138, C1 => n1851, C2 => n2132
                           , A => n810, ZN => n1561);
   U237 : AOI222_X1 port map( A1 => n2126, A2 => n30, B1 => n2120, B2 => n640, 
                           C1 => n2114, C2 => n94, ZN => n810);
   U238 : OAI221_X1 port map( B1 => n641, B2 => n2138, C1 => n1850, C2 => n2132
                           , A => n812, ZN => n1559);
   U239 : AOI222_X1 port map( A1 => n2126, A2 => n29, B1 => n2120, B2 => n643, 
                           C1 => n2114, C2 => n93, ZN => n812);
   U240 : OAI221_X1 port map( B1 => n644, B2 => n2138, C1 => n1849, C2 => n2133
                           , A => n814, ZN => n1557);
   U241 : AOI222_X1 port map( A1 => n2126, A2 => n28, B1 => n2120, B2 => n646, 
                           C1 => n2114, C2 => n92, ZN => n814);
   U242 : OAI221_X1 port map( B1 => n647, B2 => n2138, C1 => n1848, C2 => n2133
                           , A => n816, ZN => n1555);
   U243 : AOI222_X1 port map( A1 => n2126, A2 => n27, B1 => n2120, B2 => n649, 
                           C1 => n2114, C2 => n91, ZN => n816);
   U244 : OAI221_X1 port map( B1 => n650, B2 => n2138, C1 => n1847, C2 => n2133
                           , A => n818, ZN => n1553);
   U245 : AOI222_X1 port map( A1 => n2126, A2 => n26, B1 => n2120, B2 => n652, 
                           C1 => n2114, C2 => n90, ZN => n818);
   U246 : OAI221_X1 port map( B1 => n653, B2 => n2138, C1 => n1846, C2 => n2133
                           , A => n820, ZN => n1551);
   U247 : AOI222_X1 port map( A1 => n2126, A2 => n25, B1 => n2120, B2 => n655, 
                           C1 => n2114, C2 => n89, ZN => n820);
   U248 : OAI221_X1 port map( B1 => n656, B2 => n2137, C1 => n1845, C2 => n2133
                           , A => n822, ZN => n1549);
   U249 : AOI222_X1 port map( A1 => n2125, A2 => n24, B1 => n2119, B2 => n658, 
                           C1 => n2113, C2 => n88, ZN => n822);
   U250 : OAI221_X1 port map( B1 => n659, B2 => n2137, C1 => n1844, C2 => n2133
                           , A => n824, ZN => n1547);
   U251 : AOI222_X1 port map( A1 => n2125, A2 => n23, B1 => n2119, B2 => n661, 
                           C1 => n2113, C2 => n87, ZN => n824);
   U252 : OAI221_X1 port map( B1 => n662, B2 => n2137, C1 => n1843, C2 => n2133
                           , A => n826, ZN => n1545);
   U253 : AOI222_X1 port map( A1 => n2125, A2 => n22, B1 => n2119, B2 => n664, 
                           C1 => n2113, C2 => n86, ZN => n826);
   U254 : OAI221_X1 port map( B1 => n665, B2 => n2137, C1 => n1842, C2 => n2133
                           , A => n828, ZN => n1543);
   U255 : AOI222_X1 port map( A1 => n2125, A2 => n21, B1 => n2119, B2 => n667, 
                           C1 => n2113, C2 => n85, ZN => n828);
   U256 : OAI221_X1 port map( B1 => n668, B2 => n2137, C1 => n1841, C2 => n2133
                           , A => n830, ZN => n1541);
   U257 : AOI222_X1 port map( A1 => n2125, A2 => n20, B1 => n2119, B2 => n670, 
                           C1 => n2113, C2 => n84, ZN => n830);
   U258 : OAI221_X1 port map( B1 => n671, B2 => n2137, C1 => n1840, C2 => n2133
                           , A => n832, ZN => n1539);
   U259 : AOI222_X1 port map( A1 => n2125, A2 => n19, B1 => n2119, B2 => n673, 
                           C1 => n2113, C2 => n83, ZN => n832);
   U260 : OAI221_X1 port map( B1 => n674, B2 => n2137, C1 => n1839, C2 => n2133
                           , A => n834, ZN => n1537);
   U261 : AOI222_X1 port map( A1 => n2125, A2 => n18, B1 => n2119, B2 => n676, 
                           C1 => n2113, C2 => n82, ZN => n834);
   U262 : OAI221_X1 port map( B1 => n677, B2 => n2137, C1 => n1838, C2 => n2133
                           , A => n836, ZN => n1535);
   U263 : AOI222_X1 port map( A1 => n2125, A2 => n17, B1 => n2119, B2 => n679, 
                           C1 => n2113, C2 => n81, ZN => n836);
   U264 : OAI221_X1 port map( B1 => n680, B2 => n2137, C1 => n1837, C2 => n2134
                           , A => n838, ZN => n1533);
   U265 : AOI222_X1 port map( A1 => n2125, A2 => n16, B1 => n2119, B2 => n682, 
                           C1 => n2113, C2 => n80, ZN => n838);
   U266 : OAI221_X1 port map( B1 => n683, B2 => n2137, C1 => n1836, C2 => n2134
                           , A => n840, ZN => n1531);
   U267 : AOI222_X1 port map( A1 => n2125, A2 => n15, B1 => n2119, B2 => n685, 
                           C1 => n2113, C2 => n79, ZN => n840);
   U268 : OAI221_X1 port map( B1 => n686, B2 => n2137, C1 => n1835, C2 => n2134
                           , A => n842, ZN => n1529);
   U269 : AOI222_X1 port map( A1 => n2125, A2 => n14, B1 => n2119, B2 => n688, 
                           C1 => n2113, C2 => n78, ZN => n842);
   U270 : OAI221_X1 port map( B1 => n689, B2 => n2137, C1 => n1834, C2 => n2134
                           , A => n844, ZN => n1527);
   U271 : AOI222_X1 port map( A1 => n2125, A2 => n13, B1 => n2119, B2 => n691, 
                           C1 => n2113, C2 => n77, ZN => n844);
   U272 : OAI221_X1 port map( B1 => n692, B2 => n2136, C1 => n1833, C2 => n2134
                           , A => n846, ZN => n1525);
   U273 : AOI222_X1 port map( A1 => n2124, A2 => n694, B1 => n2118, B2 => n695,
                           C1 => n2112, C2 => n76, ZN => n846);
   U274 : OAI221_X1 port map( B1 => n696, B2 => n2136, C1 => n1832, C2 => n2134
                           , A => n848, ZN => n1523);
   U275 : AOI222_X1 port map( A1 => n2124, A2 => n698, B1 => n2118, B2 => n699,
                           C1 => n2112, C2 => n75, ZN => n848);
   U276 : OAI221_X1 port map( B1 => n700, B2 => n2136, C1 => n1831, C2 => n2134
                           , A => n850, ZN => n1521);
   U277 : AOI222_X1 port map( A1 => n2124, A2 => n702, B1 => n2118, B2 => n703,
                           C1 => n2112, C2 => n74, ZN => n850);
   U278 : OAI221_X1 port map( B1 => n704, B2 => n2136, C1 => n1830, C2 => n2134
                           , A => n852, ZN => n1519);
   U279 : AOI222_X1 port map( A1 => n2124, A2 => n9, B1 => n2118, B2 => n706, 
                           C1 => n2112, C2 => n73, ZN => n852);
   U280 : OAI221_X1 port map( B1 => n707, B2 => n2136, C1 => n1829, C2 => n2134
                           , A => n854, ZN => n1517);
   U281 : AOI222_X1 port map( A1 => n2124, A2 => n8, B1 => n2118, B2 => n709, 
                           C1 => n2112, C2 => n72, ZN => n854);
   U282 : OAI221_X1 port map( B1 => n710, B2 => n2136, C1 => n1828, C2 => n2134
                           , A => n856, ZN => n1515);
   U283 : AOI222_X1 port map( A1 => n2124, A2 => n7, B1 => n2118, B2 => n712, 
                           C1 => n2112, C2 => n71, ZN => n856);
   U284 : OAI221_X1 port map( B1 => n713, B2 => n2136, C1 => n1827, C2 => n2134
                           , A => n858, ZN => n1513);
   U285 : AOI222_X1 port map( A1 => n2124, A2 => n6, B1 => n2118, B2 => n715, 
                           C1 => n2112, C2 => n70, ZN => n858);
   U286 : OAI221_X1 port map( B1 => n716, B2 => n2136, C1 => n1826, C2 => n2135
                           , A => n860, ZN => n1511);
   U287 : AOI222_X1 port map( A1 => n2124, A2 => n5, B1 => n2118, B2 => n718, 
                           C1 => n2112, C2 => n69, ZN => n860);
   U288 : OAI221_X1 port map( B1 => n719, B2 => n2136, C1 => n1825, C2 => n2134
                           , A => n862, ZN => n1509);
   U289 : AOI222_X1 port map( A1 => n2124, A2 => n4, B1 => n2118, B2 => n721, 
                           C1 => n2112, C2 => n68, ZN => n862);
   U290 : OAI221_X1 port map( B1 => n722, B2 => n2136, C1 => n1824, C2 => n2135
                           , A => n864, ZN => n1507);
   U291 : AOI222_X1 port map( A1 => n2124, A2 => n3, B1 => n2118, B2 => n724, 
                           C1 => n2112, C2 => n67, ZN => n864);
   U292 : OAI221_X1 port map( B1 => n725, B2 => n2136, C1 => n1823, C2 => n2135
                           , A => n866, ZN => n1505);
   U293 : AOI222_X1 port map( A1 => n2124, A2 => n2, B1 => n2118, B2 => n727, 
                           C1 => n2112, C2 => n66, ZN => n866);
   U294 : OAI221_X1 port map( B1 => n728, B2 => n2136, C1 => n1822, C2 => n2135
                           , A => n868, ZN => n1503);
   U295 : AOI222_X1 port map( A1 => n2124, A2 => n730, B1 => n2118, B2 => n731,
                           C1 => n2112, C2 => n65, ZN => n868);
   U296 : INV_X1 port map( A => RESET, ZN => n734);
   U297 : OAI221_X1 port map( B1 => n2170, B2 => n522, C1 => n1949, C2 => n2159
                           , A => n524, ZN => n1693);
   U298 : AOI222_X1 port map( A1 => n64, A2 => n2155, B1 => n192, B2 => n2148, 
                           C1 => n2147, C2 => n528, ZN => n524);
   U299 : OAI221_X1 port map( B1 => n2170, B2 => n529, C1 => n1948, C2 => n2159
                           , A => n530, ZN => n1692);
   U300 : AOI222_X1 port map( A1 => n63, A2 => n2153, B1 => n191, B2 => n2148, 
                           C1 => n2147, C2 => n531, ZN => n530);
   U301 : OAI221_X1 port map( B1 => n2170, B2 => n532, C1 => n1947, C2 => n2159
                           , A => n533, ZN => n1691);
   U302 : AOI222_X1 port map( A1 => n62, A2 => n2153, B1 => n190, B2 => n2148, 
                           C1 => n2146, C2 => n534, ZN => n533);
   U303 : OAI221_X1 port map( B1 => n2170, B2 => n535, C1 => n1946, C2 => n2159
                           , A => n536, ZN => n1690);
   U304 : AOI222_X1 port map( A1 => n61, A2 => n2153, B1 => n189, B2 => n2148, 
                           C1 => n2146, C2 => n537, ZN => n536);
   U305 : OAI221_X1 port map( B1 => n2167, B2 => n619, C1 => n1921, C2 => n2161
                           , A => n620, ZN => n1665);
   U306 : AOI222_X1 port map( A1 => n36, A2 => n2155, B1 => n2150, B2 => n621, 
                           C1 => n2144, C2 => n622, ZN => n620);
   U307 : OAI221_X1 port map( B1 => n2167, B2 => n623, C1 => n1920, C2 => n2161
                           , A => n624, ZN => n1664);
   U308 : AOI222_X1 port map( A1 => n35, A2 => n2155, B1 => n2150, B2 => n625, 
                           C1 => n99, C2 => n2144, ZN => n624);
   U309 : OAI221_X1 port map( B1 => n2167, B2 => n626, C1 => n1919, C2 => n2161
                           , A => n627, ZN => n1663);
   U310 : AOI222_X1 port map( A1 => n34, A2 => n2155, B1 => n2150, B2 => n628, 
                           C1 => n98, C2 => n2144, ZN => n627);
   U311 : OAI221_X1 port map( B1 => n2167, B2 => n629, C1 => n1918, C2 => n2161
                           , A => n630, ZN => n1662);
   U312 : AOI222_X1 port map( A1 => n33, A2 => n2155, B1 => n2150, B2 => n631, 
                           C1 => n97, C2 => n2144, ZN => n630);
   U313 : OAI221_X1 port map( B1 => n2167, B2 => n632, C1 => n1917, C2 => n2161
                           , A => n633, ZN => n1661);
   U314 : AOI222_X1 port map( A1 => n32, A2 => n2155, B1 => n2150, B2 => n634, 
                           C1 => n96, C2 => n2144, ZN => n633);
   U315 : OAI221_X1 port map( B1 => n2167, B2 => n635, C1 => n1916, C2 => n2161
                           , A => n636, ZN => n1660);
   U316 : AOI222_X1 port map( A1 => n31, A2 => n2155, B1 => n2150, B2 => n637, 
                           C1 => n95, C2 => n2144, ZN => n636);
   U317 : OAI221_X1 port map( B1 => n2167, B2 => n638, C1 => n1915, C2 => n2161
                           , A => n639, ZN => n1659);
   U318 : AOI222_X1 port map( A1 => n30, A2 => n2155, B1 => n2150, B2 => n640, 
                           C1 => n94, C2 => n2144, ZN => n639);
   U319 : OAI221_X1 port map( B1 => n2167, B2 => n641, C1 => n1914, C2 => n2161
                           , A => n642, ZN => n1658);
   U320 : AOI222_X1 port map( A1 => n29, A2 => n2155, B1 => n2150, B2 => n643, 
                           C1 => n93, C2 => n2144, ZN => n642);
   U321 : OAI221_X1 port map( B1 => n2167, B2 => n644, C1 => n1913, C2 => n2162
                           , A => n645, ZN => n1657);
   U322 : AOI222_X1 port map( A1 => n28, A2 => n2156, B1 => n2150, B2 => n646, 
                           C1 => n92, C2 => n2144, ZN => n645);
   U323 : OAI221_X1 port map( B1 => n2167, B2 => n647, C1 => n1912, C2 => n2162
                           , A => n648, ZN => n1656);
   U324 : AOI222_X1 port map( A1 => n27, A2 => n2156, B1 => n2151, B2 => n649, 
                           C1 => n91, C2 => n2144, ZN => n648);
   U325 : OAI221_X1 port map( B1 => n2167, B2 => n650, C1 => n1911, C2 => n2162
                           , A => n651, ZN => n1655);
   U326 : AOI222_X1 port map( A1 => n26, A2 => n2156, B1 => n2151, B2 => n652, 
                           C1 => n90, C2 => n2144, ZN => n651);
   U327 : OAI221_X1 port map( B1 => n2167, B2 => n653, C1 => n1910, C2 => n2162
                           , A => n654, ZN => n1654);
   U328 : AOI222_X1 port map( A1 => n25, A2 => n2156, B1 => n2151, B2 => n655, 
                           C1 => n89, C2 => n2144, ZN => n654);
   U329 : OAI221_X1 port map( B1 => n2166, B2 => n656, C1 => n1909, C2 => n2162
                           , A => n657, ZN => n1653);
   U330 : AOI222_X1 port map( A1 => n24, A2 => n2156, B1 => n2151, B2 => n658, 
                           C1 => n88, C2 => n2143, ZN => n657);
   U331 : OAI221_X1 port map( B1 => n2166, B2 => n659, C1 => n1908, C2 => n2162
                           , A => n660, ZN => n1652);
   U332 : AOI222_X1 port map( A1 => n23, A2 => n2156, B1 => n2151, B2 => n661, 
                           C1 => n87, C2 => n2143, ZN => n660);
   U333 : OAI221_X1 port map( B1 => n2166, B2 => n662, C1 => n1907, C2 => n2162
                           , A => n663, ZN => n1651);
   U334 : AOI222_X1 port map( A1 => n22, A2 => n2156, B1 => n2151, B2 => n664, 
                           C1 => n86, C2 => n2143, ZN => n663);
   U335 : OAI221_X1 port map( B1 => n2166, B2 => n665, C1 => n1906, C2 => n2162
                           , A => n666, ZN => n1650);
   U336 : AOI222_X1 port map( A1 => n21, A2 => n2156, B1 => n2151, B2 => n667, 
                           C1 => n85, C2 => n2143, ZN => n666);
   U337 : OAI221_X1 port map( B1 => n2166, B2 => n668, C1 => n1905, C2 => n2162
                           , A => n669, ZN => n1649);
   U338 : AOI222_X1 port map( A1 => n20, A2 => n2156, B1 => n2151, B2 => n670, 
                           C1 => n84, C2 => n2143, ZN => n669);
   U339 : OAI221_X1 port map( B1 => n2166, B2 => n671, C1 => n1904, C2 => n2162
                           , A => n672, ZN => n1648);
   U340 : AOI222_X1 port map( A1 => n19, A2 => n2156, B1 => n2151, B2 => n673, 
                           C1 => n83, C2 => n2143, ZN => n672);
   U341 : OAI221_X1 port map( B1 => n2166, B2 => n674, C1 => n1903, C2 => n2162
                           , A => n675, ZN => n1647);
   U342 : AOI222_X1 port map( A1 => n18, A2 => n2156, B1 => n2151, B2 => n676, 
                           C1 => n82, C2 => n2143, ZN => n675);
   U343 : OAI221_X1 port map( B1 => n2166, B2 => n677, C1 => n1902, C2 => n2162
                           , A => n678, ZN => n1646);
   U344 : AOI222_X1 port map( A1 => n17, A2 => n2156, B1 => n2151, B2 => n679, 
                           C1 => n81, C2 => n2143, ZN => n678);
   U345 : OAI221_X1 port map( B1 => n2166, B2 => n680, C1 => n1901, C2 => n2163
                           , A => n681, ZN => n1645);
   U346 : AOI222_X1 port map( A1 => n16, A2 => n2157, B1 => n2151, B2 => n682, 
                           C1 => n80, C2 => n2143, ZN => n681);
   U347 : OAI221_X1 port map( B1 => n2166, B2 => n683, C1 => n1900, C2 => n2163
                           , A => n684, ZN => n1644);
   U348 : AOI222_X1 port map( A1 => n15, A2 => n2157, B1 => n2151, B2 => n685, 
                           C1 => n79, C2 => n2143, ZN => n684);
   U349 : OAI221_X1 port map( B1 => n2166, B2 => n686, C1 => n1899, C2 => n2163
                           , A => n687, ZN => n1643);
   U350 : AOI222_X1 port map( A1 => n14, A2 => n2157, B1 => n2152, B2 => n688, 
                           C1 => n78, C2 => n2143, ZN => n687);
   U351 : OAI221_X1 port map( B1 => n2166, B2 => n689, C1 => n1898, C2 => n2163
                           , A => n690, ZN => n1642);
   U352 : AOI222_X1 port map( A1 => n13, A2 => n2157, B1 => n2152, B2 => n691, 
                           C1 => n77, C2 => n2143, ZN => n690);
   U353 : OAI221_X1 port map( B1 => n2165, B2 => n692, C1 => n1897, C2 => n2163
                           , A => n693, ZN => n1641);
   U354 : AOI222_X1 port map( A1 => n2158, A2 => n694, B1 => n2152, B2 => n695,
                           C1 => n76, C2 => n2142, ZN => n693);
   U355 : OAI221_X1 port map( B1 => n2165, B2 => n696, C1 => n1896, C2 => n2163
                           , A => n697, ZN => n1640);
   U356 : AOI222_X1 port map( A1 => n2158, A2 => n698, B1 => n2152, B2 => n699,
                           C1 => n75, C2 => n2142, ZN => n697);
   U357 : OAI221_X1 port map( B1 => n2165, B2 => n700, C1 => n1895, C2 => n2163
                           , A => n701, ZN => n1639);
   U358 : AOI222_X1 port map( A1 => n2158, A2 => n702, B1 => n2152, B2 => n703,
                           C1 => n74, C2 => n2142, ZN => n701);
   U359 : OAI221_X1 port map( B1 => n2165, B2 => n704, C1 => n1894, C2 => n2163
                           , A => n705, ZN => n1638);
   U360 : AOI222_X1 port map( A1 => n9, A2 => n2157, B1 => n2152, B2 => n706, 
                           C1 => n73, C2 => n2142, ZN => n705);
   U361 : OAI221_X1 port map( B1 => n2165, B2 => n707, C1 => n1893, C2 => n2163
                           , A => n708, ZN => n1637);
   U362 : AOI222_X1 port map( A1 => n8, A2 => n2157, B1 => n2152, B2 => n709, 
                           C1 => n72, C2 => n2142, ZN => n708);
   U363 : OAI221_X1 port map( B1 => n2165, B2 => n710, C1 => n1892, C2 => n2163
                           , A => n711, ZN => n1636);
   U364 : AOI222_X1 port map( A1 => n7, A2 => n2157, B1 => n2152, B2 => n712, 
                           C1 => n71, C2 => n2142, ZN => n711);
   U365 : OAI221_X1 port map( B1 => n2165, B2 => n713, C1 => n1891, C2 => n2163
                           , A => n714, ZN => n1635);
   U366 : AOI222_X1 port map( A1 => n6, A2 => n2157, B1 => n2152, B2 => n715, 
                           C1 => n70, C2 => n2142, ZN => n714);
   U367 : OAI221_X1 port map( B1 => n2165, B2 => n719, C1 => n1889, C2 => n2163
                           , A => n720, ZN => n1633);
   U368 : AOI222_X1 port map( A1 => n4, A2 => n2157, B1 => n2152, B2 => n721, 
                           C1 => n68, C2 => n2142, ZN => n720);
   U369 : OAI221_X1 port map( B1 => n522, B2 => n2141, C1 => n1885, C2 => n2130
                           , A => n737, ZN => n1629);
   U370 : AOI222_X1 port map( A1 => n2129, A2 => n64, B1 => n2123, B2 => n192, 
                           C1 => n2117, C2 => n528, ZN => n737);
   U371 : OAI221_X1 port map( B1 => n529, B2 => n2141, C1 => n1884, C2 => n2130
                           , A => n744, ZN => n1627);
   U372 : AOI222_X1 port map( A1 => n2129, A2 => n63, B1 => n2123, B2 => n191, 
                           C1 => n2117, C2 => n531, ZN => n744);
   U373 : OAI221_X1 port map( B1 => n532, B2 => n2141, C1 => n1883, C2 => n2130
                           , A => n746, ZN => n1625);
   U374 : AOI222_X1 port map( A1 => n2129, A2 => n62, B1 => n2123, B2 => n190, 
                           C1 => n2117, C2 => n534, ZN => n746);
   U375 : OAI221_X1 port map( B1 => n535, B2 => n2141, C1 => n1882, C2 => n2130
                           , A => n748, ZN => n1623);
   U376 : AOI222_X1 port map( A1 => n2129, A2 => n61, B1 => n2123, B2 => n189, 
                           C1 => n2117, C2 => n537, ZN => n748);
   U377 : OAI221_X1 port map( B1 => n583, B2 => n2139, C1 => n1866, C2 => n2131
                           , A => n780, ZN => n1591);
   U378 : AOI222_X1 port map( A1 => n2127, A2 => n45, B1 => n2121, B2 => n585, 
                           C1 => n2115, C2 => n586, ZN => n780);
   U379 : OAI221_X1 port map( B1 => n587, B2 => n2139, C1 => n1865, C2 => n2131
                           , A => n782, ZN => n1589);
   U380 : AOI222_X1 port map( A1 => n2127, A2 => n44, B1 => n2121, B2 => n589, 
                           C1 => n2115, C2 => n590, ZN => n782);
   U381 : OAI221_X1 port map( B1 => n591, B2 => n2139, C1 => n1864, C2 => n2131
                           , A => n784, ZN => n1587);
   U382 : AOI222_X1 port map( A1 => n2127, A2 => n43, B1 => n2121, B2 => n593, 
                           C1 => n2115, C2 => n594, ZN => n784);
   U383 : OAI221_X1 port map( B1 => n595, B2 => n2139, C1 => n1863, C2 => n2131
                           , A => n786, ZN => n1585);
   U384 : AOI222_X1 port map( A1 => n2127, A2 => n42, B1 => n2121, B2 => n597, 
                           C1 => n2115, C2 => n598, ZN => n786);
   U385 : OAI221_X1 port map( B1 => n599, B2 => n2139, C1 => n1862, C2 => n2131
                           , A => n788, ZN => n1583);
   U386 : AOI222_X1 port map( A1 => n2127, A2 => n41, B1 => n2121, B2 => n601, 
                           C1 => n2115, C2 => n602, ZN => n788);
   U387 : OAI221_X1 port map( B1 => n603, B2 => n2139, C1 => n1861, C2 => n2131
                           , A => n790, ZN => n1581);
   U388 : AOI222_X1 port map( A1 => n2127, A2 => n40, B1 => n2121, B2 => n605, 
                           C1 => n2115, C2 => n606, ZN => n790);
   U389 : OAI221_X1 port map( B1 => n607, B2 => n2139, C1 => n1860, C2 => n2132
                           , A => n792, ZN => n1579);
   U390 : AOI222_X1 port map( A1 => n2127, A2 => n39, B1 => n2121, B2 => n609, 
                           C1 => n2115, C2 => n610, ZN => n792);
   U391 : OAI221_X1 port map( B1 => n611, B2 => n2139, C1 => n1859, C2 => n2132
                           , A => n794, ZN => n1577);
   U392 : AOI222_X1 port map( A1 => n2127, A2 => n38, B1 => n2121, B2 => n613, 
                           C1 => n2115, C2 => n614, ZN => n794);
   U393 : OAI221_X1 port map( B1 => n615, B2 => n2139, C1 => n1858, C2 => n2132
                           , A => n796, ZN => n1575);
   U394 : AOI222_X1 port map( A1 => n2127, A2 => n37, B1 => n2121, B2 => n617, 
                           C1 => n2115, C2 => n618, ZN => n796);
   U395 : OAI221_X1 port map( B1 => n619, B2 => n2138, C1 => n1857, C2 => n2132
                           , A => n798, ZN => n1573);
   U396 : AOI222_X1 port map( A1 => n2126, A2 => n36, B1 => n2120, B2 => n621, 
                           C1 => n2114, C2 => n622, ZN => n798);
   U397 : OAI221_X1 port map( B1 => n2169, B2 => n538, C1 => n1945, C2 => n2159
                           , A => n539, ZN => n1689);
   U398 : AOI222_X1 port map( A1 => n60, A2 => n2153, B1 => n188, B2 => n2148, 
                           C1 => n2146, C2 => n540, ZN => n539);
   U399 : OAI221_X1 port map( B1 => n2169, B2 => n541, C1 => n1944, C2 => n2159
                           , A => n542, ZN => n1688);
   U400 : AOI222_X1 port map( A1 => n59, A2 => n2153, B1 => n187, B2 => n2148, 
                           C1 => n2146, C2 => n543, ZN => n542);
   U401 : OAI221_X1 port map( B1 => n2169, B2 => n544, C1 => n1943, C2 => n2159
                           , A => n545, ZN => n1687);
   U402 : AOI222_X1 port map( A1 => n58, A2 => n2153, B1 => n186, B2 => n2148, 
                           C1 => n2146, C2 => n546, ZN => n545);
   U403 : OAI221_X1 port map( B1 => n2169, B2 => n547, C1 => n1942, C2 => n2159
                           , A => n548, ZN => n1686);
   U404 : AOI222_X1 port map( A1 => n57, A2 => n2153, B1 => n185, B2 => n2148, 
                           C1 => n2146, C2 => n549, ZN => n548);
   U405 : OAI221_X1 port map( B1 => n2169, B2 => n550, C1 => n1941, C2 => n2159
                           , A => n551, ZN => n1685);
   U406 : AOI222_X1 port map( A1 => n56, A2 => n2153, B1 => n184, B2 => n2148, 
                           C1 => n2146, C2 => n552, ZN => n551);
   U407 : OAI221_X1 port map( B1 => n2169, B2 => n553, C1 => n1940, C2 => n2159
                           , A => n554, ZN => n1684);
   U408 : AOI222_X1 port map( A1 => n55, A2 => n2153, B1 => n183, B2 => n2148, 
                           C1 => n2146, C2 => n555, ZN => n554);
   U409 : OAI221_X1 port map( B1 => n2169, B2 => n556, C1 => n1939, C2 => n2159
                           , A => n557, ZN => n1683);
   U410 : AOI222_X1 port map( A1 => n54, A2 => n2153, B1 => n182, B2 => n2148, 
                           C1 => n2146, C2 => n558, ZN => n557);
   U411 : OAI221_X1 port map( B1 => n2169, B2 => n559, C1 => n1938, C2 => n2159
                           , A => n560, ZN => n1682);
   U412 : AOI222_X1 port map( A1 => n53, A2 => n2153, B1 => n181, B2 => n2148, 
                           C1 => n2146, C2 => n561, ZN => n560);
   U413 : OAI221_X1 port map( B1 => n2168, B2 => n583, C1 => n1930, C2 => n2160
                           , A => n584, ZN => n1674);
   U414 : AOI222_X1 port map( A1 => n45, A2 => n2154, B1 => n2149, B2 => n585, 
                           C1 => n2145, C2 => n586, ZN => n584);
   U415 : OAI221_X1 port map( B1 => n2168, B2 => n587, C1 => n1929, C2 => n2160
                           , A => n588, ZN => n1673);
   U416 : AOI222_X1 port map( A1 => n44, A2 => n2154, B1 => n2149, B2 => n589, 
                           C1 => n2145, C2 => n590, ZN => n588);
   U417 : OAI221_X1 port map( B1 => n2168, B2 => n591, C1 => n1928, C2 => n2160
                           , A => n592, ZN => n1672);
   U418 : AOI222_X1 port map( A1 => n43, A2 => n2154, B1 => n2149, B2 => n593, 
                           C1 => n2145, C2 => n594, ZN => n592);
   U419 : OAI221_X1 port map( B1 => n2168, B2 => n595, C1 => n1927, C2 => n2160
                           , A => n596, ZN => n1671);
   U420 : AOI222_X1 port map( A1 => n42, A2 => n2154, B1 => n2149, B2 => n597, 
                           C1 => n2145, C2 => n598, ZN => n596);
   U421 : OAI221_X1 port map( B1 => n2168, B2 => n599, C1 => n1926, C2 => n2160
                           , A => n600, ZN => n1670);
   U422 : AOI222_X1 port map( A1 => n41, A2 => n2154, B1 => n2149, B2 => n601, 
                           C1 => n2145, C2 => n602, ZN => n600);
   U423 : OAI221_X1 port map( B1 => n2168, B2 => n603, C1 => n1925, C2 => n2160
                           , A => n604, ZN => n1669);
   U424 : AOI222_X1 port map( A1 => n40, A2 => n2154, B1 => n2150, B2 => n605, 
                           C1 => n2145, C2 => n606, ZN => n604);
   U425 : OAI221_X1 port map( B1 => n2168, B2 => n607, C1 => n1924, C2 => n2161
                           , A => n608, ZN => n1668);
   U426 : AOI222_X1 port map( A1 => n39, A2 => n2155, B1 => n2150, B2 => n609, 
                           C1 => n2145, C2 => n610, ZN => n608);
   U427 : OAI221_X1 port map( B1 => n2168, B2 => n611, C1 => n1923, C2 => n2161
                           , A => n612, ZN => n1667);
   U428 : AOI222_X1 port map( A1 => n38, A2 => n2155, B1 => n2150, B2 => n613, 
                           C1 => n2145, C2 => n614, ZN => n612);
   U429 : OAI221_X1 port map( B1 => n2168, B2 => n615, C1 => n1922, C2 => n2161
                           , A => n616, ZN => n1666);
   U430 : AOI222_X1 port map( A1 => n37, A2 => n2155, B1 => n2150, B2 => n617, 
                           C1 => n2145, C2 => n618, ZN => n616);
   U431 : OAI22_X1 port map( A1 => n1950, A2 => n2099, B1 => n743, B2 => n2093,
                           ZN => n1501);
   U432 : OAI22_X1 port map( A1 => n1951, A2 => n2099, B1 => n745, B2 => n2093,
                           ZN => n1500);
   U433 : OAI22_X1 port map( A1 => n1952, A2 => n2099, B1 => n747, B2 => n2093,
                           ZN => n1499);
   U434 : OAI22_X1 port map( A1 => n1953, A2 => n2099, B1 => n749, B2 => n2093,
                           ZN => n1498);
   U435 : OAI22_X1 port map( A1 => n1821, A2 => n2087, B1 => n743, B2 => n2081,
                           ZN => n1437);
   U436 : OAI22_X1 port map( A1 => n1820, A2 => n2087, B1 => n745, B2 => n2081,
                           ZN => n1436);
   U437 : OAI22_X1 port map( A1 => n1819, A2 => n2087, B1 => n747, B2 => n2081,
                           ZN => n1435);
   U438 : OAI22_X1 port map( A1 => n1818, A2 => n2087, B1 => n749, B2 => n2081,
                           ZN => n1434);
   U439 : OAI22_X1 port map( A1 => n2010, A2 => n2075, B1 => n743, B2 => n2069,
                           ZN => n1373);
   U440 : OAI22_X1 port map( A1 => n2011, A2 => n2075, B1 => n745, B2 => n2069,
                           ZN => n1372);
   U441 : OAI22_X1 port map( A1 => n2012, A2 => n2075, B1 => n747, B2 => n2069,
                           ZN => n1371);
   U442 : OAI22_X1 port map( A1 => n2013, A2 => n2075, B1 => n749, B2 => n2069,
                           ZN => n1370);
   U443 : OAI22_X1 port map( A1 => n1954, A2 => n2099, B1 => n751, B2 => n2092,
                           ZN => n1497);
   U444 : OAI22_X1 port map( A1 => n1955, A2 => n2098, B1 => n753, B2 => n2092,
                           ZN => n1496);
   U445 : OAI22_X1 port map( A1 => n1956, A2 => n2098, B1 => n755, B2 => n2092,
                           ZN => n1495);
   U446 : OAI22_X1 port map( A1 => n1957, A2 => n2098, B1 => n757, B2 => n2092,
                           ZN => n1494);
   U447 : OAI22_X1 port map( A1 => n1958, A2 => n2098, B1 => n759, B2 => n2092,
                           ZN => n1493);
   U448 : OAI22_X1 port map( A1 => n1959, A2 => n2098, B1 => n761, B2 => n2092,
                           ZN => n1492);
   U449 : OAI22_X1 port map( A1 => n1960, A2 => n2098, B1 => n763, B2 => n2092,
                           ZN => n1491);
   U450 : OAI22_X1 port map( A1 => n1961, A2 => n2098, B1 => n765, B2 => n2092,
                           ZN => n1490);
   U451 : OAI22_X1 port map( A1 => n1962, A2 => n2098, B1 => n767, B2 => n2092,
                           ZN => n1489);
   U452 : OAI22_X1 port map( A1 => n1963, A2 => n2098, B1 => n769, B2 => n2092,
                           ZN => n1488);
   U453 : OAI22_X1 port map( A1 => n1964, A2 => n2098, B1 => n771, B2 => n2092,
                           ZN => n1487);
   U454 : OAI22_X1 port map( A1 => n1965, A2 => n2098, B1 => n773, B2 => n2092,
                           ZN => n1486);
   U455 : OAI22_X1 port map( A1 => n1966, A2 => n2098, B1 => n775, B2 => n2091,
                           ZN => n1485);
   U456 : OAI22_X1 port map( A1 => n1967, A2 => n2097, B1 => n777, B2 => n2091,
                           ZN => n1484);
   U457 : OAI22_X1 port map( A1 => n1968, A2 => n2097, B1 => n779, B2 => n2091,
                           ZN => n1483);
   U458 : OAI22_X1 port map( A1 => n1969, A2 => n2097, B1 => n781, B2 => n2091,
                           ZN => n1482);
   U459 : OAI22_X1 port map( A1 => n1970, A2 => n2097, B1 => n783, B2 => n2091,
                           ZN => n1481);
   U460 : OAI22_X1 port map( A1 => n1971, A2 => n2097, B1 => n785, B2 => n2091,
                           ZN => n1480);
   U461 : OAI22_X1 port map( A1 => n1972, A2 => n2097, B1 => n787, B2 => n2091,
                           ZN => n1479);
   U462 : OAI22_X1 port map( A1 => n1973, A2 => n2097, B1 => n789, B2 => n2091,
                           ZN => n1478);
   U463 : OAI22_X1 port map( A1 => n1974, A2 => n2097, B1 => n791, B2 => n2091,
                           ZN => n1477);
   U464 : OAI22_X1 port map( A1 => n1975, A2 => n2097, B1 => n793, B2 => n2091,
                           ZN => n1476);
   U465 : OAI22_X1 port map( A1 => n1976, A2 => n2097, B1 => n795, B2 => n2091,
                           ZN => n1475);
   U466 : OAI22_X1 port map( A1 => n1977, A2 => n2097, B1 => n797, B2 => n2091,
                           ZN => n1474);
   U467 : OAI22_X1 port map( A1 => n1978, A2 => n2097, B1 => n799, B2 => n2090,
                           ZN => n1473);
   U468 : OAI22_X1 port map( A1 => n1979, A2 => n2096, B1 => n801, B2 => n2090,
                           ZN => n1472);
   U469 : OAI22_X1 port map( A1 => n1980, A2 => n2096, B1 => n803, B2 => n2090,
                           ZN => n1471);
   U470 : OAI22_X1 port map( A1 => n1981, A2 => n2096, B1 => n805, B2 => n2090,
                           ZN => n1470);
   U471 : OAI22_X1 port map( A1 => n1982, A2 => n2096, B1 => n807, B2 => n2090,
                           ZN => n1469);
   U472 : OAI22_X1 port map( A1 => n1983, A2 => n2096, B1 => n809, B2 => n2090,
                           ZN => n1468);
   U473 : OAI22_X1 port map( A1 => n1984, A2 => n2096, B1 => n811, B2 => n2090,
                           ZN => n1467);
   U474 : OAI22_X1 port map( A1 => n1985, A2 => n2096, B1 => n813, B2 => n2090,
                           ZN => n1466);
   U475 : OAI22_X1 port map( A1 => n1986, A2 => n2096, B1 => n815, B2 => n2090,
                           ZN => n1465);
   U476 : OAI22_X1 port map( A1 => n1987, A2 => n2096, B1 => n817, B2 => n2090,
                           ZN => n1464);
   U477 : OAI22_X1 port map( A1 => n1988, A2 => n2096, B1 => n819, B2 => n2090,
                           ZN => n1463);
   U478 : OAI22_X1 port map( A1 => n1989, A2 => n2096, B1 => n821, B2 => n2090,
                           ZN => n1462);
   U479 : OAI22_X1 port map( A1 => n1990, A2 => n2096, B1 => n823, B2 => n2089,
                           ZN => n1461);
   U480 : OAI22_X1 port map( A1 => n1991, A2 => n2095, B1 => n825, B2 => n2089,
                           ZN => n1460);
   U481 : OAI22_X1 port map( A1 => n1992, A2 => n2095, B1 => n827, B2 => n2089,
                           ZN => n1459);
   U482 : OAI22_X1 port map( A1 => n1993, A2 => n2095, B1 => n829, B2 => n2089,
                           ZN => n1458);
   U483 : OAI22_X1 port map( A1 => n1994, A2 => n2095, B1 => n831, B2 => n2089,
                           ZN => n1457);
   U484 : OAI22_X1 port map( A1 => n1995, A2 => n2095, B1 => n833, B2 => n2089,
                           ZN => n1456);
   U485 : OAI22_X1 port map( A1 => n1996, A2 => n2095, B1 => n835, B2 => n2089,
                           ZN => n1455);
   U486 : OAI22_X1 port map( A1 => n1997, A2 => n2095, B1 => n837, B2 => n2089,
                           ZN => n1454);
   U487 : OAI22_X1 port map( A1 => n1998, A2 => n2095, B1 => n839, B2 => n2089,
                           ZN => n1453);
   U488 : OAI22_X1 port map( A1 => n1999, A2 => n2095, B1 => n841, B2 => n2089,
                           ZN => n1452);
   U489 : OAI22_X1 port map( A1 => n2000, A2 => n2095, B1 => n843, B2 => n2089,
                           ZN => n1451);
   U490 : OAI22_X1 port map( A1 => n2001, A2 => n2095, B1 => n845, B2 => n2089,
                           ZN => n1450);
   U491 : OAI22_X1 port map( A1 => n1204, A2 => n2095, B1 => n847, B2 => n2088,
                           ZN => n1449);
   U492 : OAI22_X1 port map( A1 => n1202, A2 => n2094, B1 => n849, B2 => n2088,
                           ZN => n1448);
   U493 : OAI22_X1 port map( A1 => n1200, A2 => n2094, B1 => n851, B2 => n2088,
                           ZN => n1447);
   U494 : OAI22_X1 port map( A1 => n2002, A2 => n2094, B1 => n853, B2 => n2088,
                           ZN => n1446);
   U495 : OAI22_X1 port map( A1 => n2003, A2 => n2094, B1 => n855, B2 => n2088,
                           ZN => n1445);
   U496 : OAI22_X1 port map( A1 => n2004, A2 => n2094, B1 => n857, B2 => n2088,
                           ZN => n1444);
   U497 : OAI22_X1 port map( A1 => n2005, A2 => n2094, B1 => n859, B2 => n2088,
                           ZN => n1443);
   U498 : OAI22_X1 port map( A1 => n2006, A2 => n2094, B1 => n861, B2 => n2088,
                           ZN => n1442);
   U499 : OAI22_X1 port map( A1 => n2007, A2 => n2094, B1 => n863, B2 => n2088,
                           ZN => n1441);
   U500 : OAI22_X1 port map( A1 => n2008, A2 => n2094, B1 => n865, B2 => n2088,
                           ZN => n1440);
   U501 : OAI22_X1 port map( A1 => n2009, A2 => n2094, B1 => n867, B2 => n2088,
                           ZN => n1439);
   U502 : OAI22_X1 port map( A1 => n415, A2 => n2094, B1 => n871, B2 => n2088, 
                           ZN => n1438);
   U503 : OAI22_X1 port map( A1 => n1817, A2 => n2087, B1 => n751, B2 => n2080,
                           ZN => n1433);
   U504 : OAI22_X1 port map( A1 => n1816, A2 => n2086, B1 => n753, B2 => n2080,
                           ZN => n1432);
   U505 : OAI22_X1 port map( A1 => n1815, A2 => n2086, B1 => n755, B2 => n2080,
                           ZN => n1431);
   U506 : OAI22_X1 port map( A1 => n1814, A2 => n2086, B1 => n757, B2 => n2080,
                           ZN => n1430);
   U507 : OAI22_X1 port map( A1 => n1813, A2 => n2086, B1 => n759, B2 => n2080,
                           ZN => n1429);
   U508 : OAI22_X1 port map( A1 => n1812, A2 => n2086, B1 => n761, B2 => n2080,
                           ZN => n1428);
   U509 : OAI22_X1 port map( A1 => n1811, A2 => n2086, B1 => n763, B2 => n2080,
                           ZN => n1427);
   U510 : OAI22_X1 port map( A1 => n1810, A2 => n2086, B1 => n765, B2 => n2080,
                           ZN => n1426);
   U511 : OAI22_X1 port map( A1 => n1809, A2 => n2086, B1 => n767, B2 => n2080,
                           ZN => n1425);
   U512 : OAI22_X1 port map( A1 => n1808, A2 => n2086, B1 => n769, B2 => n2080,
                           ZN => n1424);
   U513 : OAI22_X1 port map( A1 => n1807, A2 => n2086, B1 => n771, B2 => n2080,
                           ZN => n1423);
   U514 : OAI22_X1 port map( A1 => n1806, A2 => n2086, B1 => n773, B2 => n2080,
                           ZN => n1422);
   U515 : OAI22_X1 port map( A1 => n1805, A2 => n2086, B1 => n775, B2 => n2079,
                           ZN => n1421);
   U516 : OAI22_X1 port map( A1 => n1804, A2 => n2085, B1 => n777, B2 => n2079,
                           ZN => n1420);
   U517 : OAI22_X1 port map( A1 => n1803, A2 => n2085, B1 => n779, B2 => n2079,
                           ZN => n1419);
   U518 : OAI22_X1 port map( A1 => n1802, A2 => n2085, B1 => n781, B2 => n2079,
                           ZN => n1418);
   U519 : OAI22_X1 port map( A1 => n1801, A2 => n2085, B1 => n783, B2 => n2079,
                           ZN => n1417);
   U520 : OAI22_X1 port map( A1 => n1800, A2 => n2085, B1 => n785, B2 => n2079,
                           ZN => n1416);
   U521 : OAI22_X1 port map( A1 => n1799, A2 => n2085, B1 => n787, B2 => n2079,
                           ZN => n1415);
   U522 : OAI22_X1 port map( A1 => n1798, A2 => n2085, B1 => n789, B2 => n2079,
                           ZN => n1414);
   U523 : OAI22_X1 port map( A1 => n1797, A2 => n2085, B1 => n791, B2 => n2079,
                           ZN => n1413);
   U524 : OAI22_X1 port map( A1 => n1796, A2 => n2085, B1 => n793, B2 => n2079,
                           ZN => n1412);
   U525 : OAI22_X1 port map( A1 => n1795, A2 => n2085, B1 => n795, B2 => n2079,
                           ZN => n1411);
   U526 : OAI22_X1 port map( A1 => n1794, A2 => n2085, B1 => n797, B2 => n2079,
                           ZN => n1410);
   U527 : OAI22_X1 port map( A1 => n1793, A2 => n2085, B1 => n799, B2 => n2078,
                           ZN => n1409);
   U528 : OAI22_X1 port map( A1 => n2029, A2 => n2084, B1 => n801, B2 => n2078,
                           ZN => n1408);
   U529 : OAI22_X1 port map( A1 => n2030, A2 => n2084, B1 => n803, B2 => n2078,
                           ZN => n1407);
   U530 : OAI22_X1 port map( A1 => n2031, A2 => n2084, B1 => n805, B2 => n2078,
                           ZN => n1406);
   U531 : OAI22_X1 port map( A1 => n2032, A2 => n2084, B1 => n807, B2 => n2078,
                           ZN => n1405);
   U532 : OAI22_X1 port map( A1 => n2033, A2 => n2084, B1 => n809, B2 => n2078,
                           ZN => n1404);
   U533 : OAI22_X1 port map( A1 => n2034, A2 => n2084, B1 => n811, B2 => n2078,
                           ZN => n1403);
   U534 : OAI22_X1 port map( A1 => n2035, A2 => n2084, B1 => n813, B2 => n2078,
                           ZN => n1402);
   U535 : OAI22_X1 port map( A1 => n2036, A2 => n2084, B1 => n815, B2 => n2078,
                           ZN => n1401);
   U536 : OAI22_X1 port map( A1 => n2037, A2 => n2084, B1 => n817, B2 => n2078,
                           ZN => n1400);
   U537 : OAI22_X1 port map( A1 => n2038, A2 => n2084, B1 => n819, B2 => n2078,
                           ZN => n1399);
   U538 : OAI22_X1 port map( A1 => n2039, A2 => n2084, B1 => n821, B2 => n2078,
                           ZN => n1398);
   U539 : OAI22_X1 port map( A1 => n2040, A2 => n2084, B1 => n823, B2 => n2077,
                           ZN => n1397);
   U540 : OAI22_X1 port map( A1 => n2041, A2 => n2083, B1 => n825, B2 => n2077,
                           ZN => n1396);
   U541 : OAI22_X1 port map( A1 => n2042, A2 => n2083, B1 => n827, B2 => n2077,
                           ZN => n1395);
   U542 : OAI22_X1 port map( A1 => n2043, A2 => n2083, B1 => n829, B2 => n2077,
                           ZN => n1394);
   U543 : OAI22_X1 port map( A1 => n2044, A2 => n2083, B1 => n831, B2 => n2077,
                           ZN => n1393);
   U544 : OAI22_X1 port map( A1 => n2045, A2 => n2083, B1 => n833, B2 => n2077,
                           ZN => n1392);
   U545 : OAI22_X1 port map( A1 => n2046, A2 => n2083, B1 => n835, B2 => n2077,
                           ZN => n1391);
   U546 : OAI22_X1 port map( A1 => n2047, A2 => n2083, B1 => n837, B2 => n2077,
                           ZN => n1390);
   U547 : OAI22_X1 port map( A1 => n2048, A2 => n2083, B1 => n839, B2 => n2077,
                           ZN => n1389);
   U548 : OAI22_X1 port map( A1 => n2049, A2 => n2083, B1 => n841, B2 => n2077,
                           ZN => n1388);
   U549 : OAI22_X1 port map( A1 => n2050, A2 => n2083, B1 => n843, B2 => n2077,
                           ZN => n1387);
   U550 : OAI22_X1 port map( A1 => n2051, A2 => n2083, B1 => n845, B2 => n2077,
                           ZN => n1386);
   U551 : OAI22_X1 port map( A1 => n2052, A2 => n2083, B1 => n847, B2 => n2076,
                           ZN => n1385);
   U552 : OAI22_X1 port map( A1 => n2053, A2 => n2082, B1 => n849, B2 => n2076,
                           ZN => n1384);
   U553 : OAI22_X1 port map( A1 => n2054, A2 => n2082, B1 => n851, B2 => n2076,
                           ZN => n1383);
   U554 : OAI22_X1 port map( A1 => n2055, A2 => n2082, B1 => n853, B2 => n2076,
                           ZN => n1382);
   U555 : OAI22_X1 port map( A1 => n2056, A2 => n2082, B1 => n855, B2 => n2076,
                           ZN => n1381);
   U556 : OAI22_X1 port map( A1 => n2057, A2 => n2082, B1 => n857, B2 => n2076,
                           ZN => n1380);
   U557 : OAI22_X1 port map( A1 => n2058, A2 => n2082, B1 => n859, B2 => n2076,
                           ZN => n1379);
   U558 : OAI22_X1 port map( A1 => n2059, A2 => n2082, B1 => n861, B2 => n2076,
                           ZN => n1378);
   U559 : OAI22_X1 port map( A1 => n2060, A2 => n2082, B1 => n863, B2 => n2076,
                           ZN => n1377);
   U560 : OAI22_X1 port map( A1 => n2061, A2 => n2082, B1 => n865, B2 => n2076,
                           ZN => n1376);
   U561 : OAI22_X1 port map( A1 => n2062, A2 => n2082, B1 => n867, B2 => n2076,
                           ZN => n1375);
   U562 : OAI22_X1 port map( A1 => n2063, A2 => n2082, B1 => n871, B2 => n2076,
                           ZN => n1374);
   U563 : OAI22_X1 port map( A1 => n2014, A2 => n2075, B1 => n751, B2 => n2068,
                           ZN => n1369);
   U564 : OAI22_X1 port map( A1 => n2015, A2 => n2074, B1 => n753, B2 => n2068,
                           ZN => n1368);
   U565 : OAI22_X1 port map( A1 => n2016, A2 => n2074, B1 => n755, B2 => n2068,
                           ZN => n1367);
   U566 : OAI22_X1 port map( A1 => n2017, A2 => n2074, B1 => n757, B2 => n2068,
                           ZN => n1366);
   U567 : OAI22_X1 port map( A1 => n2018, A2 => n2074, B1 => n759, B2 => n2068,
                           ZN => n1365);
   U568 : OAI22_X1 port map( A1 => n2019, A2 => n2074, B1 => n761, B2 => n2068,
                           ZN => n1364);
   U569 : OAI22_X1 port map( A1 => n2020, A2 => n2074, B1 => n763, B2 => n2068,
                           ZN => n1363);
   U570 : OAI22_X1 port map( A1 => n2021, A2 => n2074, B1 => n765, B2 => n2068,
                           ZN => n1362);
   U571 : OAI22_X1 port map( A1 => n2022, A2 => n2074, B1 => n767, B2 => n2068,
                           ZN => n1361);
   U572 : OAI22_X1 port map( A1 => n2023, A2 => n2074, B1 => n769, B2 => n2068,
                           ZN => n1360);
   U573 : OAI22_X1 port map( A1 => n2024, A2 => n2074, B1 => n771, B2 => n2068,
                           ZN => n1359);
   U574 : OAI22_X1 port map( A1 => n2025, A2 => n2074, B1 => n773, B2 => n2068,
                           ZN => n1358);
   U575 : OAI22_X1 port map( A1 => n2026, A2 => n2074, B1 => n775, B2 => n2067,
                           ZN => n1357);
   U576 : OAI22_X1 port map( A1 => n2027, A2 => n2073, B1 => n777, B2 => n2067,
                           ZN => n1356);
   U577 : OAI22_X1 port map( A1 => n2028, A2 => n2073, B1 => n779, B2 => n2067,
                           ZN => n1355);
   U578 : OAI22_X1 port map( A1 => n1738, A2 => n2073, B1 => n781, B2 => n2067,
                           ZN => n1354);
   U579 : OAI22_X1 port map( A1 => n1737, A2 => n2073, B1 => n783, B2 => n2067,
                           ZN => n1353);
   U580 : OAI22_X1 port map( A1 => n1736, A2 => n2073, B1 => n785, B2 => n2067,
                           ZN => n1352);
   U581 : OAI22_X1 port map( A1 => n1735, A2 => n2073, B1 => n787, B2 => n2067,
                           ZN => n1351);
   U582 : OAI22_X1 port map( A1 => n1734, A2 => n2073, B1 => n789, B2 => n2067,
                           ZN => n1350);
   U583 : OAI22_X1 port map( A1 => n1733, A2 => n2073, B1 => n791, B2 => n2067,
                           ZN => n1349);
   U584 : OAI22_X1 port map( A1 => n1732, A2 => n2073, B1 => n793, B2 => n2067,
                           ZN => n1348);
   U585 : OAI22_X1 port map( A1 => n1731, A2 => n2073, B1 => n795, B2 => n2067,
                           ZN => n1347);
   U586 : OAI22_X1 port map( A1 => n1730, A2 => n2073, B1 => n797, B2 => n2067,
                           ZN => n1346);
   U587 : OAI22_X1 port map( A1 => n1729, A2 => n2073, B1 => n799, B2 => n2066,
                           ZN => n1345);
   U588 : OAI22_X1 port map( A1 => n1728, A2 => n2072, B1 => n801, B2 => n2066,
                           ZN => n1344);
   U589 : OAI22_X1 port map( A1 => n1727, A2 => n2072, B1 => n803, B2 => n2066,
                           ZN => n1343);
   U590 : OAI22_X1 port map( A1 => n1726, A2 => n2072, B1 => n805, B2 => n2066,
                           ZN => n1342);
   U591 : OAI22_X1 port map( A1 => n1725, A2 => n2072, B1 => n807, B2 => n2066,
                           ZN => n1341);
   U592 : OAI22_X1 port map( A1 => n1724, A2 => n2072, B1 => n809, B2 => n2066,
                           ZN => n1340);
   U593 : OAI22_X1 port map( A1 => n1723, A2 => n2072, B1 => n811, B2 => n2066,
                           ZN => n1339);
   U594 : OAI22_X1 port map( A1 => n1722, A2 => n2072, B1 => n813, B2 => n2066,
                           ZN => n1338);
   U595 : OAI22_X1 port map( A1 => n1721, A2 => n2072, B1 => n815, B2 => n2066,
                           ZN => n1337);
   U596 : OAI22_X1 port map( A1 => n1720, A2 => n2072, B1 => n817, B2 => n2066,
                           ZN => n1336);
   U597 : OAI22_X1 port map( A1 => n1719, A2 => n2072, B1 => n819, B2 => n2066,
                           ZN => n1335);
   U598 : OAI22_X1 port map( A1 => n1718, A2 => n2072, B1 => n821, B2 => n2066,
                           ZN => n1334);
   U599 : OAI22_X1 port map( A1 => n1717, A2 => n2072, B1 => n823, B2 => n2065,
                           ZN => n1333);
   U600 : OAI22_X1 port map( A1 => n1716, A2 => n2071, B1 => n825, B2 => n2065,
                           ZN => n1332);
   U601 : OAI22_X1 port map( A1 => n1715, A2 => n2071, B1 => n827, B2 => n2065,
                           ZN => n1331);
   U602 : OAI22_X1 port map( A1 => n1714, A2 => n2071, B1 => n829, B2 => n2065,
                           ZN => n1330);
   U603 : OAI22_X1 port map( A1 => n1713, A2 => n2071, B1 => n831, B2 => n2065,
                           ZN => n1329);
   U604 : OAI22_X1 port map( A1 => n1712, A2 => n2071, B1 => n833, B2 => n2065,
                           ZN => n1328);
   U605 : OAI22_X1 port map( A1 => n1711, A2 => n2071, B1 => n835, B2 => n2065,
                           ZN => n1327);
   U606 : OAI22_X1 port map( A1 => n1710, A2 => n2071, B1 => n837, B2 => n2065,
                           ZN => n1326);
   U607 : OAI22_X1 port map( A1 => n1709, A2 => n2071, B1 => n839, B2 => n2065,
                           ZN => n1325);
   U608 : OAI22_X1 port map( A1 => n1708, A2 => n2071, B1 => n841, B2 => n2065,
                           ZN => n1324);
   U609 : OAI22_X1 port map( A1 => n1707, A2 => n2071, B1 => n843, B2 => n2065,
                           ZN => n1323);
   U610 : OAI22_X1 port map( A1 => n1706, A2 => n2071, B1 => n845, B2 => n2065,
                           ZN => n1322);
   U611 : OAI22_X1 port map( A1 => n1705, A2 => n2071, B1 => n847, B2 => n2064,
                           ZN => n1321);
   U612 : OAI22_X1 port map( A1 => n1704, A2 => n2070, B1 => n849, B2 => n2064,
                           ZN => n1320);
   U613 : OAI22_X1 port map( A1 => n1703, A2 => n2070, B1 => n851, B2 => n2064,
                           ZN => n1319);
   U614 : OAI22_X1 port map( A1 => n1702, A2 => n2070, B1 => n853, B2 => n2064,
                           ZN => n1318);
   U615 : OAI22_X1 port map( A1 => n1701, A2 => n2070, B1 => n855, B2 => n2064,
                           ZN => n1317);
   U616 : OAI22_X1 port map( A1 => n1700, A2 => n2070, B1 => n857, B2 => n2064,
                           ZN => n1316);
   U617 : OAI22_X1 port map( A1 => n1699, A2 => n2070, B1 => n859, B2 => n2064,
                           ZN => n1315);
   U618 : OAI22_X1 port map( A1 => n1698, A2 => n2070, B1 => n861, B2 => n2064,
                           ZN => n1314);
   U619 : OAI22_X1 port map( A1 => n1697, A2 => n2070, B1 => n863, B2 => n2064,
                           ZN => n1313);
   U620 : OAI22_X1 port map( A1 => n1696, A2 => n2070, B1 => n865, B2 => n2064,
                           ZN => n1312);
   U621 : OAI22_X1 port map( A1 => n1695, A2 => n2070, B1 => n867, B2 => n2064,
                           ZN => n1311);
   U622 : OAI22_X1 port map( A1 => n1694, A2 => n2070, B1 => n871, B2 => n2064,
                           ZN => n1310);
   U623 : INV_X1 port map( A => DATAIN(0), ZN => n743);
   U624 : INV_X1 port map( A => DATAIN(1), ZN => n745);
   U625 : INV_X1 port map( A => DATAIN(2), ZN => n747);
   U626 : INV_X1 port map( A => DATAIN(3), ZN => n749);
   U627 : INV_X1 port map( A => DATAIN(4), ZN => n751);
   U628 : INV_X1 port map( A => DATAIN(5), ZN => n753);
   U629 : INV_X1 port map( A => DATAIN(6), ZN => n755);
   U630 : INV_X1 port map( A => DATAIN(7), ZN => n757);
   U631 : INV_X1 port map( A => DATAIN(8), ZN => n759);
   U632 : INV_X1 port map( A => DATAIN(9), ZN => n761);
   U633 : INV_X1 port map( A => DATAIN(10), ZN => n763);
   U634 : INV_X1 port map( A => DATAIN(11), ZN => n765);
   U635 : INV_X1 port map( A => DATAIN(12), ZN => n767);
   U636 : INV_X1 port map( A => DATAIN(13), ZN => n769);
   U637 : INV_X1 port map( A => DATAIN(14), ZN => n771);
   U638 : INV_X1 port map( A => DATAIN(15), ZN => n773);
   U639 : INV_X1 port map( A => DATAIN(16), ZN => n775);
   U640 : INV_X1 port map( A => DATAIN(17), ZN => n777);
   U641 : INV_X1 port map( A => DATAIN(18), ZN => n779);
   U642 : INV_X1 port map( A => DATAIN(19), ZN => n781);
   U643 : INV_X1 port map( A => DATAIN(20), ZN => n783);
   U644 : INV_X1 port map( A => DATAIN(21), ZN => n785);
   U645 : INV_X1 port map( A => DATAIN(22), ZN => n787);
   U646 : INV_X1 port map( A => DATAIN(23), ZN => n789);
   U647 : INV_X1 port map( A => DATAIN(24), ZN => n791);
   U648 : INV_X1 port map( A => DATAIN(25), ZN => n793);
   U649 : INV_X1 port map( A => DATAIN(26), ZN => n795);
   U650 : INV_X1 port map( A => DATAIN(27), ZN => n797);
   U651 : INV_X1 port map( A => DATAIN(28), ZN => n799);
   U652 : INV_X1 port map( A => DATAIN(29), ZN => n801);
   U653 : INV_X1 port map( A => DATAIN(30), ZN => n803);
   U654 : INV_X1 port map( A => DATAIN(31), ZN => n805);
   U655 : INV_X1 port map( A => DATAIN(32), ZN => n807);
   U656 : INV_X1 port map( A => DATAIN(33), ZN => n809);
   U657 : INV_X1 port map( A => DATAIN(34), ZN => n811);
   U658 : INV_X1 port map( A => DATAIN(35), ZN => n813);
   U659 : INV_X1 port map( A => DATAIN(36), ZN => n815);
   U660 : INV_X1 port map( A => DATAIN(37), ZN => n817);
   U661 : INV_X1 port map( A => DATAIN(38), ZN => n819);
   U662 : INV_X1 port map( A => DATAIN(39), ZN => n821);
   U663 : INV_X1 port map( A => DATAIN(40), ZN => n823);
   U664 : INV_X1 port map( A => DATAIN(41), ZN => n825);
   U665 : INV_X1 port map( A => DATAIN(42), ZN => n827);
   U666 : INV_X1 port map( A => DATAIN(43), ZN => n829);
   U667 : INV_X1 port map( A => DATAIN(44), ZN => n831);
   U668 : INV_X1 port map( A => DATAIN(45), ZN => n833);
   U669 : INV_X1 port map( A => DATAIN(46), ZN => n835);
   U670 : INV_X1 port map( A => DATAIN(47), ZN => n837);
   U671 : INV_X1 port map( A => DATAIN(48), ZN => n839);
   U672 : INV_X1 port map( A => DATAIN(49), ZN => n841);
   U673 : INV_X1 port map( A => DATAIN(50), ZN => n843);
   U674 : INV_X1 port map( A => DATAIN(51), ZN => n845);
   U675 : INV_X1 port map( A => DATAIN(52), ZN => n847);
   U676 : INV_X1 port map( A => DATAIN(53), ZN => n849);
   U677 : INV_X1 port map( A => DATAIN(54), ZN => n851);
   U678 : INV_X1 port map( A => DATAIN(55), ZN => n853);
   U679 : INV_X1 port map( A => DATAIN(56), ZN => n855);
   U680 : INV_X1 port map( A => DATAIN(57), ZN => n857);
   U681 : INV_X1 port map( A => DATAIN(58), ZN => n859);
   U682 : INV_X1 port map( A => DATAIN(59), ZN => n861);
   U683 : INV_X1 port map( A => DATAIN(60), ZN => n863);
   U684 : INV_X1 port map( A => DATAIN(61), ZN => n865);
   U685 : INV_X1 port map( A => DATAIN(62), ZN => n867);
   U686 : INV_X1 port map( A => DATAIN(63), ZN => n871);
   U687 : CLKBUF_X1 port map( A => n979, Z => n2069);
   U688 : CLKBUF_X1 port map( A => n978, Z => n2075);
   U689 : CLKBUF_X1 port map( A => n939, Z => n2081);
   U690 : CLKBUF_X1 port map( A => n938, Z => n2087);
   U691 : CLKBUF_X1 port map( A => n876, Z => n2093);
   U692 : CLKBUF_X1 port map( A => n875, Z => n2099);
   U693 : CLKBUF_X1 port map( A => n742, Z => n2105);
   U694 : CLKBUF_X1 port map( A => n741, Z => n2111);
   U695 : CLKBUF_X1 port map( A => n740, Z => n2117);
   U696 : CLKBUF_X1 port map( A => n739, Z => n2123);
   U697 : CLKBUF_X1 port map( A => n738, Z => n2129);
   U698 : CLKBUF_X1 port map( A => n736, Z => n2135);
   U699 : CLKBUF_X1 port map( A => n735, Z => n2141);
   U700 : CLKBUF_X1 port map( A => n527, Z => n2147);
   U701 : CLKBUF_X1 port map( A => n525, Z => n2158);
   U702 : CLKBUF_X1 port map( A => n523, Z => n2164);
   U703 : CLKBUF_X1 port map( A => n521, Z => n2170);
   U704 : INV_X1 port map( A => ADD_RD2(0), ZN => n2171);
   U705 : INV_X1 port map( A => ADD_RD2(1), ZN => n2172);
   U706 : INV_X1 port map( A => ADD_RD1(0), ZN => n2173);
   U707 : INV_X1 port map( A => ADD_RD1(1), ZN => n2174);
   U708 : INV_X1 port map( A => ADD_WR(0), ZN => n2175);
   U709 : INV_X1 port map( A => ADD_WR(1), ZN => n2176);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4.all;

entity register_file_reg_size64_file_size4_0 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
         std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector (63
         downto 0));

end register_file_reg_size64_file_size4_0;

architecture SYN_BEHAVIORAL of register_file_reg_size64_file_size4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426, 
      n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, 
      n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, 
      n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, 
      n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, 
      n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486, 
      n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, 
      n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510, 
      n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, 
      n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, 
      n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, 
      n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558, 
      n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, 
      n571, n572, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, 
      n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, 
      n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, 
      n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653, 
      n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664, n665, 
      n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, 
      n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, 
      n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, 
      n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, 
      n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, 
      n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, 
      n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, 
      n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761, 
      n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, 
      n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785, 
      n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796, n797, 
      n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, 
      n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, 
      n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833, 
      n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, 
      n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, 
      n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, 
      n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, 
      n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893, 
      n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, 
      n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, 
      n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929, 
      n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, 
      n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, 
      n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965, 
      n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, 
      n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, 
      n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
      n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, 
      n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, 
      n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, 
      n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, 
      n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, 
      n1052, n1053, n1054, n1055, n1163, n1165, n1183, n2, n3, n4, n5, n6, n7, 
      n8, n9, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, 
      n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39
      , n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, 
      n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68
      , n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, 
      n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97
      , n98, n99, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296
      , n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, 
      n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, 
      n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, 
      n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, 
      n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, 
      n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, 
      n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, 
      n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, 
      n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, 
      n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1395, n1396, n1397, 
      n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, 
      n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, 
      n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, 
      n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, 
      n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, 
      n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, 
      n1458, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, 
      n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, 
      n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, 
      n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, 
      n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, 
      n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, 
      n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, 
      n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, 
      n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, 
      n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, 
      n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, 
      n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, 
      n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, 
      n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, 
      n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, 
      n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, 
      n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, 
      n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, 
      n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, 
      n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, 
      n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, 
      n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, 
      n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, 
      n1689, n1690, n1691, n1694, n1695, n1696, n1697, n1698, n1699, n1700, 
      n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, 
      n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, 
      n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, 
      n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, 
      n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, 
      n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, 
      n1761, n1762, n1765, n1799, n1800, n1801, n1802, n1803, n1804, n1805, 
      n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, 
      n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, 
      n1826, n1827, n1828, n1829, n415, n573, n574, n575, n576, n577, n578, 
      n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, 
      n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, 
      n603, n604, n605, n606, n607, n1056, n1057, n1058, n1059, n1060, n1061, 
      n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, 
      n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, 
      n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, 
      n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, 
      n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, 
      n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, 
      n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, 
      n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, 
      n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, 
      n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, 
      n1162, n1164, n1166, n1167, n1168, n1169, n1170, n1171 : std_logic;

begin
   
   OUT2_reg_63_inst : DFF_X1 port map( D => n862, CK => CLK, Q => OUT2(63), QN 
                           => n543);
   OUT2_reg_62_inst : DFF_X1 port map( D => n860, CK => CLK, Q => OUT2(62), QN 
                           => n542);
   OUT2_reg_61_inst : DFF_X1 port map( D => n858, CK => CLK, Q => OUT2(61), QN 
                           => n541);
   OUT2_reg_60_inst : DFF_X1 port map( D => n856, CK => CLK, Q => OUT2(60), QN 
                           => n540);
   OUT2_reg_59_inst : DFF_X1 port map( D => n854, CK => CLK, Q => OUT2(59), QN 
                           => n539);
   OUT2_reg_58_inst : DFF_X1 port map( D => n852, CK => CLK, Q => OUT2(58), QN 
                           => n538);
   OUT2_reg_57_inst : DFF_X1 port map( D => n850, CK => CLK, Q => OUT2(57), QN 
                           => n537);
   OUT2_reg_56_inst : DFF_X1 port map( D => n848, CK => CLK, Q => OUT2(56), QN 
                           => n536);
   OUT2_reg_55_inst : DFF_X1 port map( D => n846, CK => CLK, Q => OUT2(55), QN 
                           => n535);
   OUT2_reg_54_inst : DFF_X1 port map( D => n844, CK => CLK, Q => OUT2(54), QN 
                           => n534);
   OUT2_reg_53_inst : DFF_X1 port map( D => n842, CK => CLK, Q => OUT2(53), QN 
                           => n533);
   OUT2_reg_52_inst : DFF_X1 port map( D => n840, CK => CLK, Q => OUT2(52), QN 
                           => n532);
   OUT2_reg_51_inst : DFF_X1 port map( D => n838, CK => CLK, Q => OUT2(51), QN 
                           => n531);
   OUT2_reg_50_inst : DFF_X1 port map( D => n836, CK => CLK, Q => OUT2(50), QN 
                           => n530);
   OUT2_reg_49_inst : DFF_X1 port map( D => n834, CK => CLK, Q => OUT2(49), QN 
                           => n529);
   OUT2_reg_48_inst : DFF_X1 port map( D => n832, CK => CLK, Q => OUT2(48), QN 
                           => n528);
   OUT2_reg_47_inst : DFF_X1 port map( D => n830, CK => CLK, Q => OUT2(47), QN 
                           => n527);
   OUT2_reg_46_inst : DFF_X1 port map( D => n828, CK => CLK, Q => OUT2(46), QN 
                           => n526);
   OUT2_reg_45_inst : DFF_X1 port map( D => n826, CK => CLK, Q => OUT2(45), QN 
                           => n525);
   OUT2_reg_44_inst : DFF_X1 port map( D => n824, CK => CLK, Q => OUT2(44), QN 
                           => n524);
   OUT2_reg_43_inst : DFF_X1 port map( D => n822, CK => CLK, Q => OUT2(43), QN 
                           => n523);
   OUT2_reg_42_inst : DFF_X1 port map( D => n820, CK => CLK, Q => OUT2(42), QN 
                           => n522);
   OUT2_reg_41_inst : DFF_X1 port map( D => n818, CK => CLK, Q => OUT2(41), QN 
                           => n521);
   OUT2_reg_40_inst : DFF_X1 port map( D => n816, CK => CLK, Q => OUT2(40), QN 
                           => n520);
   OUT2_reg_39_inst : DFF_X1 port map( D => n814, CK => CLK, Q => OUT2(39), QN 
                           => n519);
   OUT2_reg_38_inst : DFF_X1 port map( D => n812, CK => CLK, Q => OUT2(38), QN 
                           => n518);
   OUT2_reg_37_inst : DFF_X1 port map( D => n810, CK => CLK, Q => OUT2(37), QN 
                           => n517);
   OUT2_reg_36_inst : DFF_X1 port map( D => n808, CK => CLK, Q => OUT2(36), QN 
                           => n516);
   OUT2_reg_35_inst : DFF_X1 port map( D => n806, CK => CLK, Q => OUT2(35), QN 
                           => n515);
   OUT2_reg_34_inst : DFF_X1 port map( D => n804, CK => CLK, Q => OUT2(34), QN 
                           => n514);
   OUT2_reg_33_inst : DFF_X1 port map( D => n802, CK => CLK, Q => OUT2(33), QN 
                           => n513);
   OUT2_reg_32_inst : DFF_X1 port map( D => n800, CK => CLK, Q => OUT2(32), QN 
                           => n512);
   OUT2_reg_31_inst : DFF_X1 port map( D => n798, CK => CLK, Q => OUT2(31), QN 
                           => n511);
   REGISTERS_reg_3_30_inst : DFF_X1 port map( D => n797, CK => CLK, Q => n1799,
                           QN => n1569);
   OUT2_reg_30_inst : DFF_X1 port map( D => n796, CK => CLK, Q => OUT2(30), QN 
                           => n510);
   REGISTERS_reg_3_29_inst : DFF_X1 port map( D => n795, CK => CLK, Q => n1800,
                           QN => n1572);
   OUT2_reg_29_inst : DFF_X1 port map( D => n794, CK => CLK, Q => OUT2(29), QN 
                           => n509);
   REGISTERS_reg_3_28_inst : DFF_X1 port map( D => n793, CK => CLK, Q => n1801,
                           QN => n1575);
   OUT2_reg_28_inst : DFF_X1 port map( D => n792, CK => CLK, Q => OUT2(28), QN 
                           => n508);
   REGISTERS_reg_3_27_inst : DFF_X1 port map( D => n791, CK => CLK, Q => n1802,
                           QN => n1579);
   OUT2_reg_27_inst : DFF_X1 port map( D => n790, CK => CLK, Q => OUT2(27), QN 
                           => n507);
   REGISTERS_reg_3_26_inst : DFF_X1 port map( D => n789, CK => CLK, Q => n1803,
                           QN => n1583);
   OUT2_reg_26_inst : DFF_X1 port map( D => n788, CK => CLK, Q => OUT2(26), QN 
                           => n506);
   REGISTERS_reg_3_25_inst : DFF_X1 port map( D => n787, CK => CLK, Q => n1804,
                           QN => n1587);
   OUT2_reg_25_inst : DFF_X1 port map( D => n786, CK => CLK, Q => OUT2(25), QN 
                           => n505);
   REGISTERS_reg_3_24_inst : DFF_X1 port map( D => n785, CK => CLK, Q => n1805,
                           QN => n1591);
   OUT2_reg_24_inst : DFF_X1 port map( D => n784, CK => CLK, Q => OUT2(24), QN 
                           => n504);
   REGISTERS_reg_3_23_inst : DFF_X1 port map( D => n783, CK => CLK, Q => n1806,
                           QN => n1595);
   OUT2_reg_23_inst : DFF_X1 port map( D => n782, CK => CLK, Q => OUT2(23), QN 
                           => n503);
   REGISTERS_reg_3_22_inst : DFF_X1 port map( D => n781, CK => CLK, Q => n1807,
                           QN => n1599);
   OUT2_reg_22_inst : DFF_X1 port map( D => n780, CK => CLK, Q => OUT2(22), QN 
                           => n502);
   REGISTERS_reg_3_21_inst : DFF_X1 port map( D => n779, CK => CLK, Q => n1808,
                           QN => n1603);
   OUT2_reg_21_inst : DFF_X1 port map( D => n778, CK => CLK, Q => OUT2(21), QN 
                           => n501);
   REGISTERS_reg_3_20_inst : DFF_X1 port map( D => n777, CK => CLK, Q => n1809,
                           QN => n1607);
   OUT2_reg_20_inst : DFF_X1 port map( D => n776, CK => CLK, Q => OUT2(20), QN 
                           => n500);
   REGISTERS_reg_3_19_inst : DFF_X1 port map( D => n775, CK => CLK, Q => n1810,
                           QN => n1611);
   OUT2_reg_19_inst : DFF_X1 port map( D => n774, CK => CLK, Q => OUT2(19), QN 
                           => n499);
   REGISTERS_reg_3_18_inst : DFF_X1 port map( D => n773, CK => CLK, Q => n1811,
                           QN => n1615);
   OUT2_reg_18_inst : DFF_X1 port map( D => n772, CK => CLK, Q => OUT2(18), QN 
                           => n498);
   REGISTERS_reg_3_17_inst : DFF_X1 port map( D => n771, CK => CLK, Q => n1812,
                           QN => n1619);
   OUT2_reg_17_inst : DFF_X1 port map( D => n770, CK => CLK, Q => OUT2(17), QN 
                           => n497);
   REGISTERS_reg_3_16_inst : DFF_X1 port map( D => n769, CK => CLK, Q => n1813,
                           QN => n1623);
   OUT2_reg_16_inst : DFF_X1 port map( D => n768, CK => CLK, Q => OUT2(16), QN 
                           => n496);
   REGISTERS_reg_3_15_inst : DFF_X1 port map( D => n767, CK => CLK, Q => n1814,
                           QN => n1627);
   OUT2_reg_15_inst : DFF_X1 port map( D => n766, CK => CLK, Q => OUT2(15), QN 
                           => n495);
   REGISTERS_reg_3_14_inst : DFF_X1 port map( D => n765, CK => CLK, Q => n1815,
                           QN => n1631);
   OUT2_reg_14_inst : DFF_X1 port map( D => n764, CK => CLK, Q => OUT2(14), QN 
                           => n494);
   REGISTERS_reg_3_13_inst : DFF_X1 port map( D => n763, CK => CLK, Q => n1816,
                           QN => n1635);
   OUT2_reg_13_inst : DFF_X1 port map( D => n762, CK => CLK, Q => OUT2(13), QN 
                           => n493);
   REGISTERS_reg_3_12_inst : DFF_X1 port map( D => n761, CK => CLK, Q => n1817,
                           QN => n1639);
   OUT2_reg_12_inst : DFF_X1 port map( D => n760, CK => CLK, Q => OUT2(12), QN 
                           => n492);
   REGISTERS_reg_3_11_inst : DFF_X1 port map( D => n759, CK => CLK, Q => n1818,
                           QN => n1643);
   OUT2_reg_11_inst : DFF_X1 port map( D => n758, CK => CLK, Q => OUT2(11), QN 
                           => n491);
   REGISTERS_reg_3_10_inst : DFF_X1 port map( D => n757, CK => CLK, Q => n1819,
                           QN => n1647);
   OUT2_reg_10_inst : DFF_X1 port map( D => n756, CK => CLK, Q => OUT2(10), QN 
                           => n490);
   REGISTERS_reg_3_9_inst : DFF_X1 port map( D => n755, CK => CLK, Q => n1820, 
                           QN => n1651);
   OUT2_reg_9_inst : DFF_X1 port map( D => n754, CK => CLK, Q => OUT2(9), QN =>
                           n489);
   REGISTERS_reg_3_8_inst : DFF_X1 port map( D => n753, CK => CLK, Q => n1821, 
                           QN => n1655);
   OUT2_reg_8_inst : DFF_X1 port map( D => n752, CK => CLK, Q => OUT2(8), QN =>
                           n488);
   REGISTERS_reg_3_7_inst : DFF_X1 port map( D => n751, CK => CLK, Q => n1822, 
                           QN => n1659);
   OUT2_reg_7_inst : DFF_X1 port map( D => n750, CK => CLK, Q => OUT2(7), QN =>
                           n487);
   REGISTERS_reg_3_6_inst : DFF_X1 port map( D => n749, CK => CLK, Q => n1823, 
                           QN => n1663);
   OUT2_reg_6_inst : DFF_X1 port map( D => n748, CK => CLK, Q => OUT2(6), QN =>
                           n486);
   REGISTERS_reg_3_5_inst : DFF_X1 port map( D => n747, CK => CLK, Q => n1824, 
                           QN => n1667);
   OUT2_reg_5_inst : DFF_X1 port map( D => n746, CK => CLK, Q => OUT2(5), QN =>
                           n485);
   REGISTERS_reg_3_4_inst : DFF_X1 port map( D => n745, CK => CLK, Q => n1825, 
                           QN => n1671);
   OUT2_reg_4_inst : DFF_X1 port map( D => n744, CK => CLK, Q => OUT2(4), QN =>
                           n484);
   REGISTERS_reg_3_3_inst : DFF_X1 port map( D => n743, CK => CLK, Q => n1826, 
                           QN => n1675);
   OUT2_reg_3_inst : DFF_X1 port map( D => n742, CK => CLK, Q => OUT2(3), QN =>
                           n483);
   REGISTERS_reg_3_2_inst : DFF_X1 port map( D => n741, CK => CLK, Q => n1827, 
                           QN => n1679);
   OUT2_reg_2_inst : DFF_X1 port map( D => n740, CK => CLK, Q => OUT2(2), QN =>
                           n482);
   REGISTERS_reg_3_1_inst : DFF_X1 port map( D => n739, CK => CLK, Q => n1828, 
                           QN => n1683);
   OUT2_reg_1_inst : DFF_X1 port map( D => n738, CK => CLK, Q => OUT2(1), QN =>
                           n481);
   REGISTERS_reg_3_0_inst : DFF_X1 port map( D => n737, CK => CLK, Q => n1829, 
                           QN => n1687);
   OUT2_reg_0_inst : DFF_X1 port map( D => n736, CK => CLK, Q => OUT2(0), QN =>
                           n480);
   OUT1_reg_63_inst : DFF_X1 port map( D => n735, CK => CLK, Q => OUT1(63), QN 
                           => n479);
   OUT1_reg_62_inst : DFF_X1 port map( D => n734, CK => CLK, Q => OUT1(62), QN 
                           => n478);
   OUT1_reg_61_inst : DFF_X1 port map( D => n733, CK => CLK, Q => OUT1(61), QN 
                           => n477);
   OUT1_reg_60_inst : DFF_X1 port map( D => n732, CK => CLK, Q => OUT1(60), QN 
                           => n476);
   OUT1_reg_59_inst : DFF_X1 port map( D => n731, CK => CLK, Q => OUT1(59), QN 
                           => n475);
   OUT1_reg_58_inst : DFF_X1 port map( D => n730, CK => CLK, Q => OUT1(58), QN 
                           => n474);
   OUT1_reg_57_inst : DFF_X1 port map( D => n729, CK => CLK, Q => OUT1(57), QN 
                           => n473);
   OUT1_reg_56_inst : DFF_X1 port map( D => n728, CK => CLK, Q => OUT1(56), QN 
                           => n472);
   OUT1_reg_55_inst : DFF_X1 port map( D => n727, CK => CLK, Q => OUT1(55), QN 
                           => n471);
   OUT1_reg_54_inst : DFF_X1 port map( D => n726, CK => CLK, Q => OUT1(54), QN 
                           => n470);
   OUT1_reg_53_inst : DFF_X1 port map( D => n725, CK => CLK, Q => OUT1(53), QN 
                           => n469);
   OUT1_reg_52_inst : DFF_X1 port map( D => n724, CK => CLK, Q => OUT1(52), QN 
                           => n468);
   OUT1_reg_51_inst : DFF_X1 port map( D => n723, CK => CLK, Q => OUT1(51), QN 
                           => n467);
   OUT1_reg_50_inst : DFF_X1 port map( D => n722, CK => CLK, Q => OUT1(50), QN 
                           => n466);
   OUT1_reg_49_inst : DFF_X1 port map( D => n721, CK => CLK, Q => OUT1(49), QN 
                           => n465);
   OUT1_reg_48_inst : DFF_X1 port map( D => n720, CK => CLK, Q => OUT1(48), QN 
                           => n464);
   OUT1_reg_47_inst : DFF_X1 port map( D => n719, CK => CLK, Q => OUT1(47), QN 
                           => n463);
   OUT1_reg_46_inst : DFF_X1 port map( D => n718, CK => CLK, Q => OUT1(46), QN 
                           => n462);
   OUT1_reg_45_inst : DFF_X1 port map( D => n717, CK => CLK, Q => OUT1(45), QN 
                           => n461);
   OUT1_reg_44_inst : DFF_X1 port map( D => n716, CK => CLK, Q => OUT1(44), QN 
                           => n460);
   OUT1_reg_43_inst : DFF_X1 port map( D => n715, CK => CLK, Q => OUT1(43), QN 
                           => n459);
   OUT1_reg_42_inst : DFF_X1 port map( D => n714, CK => CLK, Q => OUT1(42), QN 
                           => n458);
   OUT1_reg_41_inst : DFF_X1 port map( D => n713, CK => CLK, Q => OUT1(41), QN 
                           => n457);
   OUT1_reg_40_inst : DFF_X1 port map( D => n712, CK => CLK, Q => OUT1(40), QN 
                           => n456);
   OUT1_reg_39_inst : DFF_X1 port map( D => n711, CK => CLK, Q => OUT1(39), QN 
                           => n455);
   OUT1_reg_38_inst : DFF_X1 port map( D => n710, CK => CLK, Q => OUT1(38), QN 
                           => n454);
   OUT1_reg_37_inst : DFF_X1 port map( D => n709, CK => CLK, Q => OUT1(37), QN 
                           => n453);
   OUT1_reg_36_inst : DFF_X1 port map( D => n708, CK => CLK, Q => OUT1(36), QN 
                           => n452);
   OUT1_reg_35_inst : DFF_X1 port map( D => n707, CK => CLK, Q => OUT1(35), QN 
                           => n451);
   OUT1_reg_34_inst : DFF_X1 port map( D => n706, CK => CLK, Q => OUT1(34), QN 
                           => n450);
   OUT1_reg_33_inst : DFF_X1 port map( D => n705, CK => CLK, Q => OUT1(33), QN 
                           => n449);
   OUT1_reg_32_inst : DFF_X1 port map( D => n704, CK => CLK, Q => OUT1(32), QN 
                           => n448);
   OUT1_reg_31_inst : DFF_X1 port map( D => n703, CK => CLK, Q => OUT1(31), QN 
                           => n447);
   OUT1_reg_30_inst : DFF_X1 port map( D => n702, CK => CLK, Q => OUT1(30), QN 
                           => n446);
   OUT1_reg_29_inst : DFF_X1 port map( D => n701, CK => CLK, Q => OUT1(29), QN 
                           => n445);
   OUT1_reg_28_inst : DFF_X1 port map( D => n700, CK => CLK, Q => OUT1(28), QN 
                           => n444);
   OUT1_reg_27_inst : DFF_X1 port map( D => n699, CK => CLK, Q => OUT1(27), QN 
                           => n443);
   OUT1_reg_26_inst : DFF_X1 port map( D => n698, CK => CLK, Q => OUT1(26), QN 
                           => n442);
   OUT1_reg_25_inst : DFF_X1 port map( D => n697, CK => CLK, Q => OUT1(25), QN 
                           => n441);
   OUT1_reg_24_inst : DFF_X1 port map( D => n696, CK => CLK, Q => OUT1(24), QN 
                           => n440);
   OUT1_reg_23_inst : DFF_X1 port map( D => n695, CK => CLK, Q => OUT1(23), QN 
                           => n439);
   OUT1_reg_22_inst : DFF_X1 port map( D => n694, CK => CLK, Q => OUT1(22), QN 
                           => n438);
   OUT1_reg_21_inst : DFF_X1 port map( D => n693, CK => CLK, Q => OUT1(21), QN 
                           => n437);
   OUT1_reg_20_inst : DFF_X1 port map( D => n692, CK => CLK, Q => OUT1(20), QN 
                           => n436);
   OUT1_reg_19_inst : DFF_X1 port map( D => n691, CK => CLK, Q => OUT1(19), QN 
                           => n435);
   OUT1_reg_18_inst : DFF_X1 port map( D => n690, CK => CLK, Q => OUT1(18), QN 
                           => n434);
   OUT1_reg_17_inst : DFF_X1 port map( D => n689, CK => CLK, Q => OUT1(17), QN 
                           => n433);
   OUT1_reg_16_inst : DFF_X1 port map( D => n688, CK => CLK, Q => OUT1(16), QN 
                           => n432);
   OUT1_reg_15_inst : DFF_X1 port map( D => n687, CK => CLK, Q => OUT1(15), QN 
                           => n431);
   OUT1_reg_14_inst : DFF_X1 port map( D => n686, CK => CLK, Q => OUT1(14), QN 
                           => n430);
   OUT1_reg_13_inst : DFF_X1 port map( D => n685, CK => CLK, Q => OUT1(13), QN 
                           => n429);
   OUT1_reg_12_inst : DFF_X1 port map( D => n684, CK => CLK, Q => OUT1(12), QN 
                           => n428);
   OUT1_reg_11_inst : DFF_X1 port map( D => n683, CK => CLK, Q => OUT1(11), QN 
                           => n427);
   OUT1_reg_10_inst : DFF_X1 port map( D => n682, CK => CLK, Q => OUT1(10), QN 
                           => n426);
   OUT1_reg_9_inst : DFF_X1 port map( D => n681, CK => CLK, Q => OUT1(9), QN =>
                           n425);
   OUT1_reg_8_inst : DFF_X1 port map( D => n680, CK => CLK, Q => OUT1(8), QN =>
                           n424);
   OUT1_reg_7_inst : DFF_X1 port map( D => n679, CK => CLK, Q => OUT1(7), QN =>
                           n423);
   OUT1_reg_6_inst : DFF_X1 port map( D => n678, CK => CLK, Q => OUT1(6), QN =>
                           n422);
   OUT1_reg_5_inst : DFF_X1 port map( D => n677, CK => CLK, Q => OUT1(5), QN =>
                           n421);
   OUT1_reg_4_inst : DFF_X1 port map( D => n676, CK => CLK, Q => OUT1(4), QN =>
                           n420);
   OUT1_reg_3_inst : DFF_X1 port map( D => n675, CK => CLK, Q => OUT1(3), QN =>
                           n419);
   OUT1_reg_2_inst : DFF_X1 port map( D => n674, CK => CLK, Q => OUT1(2), QN =>
                           n418);
   OUT1_reg_1_inst : DFF_X1 port map( D => n673, CK => CLK, Q => OUT1(1), QN =>
                           n417);
   OUT1_reg_0_inst : DFF_X1 port map( D => n672, CK => CLK, Q => OUT1(0), QN =>
                           n416);
   U859 : NAND3_X1 port map( A1 => n1393, A2 => n1171, A3 => ADD_WR(0), ZN => 
                           n1392);
   U860 : NAND3_X1 port map( A1 => n1393, A2 => n1170, A3 => ADD_WR(1), ZN => 
                           n1458);
   U861 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n1393, A3 => ADD_WR(1), ZN 
                           => n1688);
   U862 : NAND3_X1 port map( A1 => ADD_RD2(0), A2 => n1106, A3 => ADD_RD2(1), 
                           ZN => n1463);
   U863 : NAND3_X1 port map( A1 => ADD_RD1(0), A2 => n1076, A3 => ADD_RD1(1), 
                           ZN => n1694);
   U864 : NAND3_X1 port map( A1 => n1170, A2 => n1171, A3 => n1393, ZN => n1765
                           );
   REGISTERS_reg_0_7_inst : DFF_X1 port map( D => n999, CK => CLK, Q => n1661, 
                           QN => n615);
   REGISTERS_reg_0_6_inst : DFF_X1 port map( D => n998, CK => CLK, Q => n1665, 
                           QN => n614);
   REGISTERS_reg_0_5_inst : DFF_X1 port map( D => n997, CK => CLK, Q => n1669, 
                           QN => n613);
   REGISTERS_reg_0_4_inst : DFF_X1 port map( D => n996, CK => CLK, Q => n1673, 
                           QN => n612);
   REGISTERS_reg_0_63_inst : DFF_X1 port map( D => n1055, CK => CLK, Q => n1469
                           , QN => n671);
   REGISTERS_reg_0_62_inst : DFF_X1 port map( D => n1054, CK => CLK, Q => n1473
                           , QN => n670);
   REGISTERS_reg_0_61_inst : DFF_X1 port map( D => n1053, CK => CLK, Q => n1476
                           , QN => n669);
   REGISTERS_reg_0_60_inst : DFF_X1 port map( D => n1052, CK => CLK, Q => n1479
                           , QN => n668);
   REGISTERS_reg_0_59_inst : DFF_X1 port map( D => n1051, CK => CLK, Q => n1482
                           , QN => n667);
   REGISTERS_reg_0_58_inst : DFF_X1 port map( D => n1050, CK => CLK, Q => n1485
                           , QN => n666);
   REGISTERS_reg_0_57_inst : DFF_X1 port map( D => n1049, CK => CLK, Q => n1488
                           , QN => n665);
   REGISTERS_reg_0_56_inst : DFF_X1 port map( D => n1048, CK => CLK, Q => n1491
                           , QN => n664);
   REGISTERS_reg_0_55_inst : DFF_X1 port map( D => n1047, CK => CLK, Q => n1494
                           , QN => n663);
   REGISTERS_reg_0_54_inst : DFF_X1 port map( D => n1046, CK => CLK, Q => n1498
                           , QN => n662);
   REGISTERS_reg_0_53_inst : DFF_X1 port map( D => n1045, CK => CLK, Q => n1502
                           , QN => n661);
   REGISTERS_reg_0_52_inst : DFF_X1 port map( D => n1044, CK => CLK, Q => n1505
                           , QN => n660);
   REGISTERS_reg_0_51_inst : DFF_X1 port map( D => n1043, CK => CLK, Q => n1508
                           , QN => n659);
   REGISTERS_reg_0_50_inst : DFF_X1 port map( D => n1042, CK => CLK, Q => n1511
                           , QN => n658);
   REGISTERS_reg_0_49_inst : DFF_X1 port map( D => n1041, CK => CLK, Q => n1514
                           , QN => n657);
   REGISTERS_reg_0_48_inst : DFF_X1 port map( D => n1040, CK => CLK, Q => n1517
                           , QN => n656);
   REGISTERS_reg_0_47_inst : DFF_X1 port map( D => n1039, CK => CLK, Q => n1520
                           , QN => n655);
   REGISTERS_reg_0_46_inst : DFF_X1 port map( D => n1038, CK => CLK, Q => n1523
                           , QN => n654);
   REGISTERS_reg_0_45_inst : DFF_X1 port map( D => n1037, CK => CLK, Q => n1526
                           , QN => n653);
   REGISTERS_reg_0_44_inst : DFF_X1 port map( D => n1036, CK => CLK, Q => n1529
                           , QN => n652);
   REGISTERS_reg_0_43_inst : DFF_X1 port map( D => n1035, CK => CLK, Q => n1532
                           , QN => n651);
   REGISTERS_reg_0_42_inst : DFF_X1 port map( D => n1034, CK => CLK, Q => n1535
                           , QN => n650);
   REGISTERS_reg_0_41_inst : DFF_X1 port map( D => n1033, CK => CLK, Q => n1538
                           , QN => n649);
   REGISTERS_reg_0_40_inst : DFF_X1 port map( D => n1032, CK => CLK, Q => n1541
                           , QN => n648);
   REGISTERS_reg_0_39_inst : DFF_X1 port map( D => n1031, CK => CLK, Q => n1544
                           , QN => n647);
   REGISTERS_reg_0_38_inst : DFF_X1 port map( D => n1030, CK => CLK, Q => n1547
                           , QN => n646);
   REGISTERS_reg_0_37_inst : DFF_X1 port map( D => n1029, CK => CLK, Q => n1550
                           , QN => n645);
   REGISTERS_reg_0_36_inst : DFF_X1 port map( D => n1028, CK => CLK, Q => n1553
                           , QN => n644);
   REGISTERS_reg_0_35_inst : DFF_X1 port map( D => n1027, CK => CLK, Q => n1556
                           , QN => n643);
   REGISTERS_reg_0_34_inst : DFF_X1 port map( D => n1026, CK => CLK, Q => n1559
                           , QN => n642);
   REGISTERS_reg_0_33_inst : DFF_X1 port map( D => n1025, CK => CLK, Q => n1562
                           , QN => n641);
   REGISTERS_reg_0_32_inst : DFF_X1 port map( D => n1024, CK => CLK, Q => n1565
                           , QN => n640);
   REGISTERS_reg_0_31_inst : DFF_X1 port map( D => n1023, CK => CLK, Q => n1568
                           , QN => n639);
   REGISTERS_reg_0_30_inst : DFF_X1 port map( D => n1022, CK => CLK, Q => n1571
                           , QN => n638);
   REGISTERS_reg_0_29_inst : DFF_X1 port map( D => n1021, CK => CLK, Q => n1574
                           , QN => n637);
   REGISTERS_reg_0_28_inst : DFF_X1 port map( D => n1020, CK => CLK, Q => n1577
                           , QN => n636);
   REGISTERS_reg_0_27_inst : DFF_X1 port map( D => n1019, CK => CLK, Q => n1581
                           , QN => n635);
   REGISTERS_reg_0_26_inst : DFF_X1 port map( D => n1018, CK => CLK, Q => n1585
                           , QN => n634);
   REGISTERS_reg_0_25_inst : DFF_X1 port map( D => n1017, CK => CLK, Q => n1589
                           , QN => n633);
   REGISTERS_reg_0_24_inst : DFF_X1 port map( D => n1016, CK => CLK, Q => n1593
                           , QN => n632);
   REGISTERS_reg_0_23_inst : DFF_X1 port map( D => n1015, CK => CLK, Q => n1597
                           , QN => n631);
   REGISTERS_reg_0_22_inst : DFF_X1 port map( D => n1014, CK => CLK, Q => n1601
                           , QN => n630);
   REGISTERS_reg_0_21_inst : DFF_X1 port map( D => n1013, CK => CLK, Q => n1605
                           , QN => n629);
   REGISTERS_reg_0_20_inst : DFF_X1 port map( D => n1012, CK => CLK, Q => n1609
                           , QN => n628);
   REGISTERS_reg_0_19_inst : DFF_X1 port map( D => n1011, CK => CLK, Q => n1613
                           , QN => n627);
   REGISTERS_reg_0_18_inst : DFF_X1 port map( D => n1010, CK => CLK, Q => n1617
                           , QN => n626);
   REGISTERS_reg_0_17_inst : DFF_X1 port map( D => n1009, CK => CLK, Q => n1621
                           , QN => n625);
   REGISTERS_reg_0_16_inst : DFF_X1 port map( D => n1008, CK => CLK, Q => n1625
                           , QN => n624);
   REGISTERS_reg_0_15_inst : DFF_X1 port map( D => n1007, CK => CLK, Q => n1629
                           , QN => n623);
   REGISTERS_reg_0_14_inst : DFF_X1 port map( D => n1006, CK => CLK, Q => n1633
                           , QN => n622);
   REGISTERS_reg_0_13_inst : DFF_X1 port map( D => n1005, CK => CLK, Q => n1637
                           , QN => n621);
   REGISTERS_reg_0_12_inst : DFF_X1 port map( D => n1004, CK => CLK, Q => n1641
                           , QN => n620);
   REGISTERS_reg_0_11_inst : DFF_X1 port map( D => n1003, CK => CLK, Q => n1645
                           , QN => n619);
   REGISTERS_reg_0_10_inst : DFF_X1 port map( D => n1002, CK => CLK, Q => n1649
                           , QN => n618);
   REGISTERS_reg_0_9_inst : DFF_X1 port map( D => n1001, CK => CLK, Q => n1653,
                           QN => n617);
   REGISTERS_reg_0_8_inst : DFF_X1 port map( D => n1000, CK => CLK, Q => n1657,
                           QN => n616);
   REGISTERS_reg_0_3_inst : DFF_X1 port map( D => n995, CK => CLK, Q => n1677, 
                           QN => n611);
   REGISTERS_reg_0_2_inst : DFF_X1 port map( D => n994, CK => CLK, Q => n1681, 
                           QN => n610);
   REGISTERS_reg_0_1_inst : DFF_X1 port map( D => n993, CK => CLK, Q => n1685, 
                           QN => n609);
   REGISTERS_reg_0_0_inst : DFF_X1 port map( D => n992, CK => CLK, Q => n1690, 
                           QN => n608);
   REGISTERS_reg_2_63_inst : DFF_X1 port map( D => n927, CK => CLK, Q => n1467,
                           QN => n1183);
   REGISTERS_reg_1_11_inst : DFF_X1 port map( D => n939, CK => CLK, Q => n1646,
                           QN => n555);
   REGISTERS_reg_1_10_inst : DFF_X1 port map( D => n938, CK => CLK, Q => n1650,
                           QN => n554);
   REGISTERS_reg_1_9_inst : DFF_X1 port map( D => n937, CK => CLK, Q => n1654, 
                           QN => n553);
   REGISTERS_reg_1_8_inst : DFF_X1 port map( D => n936, CK => CLK, Q => n1658, 
                           QN => n552);
   REGISTERS_reg_1_7_inst : DFF_X1 port map( D => n935, CK => CLK, Q => n1662, 
                           QN => n551);
   REGISTERS_reg_1_6_inst : DFF_X1 port map( D => n934, CK => CLK, Q => n1666, 
                           QN => n550);
   REGISTERS_reg_1_5_inst : DFF_X1 port map( D => n933, CK => CLK, Q => n1670, 
                           QN => n549);
   REGISTERS_reg_1_4_inst : DFF_X1 port map( D => n932, CK => CLK, Q => n1674, 
                           QN => n548);
   REGISTERS_reg_1_3_inst : DFF_X1 port map( D => n931, CK => CLK, Q => n1678, 
                           QN => n547);
   REGISTERS_reg_1_2_inst : DFF_X1 port map( D => n930, CK => CLK, Q => n1682, 
                           QN => n546);
   REGISTERS_reg_1_1_inst : DFF_X1 port map( D => n929, CK => CLK, Q => n1686, 
                           QN => n545);
   REGISTERS_reg_1_0_inst : DFF_X1 port map( D => n928, CK => CLK, Q => n1691, 
                           QN => n544);
   REGISTERS_reg_1_28_inst : DFF_X1 port map( D => n956, CK => CLK, Q => n1578,
                           QN => n572);
   REGISTERS_reg_1_27_inst : DFF_X1 port map( D => n955, CK => CLK, Q => n1582,
                           QN => n571);
   REGISTERS_reg_1_26_inst : DFF_X1 port map( D => n954, CK => CLK, Q => n1586,
                           QN => n570);
   REGISTERS_reg_1_25_inst : DFF_X1 port map( D => n953, CK => CLK, Q => n1590,
                           QN => n569);
   REGISTERS_reg_1_24_inst : DFF_X1 port map( D => n952, CK => CLK, Q => n1594,
                           QN => n568);
   REGISTERS_reg_1_23_inst : DFF_X1 port map( D => n951, CK => CLK, Q => n1598,
                           QN => n567);
   REGISTERS_reg_1_22_inst : DFF_X1 port map( D => n950, CK => CLK, Q => n1602,
                           QN => n566);
   REGISTERS_reg_1_21_inst : DFF_X1 port map( D => n949, CK => CLK, Q => n1606,
                           QN => n565);
   REGISTERS_reg_1_20_inst : DFF_X1 port map( D => n948, CK => CLK, Q => n1610,
                           QN => n564);
   REGISTERS_reg_1_19_inst : DFF_X1 port map( D => n947, CK => CLK, Q => n1614,
                           QN => n563);
   REGISTERS_reg_1_18_inst : DFF_X1 port map( D => n946, CK => CLK, Q => n1618,
                           QN => n562);
   REGISTERS_reg_1_17_inst : DFF_X1 port map( D => n945, CK => CLK, Q => n1622,
                           QN => n561);
   REGISTERS_reg_1_16_inst : DFF_X1 port map( D => n944, CK => CLK, Q => n1626,
                           QN => n560);
   REGISTERS_reg_1_15_inst : DFF_X1 port map( D => n943, CK => CLK, Q => n1630,
                           QN => n559);
   REGISTERS_reg_1_14_inst : DFF_X1 port map( D => n942, CK => CLK, Q => n1634,
                           QN => n558);
   REGISTERS_reg_1_13_inst : DFF_X1 port map( D => n941, CK => CLK, Q => n1638,
                           QN => n557);
   REGISTERS_reg_1_12_inst : DFF_X1 port map( D => n940, CK => CLK, Q => n1642,
                           QN => n556);
   REGISTERS_reg_2_54_inst : DFF_X1 port map( D => n918, CK => CLK, Q => n1497,
                           QN => n1165);
   REGISTERS_reg_2_53_inst : DFF_X1 port map( D => n917, CK => CLK, Q => n1501,
                           QN => n1163);
   REGISTERS_reg_2_62_inst : DFF_X1 port map( D => n926, CK => CLK, Q => n2, QN
                           => n1397);
   REGISTERS_reg_2_61_inst : DFF_X1 port map( D => n925, CK => CLK, Q => n3, QN
                           => n1398);
   REGISTERS_reg_2_60_inst : DFF_X1 port map( D => n924, CK => CLK, Q => n4, QN
                           => n1399);
   REGISTERS_reg_3_63_inst : DFF_X1 port map( D => n863, CK => CLK, Q => n604, 
                           QN => n1461);
   REGISTERS_reg_3_62_inst : DFF_X1 port map( D => n861, CK => CLK, Q => n603, 
                           QN => n1471);
   REGISTERS_reg_3_61_inst : DFF_X1 port map( D => n859, CK => CLK, Q => n602, 
                           QN => n1474);
   REGISTERS_reg_3_60_inst : DFF_X1 port map( D => n857, CK => CLK, Q => n601, 
                           QN => n1477);
   REGISTERS_reg_1_63_inst : DFF_X1 port map( D => n991, CK => CLK, Q => n65, 
                           QN => n1299);
   REGISTERS_reg_1_62_inst : DFF_X1 port map( D => n990, CK => CLK, Q => n66, 
                           QN => n1302);
   REGISTERS_reg_1_61_inst : DFF_X1 port map( D => n989, CK => CLK, Q => n67, 
                           QN => n1304);
   REGISTERS_reg_1_60_inst : DFF_X1 port map( D => n988, CK => CLK, Q => n68, 
                           QN => n1306);
   REGISTERS_reg_1_59_inst : DFF_X1 port map( D => n987, CK => CLK, Q => n69, 
                           QN => n1308);
   REGISTERS_reg_1_58_inst : DFF_X1 port map( D => n986, CK => CLK, Q => n70, 
                           QN => n1310);
   REGISTERS_reg_1_57_inst : DFF_X1 port map( D => n985, CK => CLK, Q => n71, 
                           QN => n1312);
   REGISTERS_reg_1_56_inst : DFF_X1 port map( D => n984, CK => CLK, Q => n72, 
                           QN => n1314);
   REGISTERS_reg_1_55_inst : DFF_X1 port map( D => n983, CK => CLK, Q => n73, 
                           QN => n1316);
   REGISTERS_reg_1_54_inst : DFF_X1 port map( D => n982, CK => CLK, Q => n74, 
                           QN => n1318);
   REGISTERS_reg_1_53_inst : DFF_X1 port map( D => n981, CK => CLK, Q => n75, 
                           QN => n1320);
   REGISTERS_reg_1_52_inst : DFF_X1 port map( D => n980, CK => CLK, Q => n76, 
                           QN => n1322);
   REGISTERS_reg_1_51_inst : DFF_X1 port map( D => n979, CK => CLK, Q => n77, 
                           QN => n1324);
   REGISTERS_reg_1_50_inst : DFF_X1 port map( D => n978, CK => CLK, Q => n78, 
                           QN => n1326);
   REGISTERS_reg_1_49_inst : DFF_X1 port map( D => n977, CK => CLK, Q => n79, 
                           QN => n1328);
   REGISTERS_reg_1_48_inst : DFF_X1 port map( D => n976, CK => CLK, Q => n80, 
                           QN => n1330);
   REGISTERS_reg_1_47_inst : DFF_X1 port map( D => n975, CK => CLK, Q => n81, 
                           QN => n1332);
   REGISTERS_reg_1_46_inst : DFF_X1 port map( D => n974, CK => CLK, Q => n82, 
                           QN => n1334);
   REGISTERS_reg_1_45_inst : DFF_X1 port map( D => n973, CK => CLK, Q => n83, 
                           QN => n1336);
   REGISTERS_reg_1_44_inst : DFF_X1 port map( D => n972, CK => CLK, Q => n84, 
                           QN => n1338);
   REGISTERS_reg_1_43_inst : DFF_X1 port map( D => n971, CK => CLK, Q => n85, 
                           QN => n1340);
   REGISTERS_reg_1_42_inst : DFF_X1 port map( D => n970, CK => CLK, Q => n86, 
                           QN => n1342);
   REGISTERS_reg_1_41_inst : DFF_X1 port map( D => n969, CK => CLK, Q => n87, 
                           QN => n1344);
   REGISTERS_reg_1_40_inst : DFF_X1 port map( D => n968, CK => CLK, Q => n88, 
                           QN => n1346);
   REGISTERS_reg_1_39_inst : DFF_X1 port map( D => n967, CK => CLK, Q => n89, 
                           QN => n1348);
   REGISTERS_reg_1_38_inst : DFF_X1 port map( D => n966, CK => CLK, Q => n90, 
                           QN => n1350);
   REGISTERS_reg_1_37_inst : DFF_X1 port map( D => n965, CK => CLK, Q => n91, 
                           QN => n1352);
   REGISTERS_reg_1_36_inst : DFF_X1 port map( D => n964, CK => CLK, Q => n92, 
                           QN => n1354);
   REGISTERS_reg_1_35_inst : DFF_X1 port map( D => n963, CK => CLK, Q => n93, 
                           QN => n1356);
   REGISTERS_reg_1_34_inst : DFF_X1 port map( D => n962, CK => CLK, Q => n94, 
                           QN => n1358);
   REGISTERS_reg_1_33_inst : DFF_X1 port map( D => n961, CK => CLK, Q => n95, 
                           QN => n1360);
   REGISTERS_reg_1_32_inst : DFF_X1 port map( D => n960, CK => CLK, Q => n96, 
                           QN => n1362);
   REGISTERS_reg_1_31_inst : DFF_X1 port map( D => n959, CK => CLK, Q => n97, 
                           QN => n1364);
   REGISTERS_reg_1_30_inst : DFF_X1 port map( D => n958, CK => CLK, Q => n98, 
                           QN => n1366);
   REGISTERS_reg_1_29_inst : DFF_X1 port map( D => n957, CK => CLK, Q => n99, 
                           QN => n1368);
   REGISTERS_reg_2_59_inst : DFF_X1 port map( D => n923, CK => CLK, Q => n5, QN
                           => n1400);
   REGISTERS_reg_2_58_inst : DFF_X1 port map( D => n922, CK => CLK, Q => n6, QN
                           => n1401);
   REGISTERS_reg_2_57_inst : DFF_X1 port map( D => n921, CK => CLK, Q => n7, QN
                           => n1402);
   REGISTERS_reg_2_56_inst : DFF_X1 port map( D => n920, CK => CLK, Q => n8, QN
                           => n1403);
   REGISTERS_reg_2_55_inst : DFF_X1 port map( D => n919, CK => CLK, Q => n9, QN
                           => n1404);
   REGISTERS_reg_2_52_inst : DFF_X1 port map( D => n916, CK => CLK, Q => n12, 
                           QN => n1405);
   REGISTERS_reg_2_51_inst : DFF_X1 port map( D => n915, CK => CLK, Q => n13, 
                           QN => n1406);
   REGISTERS_reg_2_50_inst : DFF_X1 port map( D => n914, CK => CLK, Q => n14, 
                           QN => n1407);
   REGISTERS_reg_2_49_inst : DFF_X1 port map( D => n913, CK => CLK, Q => n15, 
                           QN => n1408);
   REGISTERS_reg_2_48_inst : DFF_X1 port map( D => n912, CK => CLK, Q => n16, 
                           QN => n1409);
   REGISTERS_reg_2_47_inst : DFF_X1 port map( D => n911, CK => CLK, Q => n17, 
                           QN => n1410);
   REGISTERS_reg_2_46_inst : DFF_X1 port map( D => n910, CK => CLK, Q => n18, 
                           QN => n1411);
   REGISTERS_reg_2_45_inst : DFF_X1 port map( D => n909, CK => CLK, Q => n19, 
                           QN => n1412);
   REGISTERS_reg_2_44_inst : DFF_X1 port map( D => n908, CK => CLK, Q => n20, 
                           QN => n1413);
   REGISTERS_reg_2_43_inst : DFF_X1 port map( D => n907, CK => CLK, Q => n21, 
                           QN => n1414);
   REGISTERS_reg_2_42_inst : DFF_X1 port map( D => n906, CK => CLK, Q => n22, 
                           QN => n1415);
   REGISTERS_reg_2_41_inst : DFF_X1 port map( D => n905, CK => CLK, Q => n23, 
                           QN => n1416);
   REGISTERS_reg_2_40_inst : DFF_X1 port map( D => n904, CK => CLK, Q => n24, 
                           QN => n1417);
   REGISTERS_reg_2_39_inst : DFF_X1 port map( D => n903, CK => CLK, Q => n25, 
                           QN => n1418);
   REGISTERS_reg_2_38_inst : DFF_X1 port map( D => n902, CK => CLK, Q => n26, 
                           QN => n1419);
   REGISTERS_reg_2_37_inst : DFF_X1 port map( D => n901, CK => CLK, Q => n27, 
                           QN => n1420);
   REGISTERS_reg_2_36_inst : DFF_X1 port map( D => n900, CK => CLK, Q => n28, 
                           QN => n1421);
   REGISTERS_reg_2_35_inst : DFF_X1 port map( D => n899, CK => CLK, Q => n29, 
                           QN => n1422);
   REGISTERS_reg_2_34_inst : DFF_X1 port map( D => n898, CK => CLK, Q => n30, 
                           QN => n1423);
   REGISTERS_reg_2_33_inst : DFF_X1 port map( D => n897, CK => CLK, Q => n31, 
                           QN => n1424);
   REGISTERS_reg_2_32_inst : DFF_X1 port map( D => n896, CK => CLK, Q => n32, 
                           QN => n1425);
   REGISTERS_reg_2_31_inst : DFF_X1 port map( D => n895, CK => CLK, Q => n33, 
                           QN => n1426);
   REGISTERS_reg_2_30_inst : DFF_X1 port map( D => n894, CK => CLK, Q => n34, 
                           QN => n1427);
   REGISTERS_reg_2_29_inst : DFF_X1 port map( D => n893, CK => CLK, Q => n35, 
                           QN => n1428);
   REGISTERS_reg_2_28_inst : DFF_X1 port map( D => n892, CK => CLK, Q => n36, 
                           QN => n1429);
   REGISTERS_reg_2_27_inst : DFF_X1 port map( D => n891, CK => CLK, Q => n37, 
                           QN => n1430);
   REGISTERS_reg_2_26_inst : DFF_X1 port map( D => n890, CK => CLK, Q => n38, 
                           QN => n1431);
   REGISTERS_reg_2_25_inst : DFF_X1 port map( D => n889, CK => CLK, Q => n39, 
                           QN => n1432);
   REGISTERS_reg_2_24_inst : DFF_X1 port map( D => n888, CK => CLK, Q => n40, 
                           QN => n1433);
   REGISTERS_reg_2_23_inst : DFF_X1 port map( D => n887, CK => CLK, Q => n41, 
                           QN => n1434);
   REGISTERS_reg_2_22_inst : DFF_X1 port map( D => n886, CK => CLK, Q => n42, 
                           QN => n1435);
   REGISTERS_reg_2_21_inst : DFF_X1 port map( D => n885, CK => CLK, Q => n43, 
                           QN => n1436);
   REGISTERS_reg_2_20_inst : DFF_X1 port map( D => n884, CK => CLK, Q => n44, 
                           QN => n1437);
   REGISTERS_reg_2_19_inst : DFF_X1 port map( D => n883, CK => CLK, Q => n45, 
                           QN => n1438);
   REGISTERS_reg_2_18_inst : DFF_X1 port map( D => n882, CK => CLK, Q => n46, 
                           QN => n1439);
   REGISTERS_reg_2_17_inst : DFF_X1 port map( D => n881, CK => CLK, Q => n47, 
                           QN => n1440);
   REGISTERS_reg_2_16_inst : DFF_X1 port map( D => n880, CK => CLK, Q => n48, 
                           QN => n1441);
   REGISTERS_reg_2_15_inst : DFF_X1 port map( D => n879, CK => CLK, Q => n49, 
                           QN => n1442);
   REGISTERS_reg_2_14_inst : DFF_X1 port map( D => n878, CK => CLK, Q => n50, 
                           QN => n1443);
   REGISTERS_reg_2_13_inst : DFF_X1 port map( D => n877, CK => CLK, Q => n51, 
                           QN => n1444);
   REGISTERS_reg_2_12_inst : DFF_X1 port map( D => n876, CK => CLK, Q => n52, 
                           QN => n1445);
   REGISTERS_reg_2_11_inst : DFF_X1 port map( D => n875, CK => CLK, Q => n53, 
                           QN => n1446);
   REGISTERS_reg_2_10_inst : DFF_X1 port map( D => n874, CK => CLK, Q => n54, 
                           QN => n1447);
   REGISTERS_reg_2_9_inst : DFF_X1 port map( D => n873, CK => CLK, Q => n55, QN
                           => n1448);
   REGISTERS_reg_2_8_inst : DFF_X1 port map( D => n872, CK => CLK, Q => n56, QN
                           => n1449);
   REGISTERS_reg_2_7_inst : DFF_X1 port map( D => n871, CK => CLK, Q => n57, QN
                           => n1450);
   REGISTERS_reg_2_6_inst : DFF_X1 port map( D => n870, CK => CLK, Q => n58, QN
                           => n1451);
   REGISTERS_reg_2_5_inst : DFF_X1 port map( D => n869, CK => CLK, Q => n59, QN
                           => n1452);
   REGISTERS_reg_2_4_inst : DFF_X1 port map( D => n868, CK => CLK, Q => n60, QN
                           => n1453);
   REGISTERS_reg_2_3_inst : DFF_X1 port map( D => n867, CK => CLK, Q => n61, QN
                           => n1454);
   REGISTERS_reg_2_2_inst : DFF_X1 port map( D => n866, CK => CLK, Q => n62, QN
                           => n1455);
   REGISTERS_reg_2_1_inst : DFF_X1 port map( D => n865, CK => CLK, Q => n63, QN
                           => n1456);
   REGISTERS_reg_2_0_inst : DFF_X1 port map( D => n864, CK => CLK, Q => n64, QN
                           => n1457);
   REGISTERS_reg_3_59_inst : DFF_X1 port map( D => n855, CK => CLK, Q => n600, 
                           QN => n1480);
   REGISTERS_reg_3_58_inst : DFF_X1 port map( D => n853, CK => CLK, Q => n599, 
                           QN => n1483);
   REGISTERS_reg_3_57_inst : DFF_X1 port map( D => n851, CK => CLK, Q => n598, 
                           QN => n1486);
   REGISTERS_reg_3_56_inst : DFF_X1 port map( D => n849, CK => CLK, Q => n597, 
                           QN => n1489);
   REGISTERS_reg_3_55_inst : DFF_X1 port map( D => n847, CK => CLK, Q => n596, 
                           QN => n1492);
   REGISTERS_reg_3_54_inst : DFF_X1 port map( D => n845, CK => CLK, Q => n595, 
                           QN => n1495);
   REGISTERS_reg_3_53_inst : DFF_X1 port map( D => n843, CK => CLK, Q => n594, 
                           QN => n1499);
   REGISTERS_reg_3_52_inst : DFF_X1 port map( D => n841, CK => CLK, Q => n593, 
                           QN => n1503);
   REGISTERS_reg_3_51_inst : DFF_X1 port map( D => n839, CK => CLK, Q => n592, 
                           QN => n1506);
   REGISTERS_reg_3_50_inst : DFF_X1 port map( D => n837, CK => CLK, Q => n591, 
                           QN => n1509);
   REGISTERS_reg_3_49_inst : DFF_X1 port map( D => n835, CK => CLK, Q => n590, 
                           QN => n1512);
   REGISTERS_reg_3_48_inst : DFF_X1 port map( D => n833, CK => CLK, Q => n589, 
                           QN => n1515);
   REGISTERS_reg_3_47_inst : DFF_X1 port map( D => n831, CK => CLK, Q => n588, 
                           QN => n1518);
   REGISTERS_reg_3_46_inst : DFF_X1 port map( D => n829, CK => CLK, Q => n587, 
                           QN => n1521);
   REGISTERS_reg_3_45_inst : DFF_X1 port map( D => n827, CK => CLK, Q => n586, 
                           QN => n1524);
   REGISTERS_reg_3_44_inst : DFF_X1 port map( D => n825, CK => CLK, Q => n585, 
                           QN => n1527);
   REGISTERS_reg_3_43_inst : DFF_X1 port map( D => n823, CK => CLK, Q => n584, 
                           QN => n1530);
   REGISTERS_reg_3_42_inst : DFF_X1 port map( D => n821, CK => CLK, Q => n583, 
                           QN => n1533);
   REGISTERS_reg_3_41_inst : DFF_X1 port map( D => n819, CK => CLK, Q => n582, 
                           QN => n1536);
   REGISTERS_reg_3_40_inst : DFF_X1 port map( D => n817, CK => CLK, Q => n581, 
                           QN => n1539);
   REGISTERS_reg_3_39_inst : DFF_X1 port map( D => n815, CK => CLK, Q => n580, 
                           QN => n1542);
   REGISTERS_reg_3_38_inst : DFF_X1 port map( D => n813, CK => CLK, Q => n579, 
                           QN => n1545);
   REGISTERS_reg_3_37_inst : DFF_X1 port map( D => n811, CK => CLK, Q => n578, 
                           QN => n1548);
   REGISTERS_reg_3_36_inst : DFF_X1 port map( D => n809, CK => CLK, Q => n577, 
                           QN => n1551);
   REGISTERS_reg_3_35_inst : DFF_X1 port map( D => n807, CK => CLK, Q => n576, 
                           QN => n1554);
   REGISTERS_reg_3_34_inst : DFF_X1 port map( D => n805, CK => CLK, Q => n575, 
                           QN => n1557);
   REGISTERS_reg_3_33_inst : DFF_X1 port map( D => n803, CK => CLK, Q => n574, 
                           QN => n1560);
   REGISTERS_reg_3_32_inst : DFF_X1 port map( D => n801, CK => CLK, Q => n573, 
                           QN => n1563);
   REGISTERS_reg_3_31_inst : DFF_X1 port map( D => n799, CK => CLK, Q => n415, 
                           QN => n1566);
   U3 : BUF_X1 port map( A => n1463, Z => n1107);
   U4 : BUF_X1 port map( A => n1463, Z => n1108);
   U5 : BUF_X1 port map( A => n1463, Z => n1109);
   U6 : BUF_X1 port map( A => n1694, Z => n1077);
   U7 : BUF_X1 port map( A => n1694, Z => n1078);
   U8 : BUF_X1 port map( A => n1694, Z => n1079);
   U9 : BUF_X1 port map( A => n1694, Z => n1080);
   U10 : BUF_X1 port map( A => n1132, Z => n1134);
   U11 : BUF_X1 port map( A => n1139, Z => n1142);
   U12 : BUF_X1 port map( A => n1139, Z => n1143);
   U13 : BUF_X1 port map( A => n1140, Z => n1144);
   U14 : BUF_X1 port map( A => n1140, Z => n1145);
   U15 : BUF_X1 port map( A => n1463, Z => n1110);
   U16 : BUF_X1 port map( A => n1463, Z => n1111);
   U17 : BUF_X1 port map( A => n1119, Z => n1121);
   U18 : BUF_X1 port map( A => n1119, Z => n1122);
   U19 : BUF_X1 port map( A => n1119, Z => n1123);
   U20 : BUF_X1 port map( A => n1120, Z => n1124);
   U21 : BUF_X1 port map( A => n1120, Z => n1125);
   U22 : BUF_X1 port map( A => n1133, Z => n1138);
   U23 : BUF_X1 port map( A => n1133, Z => n1137);
   U24 : BUF_X1 port map( A => n1132, Z => n1136);
   U25 : BUF_X1 port map( A => n1132, Z => n1135);
   U26 : BUF_X1 port map( A => n1139, Z => n1141);
   U27 : BUF_X1 port map( A => n1694, Z => n1081);
   U28 : BUF_X1 port map( A => n1695, Z => n1075);
   U29 : BUF_X1 port map( A => n1695, Z => n1074);
   U30 : BUF_X1 port map( A => n1695, Z => n1073);
   U31 : BUF_X1 port map( A => n1695, Z => n1072);
   U32 : BUF_X1 port map( A => n1695, Z => n1071);
   U33 : BUF_X1 port map( A => n1697, Z => n1065);
   U34 : BUF_X1 port map( A => n1697, Z => n1066);
   U35 : BUF_X1 port map( A => n1697, Z => n1067);
   U36 : BUF_X1 port map( A => n1697, Z => n1068);
   U37 : BUF_X1 port map( A => n1697, Z => n1069);
   U38 : BUF_X1 port map( A => n1466, Z => n1095);
   U39 : BUF_X1 port map( A => n1466, Z => n1096);
   U40 : BUF_X1 port map( A => n1466, Z => n1097);
   U41 : BUF_X1 port map( A => n1466, Z => n1098);
   U42 : BUF_X1 port map( A => n1466, Z => n1099);
   U43 : BUF_X1 port map( A => n1289, Z => n1153);
   U44 : BUF_X1 port map( A => n1289, Z => n1154);
   U45 : BUF_X1 port map( A => n1289, Z => n1155);
   U46 : BUF_X1 port map( A => n1289, Z => n1156);
   U47 : BUF_X1 port map( A => n1698, Z => n1059);
   U48 : BUF_X1 port map( A => n1698, Z => n1060);
   U49 : BUF_X1 port map( A => n1698, Z => n1061);
   U50 : BUF_X1 port map( A => n1698, Z => n1062);
   U51 : BUF_X1 port map( A => n1698, Z => n1063);
   U52 : BUF_X1 port map( A => n1468, Z => n1089);
   U53 : BUF_X1 port map( A => n1468, Z => n1090);
   U54 : BUF_X1 port map( A => n1468, Z => n1091);
   U55 : BUF_X1 port map( A => n1468, Z => n1092);
   U56 : BUF_X1 port map( A => n1468, Z => n1093);
   U57 : BUF_X1 port map( A => n1699, Z => n605);
   U58 : BUF_X1 port map( A => n1699, Z => n606);
   U59 : BUF_X1 port map( A => n1699, Z => n607);
   U60 : BUF_X1 port map( A => n1699, Z => n1056);
   U61 : BUF_X1 port map( A => n1699, Z => n1057);
   U62 : BUF_X1 port map( A => n1470, Z => n1083);
   U63 : BUF_X1 port map( A => n1470, Z => n1084);
   U64 : BUF_X1 port map( A => n1470, Z => n1085);
   U65 : BUF_X1 port map( A => n1470, Z => n1086);
   U66 : BUF_X1 port map( A => n1470, Z => n1087);
   U67 : BUF_X1 port map( A => n1298, Z => n1148);
   U68 : BUF_X1 port map( A => n1298, Z => n1149);
   U69 : BUF_X1 port map( A => n1298, Z => n1150);
   U70 : BUF_X1 port map( A => n1298, Z => n1146);
   U71 : BUF_X1 port map( A => n1288, Z => n1158);
   U72 : BUF_X1 port map( A => n1298, Z => n1147);
   U73 : BUF_X1 port map( A => n1288, Z => n1159);
   U74 : BUF_X1 port map( A => n1288, Z => n1160);
   U75 : BUF_X1 port map( A => n1288, Z => n1161);
   U76 : BUF_X1 port map( A => n1288, Z => n1162);
   U77 : BUF_X1 port map( A => n1462, Z => n1113);
   U78 : BUF_X1 port map( A => n1462, Z => n1114);
   U79 : BUF_X1 port map( A => n1462, Z => n1115);
   U80 : BUF_X1 port map( A => n1462, Z => n1116);
   U81 : BUF_X1 port map( A => n1462, Z => n1117);
   U82 : BUF_X1 port map( A => n1396, Z => n1126);
   U83 : BUF_X1 port map( A => n1396, Z => n1127);
   U84 : BUF_X1 port map( A => n1396, Z => n1128);
   U85 : BUF_X1 port map( A => n1396, Z => n1129);
   U86 : BUF_X1 port map( A => n1396, Z => n1130);
   U87 : BUF_X1 port map( A => n1289, Z => n1152);
   U88 : BUF_X1 port map( A => n1460, Z => n1119);
   U89 : BUF_X1 port map( A => n1395, Z => n1132);
   U90 : BUF_X1 port map( A => n1300, Z => n1139);
   U91 : BUF_X1 port map( A => n1460, Z => n1120);
   U92 : BUF_X1 port map( A => n1395, Z => n1133);
   U93 : BUF_X1 port map( A => n1300, Z => n1140);
   U94 : BUF_X1 port map( A => n1464, Z => n1105);
   U95 : BUF_X1 port map( A => n1464, Z => n1104);
   U96 : BUF_X1 port map( A => n1464, Z => n1103);
   U97 : BUF_X1 port map( A => n1464, Z => n1102);
   U98 : BUF_X1 port map( A => n1464, Z => n1101);
   U99 : NAND2_X1 port map( A1 => n1391, A2 => n1121, ZN => n1462);
   U100 : NAND2_X1 port map( A1 => n1391, A2 => n1134, ZN => n1396);
   U101 : NAND2_X1 port map( A1 => n1391, A2 => n1392, ZN => n1298);
   U102 : NAND2_X1 port map( A1 => n1391, A2 => n1765, ZN => n1288);
   U103 : OAI22_X1 port map( A1 => n1125, A2 => n1477, B1 => n1307, B2 => n1118
                           , ZN => n857);
   U104 : OAI22_X1 port map( A1 => n1125, A2 => n1474, B1 => n1305, B2 => n1118
                           , ZN => n859);
   U105 : OAI22_X1 port map( A1 => n1125, A2 => n1471, B1 => n1303, B2 => n1118
                           , ZN => n861);
   U106 : OAI22_X1 port map( A1 => n1125, A2 => n1461, B1 => n1301, B2 => n1118
                           , ZN => n863);
   U107 : OAI22_X1 port map( A1 => n1121, A2 => n1687, B1 => n1297, B2 => n1113
                           , ZN => n737);
   U108 : OAI22_X1 port map( A1 => n1121, A2 => n1683, B1 => n1296, B2 => n1113
                           , ZN => n739);
   U109 : OAI22_X1 port map( A1 => n1121, A2 => n1679, B1 => n1295, B2 => n1113
                           , ZN => n741);
   U110 : OAI22_X1 port map( A1 => n1121, A2 => n1675, B1 => n1294, B2 => n1113
                           , ZN => n743);
   U111 : OAI22_X1 port map( A1 => n1121, A2 => n1671, B1 => n1293, B2 => n1113
                           , ZN => n745);
   U112 : OAI22_X1 port map( A1 => n1121, A2 => n1667, B1 => n1292, B2 => n1113
                           , ZN => n747);
   U113 : OAI22_X1 port map( A1 => n1121, A2 => n1663, B1 => n1291, B2 => n1113
                           , ZN => n749);
   U114 : OAI22_X1 port map( A1 => n1121, A2 => n1659, B1 => n1290, B2 => n1113
                           , ZN => n751);
   U115 : OAI22_X1 port map( A1 => n1121, A2 => n1655, B1 => n1390, B2 => n1113
                           , ZN => n753);
   U116 : OAI22_X1 port map( A1 => n1121, A2 => n1651, B1 => n1389, B2 => n1113
                           , ZN => n755);
   U117 : OAI22_X1 port map( A1 => n1121, A2 => n1647, B1 => n1388, B2 => n1113
                           , ZN => n757);
   U118 : OAI22_X1 port map( A1 => n1121, A2 => n1643, B1 => n1387, B2 => n1113
                           , ZN => n759);
   U119 : OAI22_X1 port map( A1 => n1122, A2 => n1639, B1 => n1386, B2 => n1114
                           , ZN => n761);
   U120 : OAI22_X1 port map( A1 => n1122, A2 => n1635, B1 => n1385, B2 => n1114
                           , ZN => n763);
   U121 : OAI22_X1 port map( A1 => n1122, A2 => n1631, B1 => n1384, B2 => n1114
                           , ZN => n765);
   U122 : OAI22_X1 port map( A1 => n1122, A2 => n1627, B1 => n1383, B2 => n1114
                           , ZN => n767);
   U123 : OAI22_X1 port map( A1 => n1122, A2 => n1623, B1 => n1382, B2 => n1114
                           , ZN => n769);
   U124 : OAI22_X1 port map( A1 => n1122, A2 => n1619, B1 => n1381, B2 => n1114
                           , ZN => n771);
   U125 : OAI22_X1 port map( A1 => n1122, A2 => n1615, B1 => n1380, B2 => n1114
                           , ZN => n773);
   U126 : OAI22_X1 port map( A1 => n1122, A2 => n1611, B1 => n1379, B2 => n1114
                           , ZN => n775);
   U127 : OAI22_X1 port map( A1 => n1122, A2 => n1607, B1 => n1378, B2 => n1114
                           , ZN => n777);
   U128 : OAI22_X1 port map( A1 => n1122, A2 => n1603, B1 => n1377, B2 => n1114
                           , ZN => n779);
   U129 : OAI22_X1 port map( A1 => n1122, A2 => n1599, B1 => n1376, B2 => n1114
                           , ZN => n781);
   U130 : OAI22_X1 port map( A1 => n1122, A2 => n1595, B1 => n1375, B2 => n1114
                           , ZN => n783);
   U131 : OAI22_X1 port map( A1 => n1122, A2 => n1591, B1 => n1374, B2 => n1115
                           , ZN => n785);
   U132 : OAI22_X1 port map( A1 => n1123, A2 => n1587, B1 => n1373, B2 => n1115
                           , ZN => n787);
   U133 : OAI22_X1 port map( A1 => n1123, A2 => n1583, B1 => n1372, B2 => n1115
                           , ZN => n789);
   U134 : OAI22_X1 port map( A1 => n1123, A2 => n1579, B1 => n1371, B2 => n1115
                           , ZN => n791);
   U135 : OAI22_X1 port map( A1 => n1123, A2 => n1575, B1 => n1370, B2 => n1115
                           , ZN => n793);
   U136 : OAI22_X1 port map( A1 => n1123, A2 => n1572, B1 => n1369, B2 => n1115
                           , ZN => n795);
   U137 : OAI22_X1 port map( A1 => n1123, A2 => n1569, B1 => n1367, B2 => n1115
                           , ZN => n797);
   U138 : OAI22_X1 port map( A1 => n1123, A2 => n1566, B1 => n1365, B2 => n1115
                           , ZN => n799);
   U139 : OAI22_X1 port map( A1 => n1123, A2 => n1563, B1 => n1363, B2 => n1115
                           , ZN => n801);
   U140 : OAI22_X1 port map( A1 => n1123, A2 => n1560, B1 => n1361, B2 => n1115
                           , ZN => n803);
   U141 : OAI22_X1 port map( A1 => n1123, A2 => n1557, B1 => n1359, B2 => n1115
                           , ZN => n805);
   U142 : OAI22_X1 port map( A1 => n1123, A2 => n1554, B1 => n1357, B2 => n1115
                           , ZN => n807);
   U143 : OAI22_X1 port map( A1 => n1123, A2 => n1551, B1 => n1355, B2 => n1116
                           , ZN => n809);
   U144 : OAI22_X1 port map( A1 => n1123, A2 => n1548, B1 => n1353, B2 => n1116
                           , ZN => n811);
   U145 : OAI22_X1 port map( A1 => n1124, A2 => n1545, B1 => n1351, B2 => n1116
                           , ZN => n813);
   U146 : OAI22_X1 port map( A1 => n1124, A2 => n1542, B1 => n1349, B2 => n1116
                           , ZN => n815);
   U147 : OAI22_X1 port map( A1 => n1124, A2 => n1539, B1 => n1347, B2 => n1116
                           , ZN => n817);
   U148 : OAI22_X1 port map( A1 => n1124, A2 => n1536, B1 => n1345, B2 => n1116
                           , ZN => n819);
   U149 : OAI22_X1 port map( A1 => n1124, A2 => n1533, B1 => n1343, B2 => n1116
                           , ZN => n821);
   U150 : OAI22_X1 port map( A1 => n1124, A2 => n1530, B1 => n1341, B2 => n1116
                           , ZN => n823);
   U151 : OAI22_X1 port map( A1 => n1124, A2 => n1527, B1 => n1339, B2 => n1116
                           , ZN => n825);
   U152 : OAI22_X1 port map( A1 => n1124, A2 => n1524, B1 => n1337, B2 => n1116
                           , ZN => n827);
   U153 : OAI22_X1 port map( A1 => n1124, A2 => n1521, B1 => n1335, B2 => n1116
                           , ZN => n829);
   U154 : OAI22_X1 port map( A1 => n1124, A2 => n1518, B1 => n1333, B2 => n1116
                           , ZN => n831);
   U155 : OAI22_X1 port map( A1 => n1124, A2 => n1515, B1 => n1331, B2 => n1117
                           , ZN => n833);
   U156 : OAI22_X1 port map( A1 => n1124, A2 => n1512, B1 => n1329, B2 => n1117
                           , ZN => n835);
   U157 : OAI22_X1 port map( A1 => n1124, A2 => n1509, B1 => n1327, B2 => n1117
                           , ZN => n837);
   U158 : OAI22_X1 port map( A1 => n1125, A2 => n1506, B1 => n1325, B2 => n1117
                           , ZN => n839);
   U159 : OAI22_X1 port map( A1 => n1125, A2 => n1503, B1 => n1323, B2 => n1117
                           , ZN => n841);
   U160 : OAI22_X1 port map( A1 => n1125, A2 => n1499, B1 => n1321, B2 => n1117
                           , ZN => n843);
   U161 : OAI22_X1 port map( A1 => n1125, A2 => n1495, B1 => n1319, B2 => n1117
                           , ZN => n845);
   U162 : OAI22_X1 port map( A1 => n1125, A2 => n1492, B1 => n1317, B2 => n1117
                           , ZN => n847);
   U163 : OAI22_X1 port map( A1 => n1125, A2 => n1489, B1 => n1315, B2 => n1117
                           , ZN => n849);
   U164 : OAI22_X1 port map( A1 => n1125, A2 => n1486, B1 => n1313, B2 => n1117
                           , ZN => n851);
   U165 : OAI22_X1 port map( A1 => n1125, A2 => n1483, B1 => n1311, B2 => n1117
                           , ZN => n853);
   U166 : OAI22_X1 port map( A1 => n1125, A2 => n1480, B1 => n1309, B2 => n1117
                           , ZN => n855);
   U167 : NAND2_X1 port map( A1 => n1391, A2 => n1158, ZN => n1289);
   U168 : AND3_X1 port map( A1 => n1076, A2 => n1169, A3 => ADD_RD1(0), ZN => 
                           n1699);
   U169 : AND3_X1 port map( A1 => n1076, A2 => n1168, A3 => ADD_RD1(1), ZN => 
                           n1697);
   U170 : AND3_X1 port map( A1 => n1106, A2 => n1167, A3 => ADD_RD2(0), ZN => 
                           n1470);
   U171 : AND3_X1 port map( A1 => n1106, A2 => n1166, A3 => ADD_RD2(1), ZN => 
                           n1466);
   U172 : AND3_X1 port map( A1 => n1168, A2 => n1169, A3 => n1076, ZN => n1698)
                           ;
   U173 : AND3_X1 port map( A1 => n1166, A2 => n1167, A3 => n1106, ZN => n1468)
                           ;
   U174 : AND2_X1 port map( A1 => RD1, A2 => n1391, ZN => n1695);
   U175 : NAND2_X1 port map( A1 => n1391, A2 => n1688, ZN => n1460);
   U176 : NAND2_X1 port map( A1 => n1391, A2 => n1458, ZN => n1395);
   U177 : NAND2_X1 port map( A1 => n1391, A2 => n1146, ZN => n1300);
   U178 : OAI221_X1 port map( B1 => n1477, B2 => n1082, C1 => n476, C2 => n1071
                           , A => n1702, ZN => n732);
   U179 : AOI222_X1 port map( A1 => n1070, A2 => n4, B1 => n1064, B2 => n1479, 
                           C1 => n1058, C2 => n68, ZN => n1702);
   U180 : OAI221_X1 port map( B1 => n1474, B2 => n1082, C1 => n477, C2 => n1071
                           , A => n1701, ZN => n733);
   U181 : AOI222_X1 port map( A1 => n1070, A2 => n3, B1 => n1064, B2 => n1476, 
                           C1 => n1058, C2 => n67, ZN => n1701);
   U182 : OAI221_X1 port map( B1 => n1471, B2 => n1082, C1 => n478, C2 => n1071
                           , A => n1700, ZN => n734);
   U183 : AOI222_X1 port map( A1 => n1070, A2 => n2, B1 => n1064, B2 => n1473, 
                           C1 => n1058, C2 => n66, ZN => n1700);
   U184 : OAI221_X1 port map( B1 => n1461, B2 => n1082, C1 => n479, C2 => n1071
                           , A => n1696, ZN => n735);
   U185 : AOI222_X1 port map( A1 => n1070, A2 => n1467, B1 => n1064, B2 => 
                           n1469, C1 => n1058, C2 => n65, ZN => n1696);
   U186 : OAI221_X1 port map( B1 => n1112, B2 => n1477, C1 => n540, C2 => n1101
                           , A => n1478, ZN => n856);
   U187 : AOI222_X1 port map( A1 => n1100, A2 => n4, B1 => n1094, B2 => n1479, 
                           C1 => n1088, C2 => n68, ZN => n1478);
   U188 : OAI221_X1 port map( B1 => n1112, B2 => n1474, C1 => n541, C2 => n1101
                           , A => n1475, ZN => n858);
   U189 : AOI222_X1 port map( A1 => n1100, A2 => n3, B1 => n1094, B2 => n1476, 
                           C1 => n1088, C2 => n67, ZN => n1475);
   U190 : OAI221_X1 port map( B1 => n1112, B2 => n1471, C1 => n542, C2 => n1101
                           , A => n1472, ZN => n860);
   U191 : AOI222_X1 port map( A1 => n1100, A2 => n2, B1 => n1094, B2 => n1473, 
                           C1 => n1088, C2 => n66, ZN => n1472);
   U192 : OAI221_X1 port map( B1 => n1461, B2 => n1112, C1 => n543, C2 => n1101
                           , A => n1465, ZN => n862);
   U193 : AOI222_X1 port map( A1 => n1100, A2 => n1467, B1 => n1094, B2 => 
                           n1469, C1 => n1088, C2 => n65, ZN => n1465);
   U194 : INV_X1 port map( A => RESET, ZN => n1391);
   U195 : OAI221_X1 port map( B1 => n1107, B2 => n1687, C1 => n480, C2 => n1106
                           , A => n1689, ZN => n736);
   U196 : AOI222_X1 port map( A1 => n1095, A2 => n64, B1 => n1089, B2 => n1690,
                           C1 => n1083, C2 => n1691, ZN => n1689);
   U197 : OAI221_X1 port map( B1 => n1107, B2 => n1683, C1 => n481, C2 => n1106
                           , A => n1684, ZN => n738);
   U198 : AOI222_X1 port map( A1 => n1095, A2 => n63, B1 => n1089, B2 => n1685,
                           C1 => n1083, C2 => n1686, ZN => n1684);
   U199 : OAI221_X1 port map( B1 => n1107, B2 => n1679, C1 => n482, C2 => n1106
                           , A => n1680, ZN => n740);
   U200 : AOI222_X1 port map( A1 => n1095, A2 => n62, B1 => n1089, B2 => n1681,
                           C1 => n1083, C2 => n1682, ZN => n1680);
   U201 : OAI221_X1 port map( B1 => n1107, B2 => n1675, C1 => n483, C2 => n1105
                           , A => n1676, ZN => n742);
   U202 : AOI222_X1 port map( A1 => n1095, A2 => n61, B1 => n1089, B2 => n1677,
                           C1 => n1083, C2 => n1678, ZN => n1676);
   U203 : OAI221_X1 port map( B1 => n1107, B2 => n1671, C1 => n484, C2 => n1106
                           , A => n1672, ZN => n744);
   U204 : AOI222_X1 port map( A1 => n1095, A2 => n60, B1 => n1089, B2 => n1673,
                           C1 => n1083, C2 => n1674, ZN => n1672);
   U205 : OAI221_X1 port map( B1 => n1107, B2 => n1667, C1 => n485, C2 => n1105
                           , A => n1668, ZN => n746);
   U206 : AOI222_X1 port map( A1 => n1095, A2 => n59, B1 => n1089, B2 => n1669,
                           C1 => n1083, C2 => n1670, ZN => n1668);
   U207 : OAI221_X1 port map( B1 => n1107, B2 => n1663, C1 => n486, C2 => n1105
                           , A => n1664, ZN => n748);
   U208 : AOI222_X1 port map( A1 => n1095, A2 => n58, B1 => n1089, B2 => n1665,
                           C1 => n1083, C2 => n1666, ZN => n1664);
   U209 : OAI221_X1 port map( B1 => n1107, B2 => n1659, C1 => n487, C2 => n1105
                           , A => n1660, ZN => n750);
   U210 : AOI222_X1 port map( A1 => n1095, A2 => n57, B1 => n1089, B2 => n1661,
                           C1 => n1083, C2 => n1662, ZN => n1660);
   U211 : OAI221_X1 port map( B1 => n1107, B2 => n1655, C1 => n488, C2 => n1105
                           , A => n1656, ZN => n752);
   U212 : AOI222_X1 port map( A1 => n1095, A2 => n56, B1 => n1089, B2 => n1657,
                           C1 => n1083, C2 => n1658, ZN => n1656);
   U213 : OAI221_X1 port map( B1 => n1107, B2 => n1651, C1 => n489, C2 => n1105
                           , A => n1652, ZN => n754);
   U214 : AOI222_X1 port map( A1 => n1095, A2 => n55, B1 => n1089, B2 => n1653,
                           C1 => n1083, C2 => n1654, ZN => n1652);
   U215 : OAI221_X1 port map( B1 => n1107, B2 => n1647, C1 => n490, C2 => n1105
                           , A => n1648, ZN => n756);
   U216 : AOI222_X1 port map( A1 => n1095, A2 => n54, B1 => n1089, B2 => n1649,
                           C1 => n1083, C2 => n1650, ZN => n1648);
   U217 : OAI221_X1 port map( B1 => n1107, B2 => n1643, C1 => n491, C2 => n1105
                           , A => n1644, ZN => n758);
   U218 : AOI222_X1 port map( A1 => n1095, A2 => n53, B1 => n1089, B2 => n1645,
                           C1 => n1083, C2 => n1646, ZN => n1644);
   U219 : OAI221_X1 port map( B1 => n1108, B2 => n1639, C1 => n492, C2 => n1105
                           , A => n1640, ZN => n760);
   U220 : AOI222_X1 port map( A1 => n1096, A2 => n52, B1 => n1090, B2 => n1641,
                           C1 => n1084, C2 => n1642, ZN => n1640);
   U221 : OAI221_X1 port map( B1 => n1108, B2 => n1635, C1 => n493, C2 => n1105
                           , A => n1636, ZN => n762);
   U222 : AOI222_X1 port map( A1 => n1096, A2 => n51, B1 => n1090, B2 => n1637,
                           C1 => n1084, C2 => n1638, ZN => n1636);
   U223 : OAI221_X1 port map( B1 => n1108, B2 => n1631, C1 => n494, C2 => n1105
                           , A => n1632, ZN => n764);
   U224 : AOI222_X1 port map( A1 => n1096, A2 => n50, B1 => n1090, B2 => n1633,
                           C1 => n1084, C2 => n1634, ZN => n1632);
   U225 : OAI221_X1 port map( B1 => n1108, B2 => n1627, C1 => n495, C2 => n1105
                           , A => n1628, ZN => n766);
   U226 : AOI222_X1 port map( A1 => n1096, A2 => n49, B1 => n1090, B2 => n1629,
                           C1 => n1084, C2 => n1630, ZN => n1628);
   U227 : OAI221_X1 port map( B1 => n1108, B2 => n1623, C1 => n496, C2 => n1104
                           , A => n1624, ZN => n768);
   U228 : AOI222_X1 port map( A1 => n1096, A2 => n48, B1 => n1090, B2 => n1625,
                           C1 => n1084, C2 => n1626, ZN => n1624);
   U229 : OAI221_X1 port map( B1 => n1108, B2 => n1619, C1 => n497, C2 => n1104
                           , A => n1620, ZN => n770);
   U230 : AOI222_X1 port map( A1 => n1096, A2 => n47, B1 => n1090, B2 => n1621,
                           C1 => n1084, C2 => n1622, ZN => n1620);
   U231 : OAI221_X1 port map( B1 => n1108, B2 => n1615, C1 => n498, C2 => n1104
                           , A => n1616, ZN => n772);
   U232 : AOI222_X1 port map( A1 => n1096, A2 => n46, B1 => n1090, B2 => n1617,
                           C1 => n1084, C2 => n1618, ZN => n1616);
   U233 : OAI221_X1 port map( B1 => n1108, B2 => n1611, C1 => n499, C2 => n1104
                           , A => n1612, ZN => n774);
   U234 : AOI222_X1 port map( A1 => n1096, A2 => n45, B1 => n1090, B2 => n1613,
                           C1 => n1084, C2 => n1614, ZN => n1612);
   U235 : OAI221_X1 port map( B1 => n1108, B2 => n1607, C1 => n500, C2 => n1104
                           , A => n1608, ZN => n776);
   U236 : AOI222_X1 port map( A1 => n1096, A2 => n44, B1 => n1090, B2 => n1609,
                           C1 => n1084, C2 => n1610, ZN => n1608);
   U237 : OAI221_X1 port map( B1 => n1108, B2 => n1603, C1 => n501, C2 => n1104
                           , A => n1604, ZN => n778);
   U238 : AOI222_X1 port map( A1 => n1096, A2 => n43, B1 => n1090, B2 => n1605,
                           C1 => n1084, C2 => n1606, ZN => n1604);
   U239 : OAI221_X1 port map( B1 => n1108, B2 => n1599, C1 => n502, C2 => n1104
                           , A => n1600, ZN => n780);
   U240 : AOI222_X1 port map( A1 => n1096, A2 => n42, B1 => n1090, B2 => n1601,
                           C1 => n1084, C2 => n1602, ZN => n1600);
   U241 : OAI221_X1 port map( B1 => n1108, B2 => n1595, C1 => n503, C2 => n1104
                           , A => n1596, ZN => n782);
   U242 : AOI222_X1 port map( A1 => n1096, A2 => n41, B1 => n1090, B2 => n1597,
                           C1 => n1084, C2 => n1598, ZN => n1596);
   U243 : OAI221_X1 port map( B1 => n1109, B2 => n1591, C1 => n504, C2 => n1104
                           , A => n1592, ZN => n784);
   U244 : AOI222_X1 port map( A1 => n1097, A2 => n40, B1 => n1091, B2 => n1593,
                           C1 => n1085, C2 => n1594, ZN => n1592);
   U245 : OAI221_X1 port map( B1 => n1109, B2 => n1587, C1 => n505, C2 => n1104
                           , A => n1588, ZN => n786);
   U246 : AOI222_X1 port map( A1 => n1097, A2 => n39, B1 => n1091, B2 => n1589,
                           C1 => n1085, C2 => n1590, ZN => n1588);
   U247 : OAI221_X1 port map( B1 => n1109, B2 => n1583, C1 => n506, C2 => n1104
                           , A => n1584, ZN => n788);
   U248 : AOI222_X1 port map( A1 => n1097, A2 => n38, B1 => n1091, B2 => n1585,
                           C1 => n1085, C2 => n1586, ZN => n1584);
   U249 : OAI221_X1 port map( B1 => n1109, B2 => n1579, C1 => n507, C2 => n1104
                           , A => n1580, ZN => n790);
   U250 : AOI222_X1 port map( A1 => n1097, A2 => n37, B1 => n1091, B2 => n1581,
                           C1 => n1085, C2 => n1582, ZN => n1580);
   U251 : OAI221_X1 port map( B1 => n1109, B2 => n1575, C1 => n508, C2 => n1103
                           , A => n1576, ZN => n792);
   U252 : AOI222_X1 port map( A1 => n1097, A2 => n36, B1 => n1091, B2 => n1577,
                           C1 => n1085, C2 => n1578, ZN => n1576);
   U253 : OAI221_X1 port map( B1 => n1109, B2 => n1572, C1 => n509, C2 => n1103
                           , A => n1573, ZN => n794);
   U254 : AOI222_X1 port map( A1 => n1097, A2 => n35, B1 => n1091, B2 => n1574,
                           C1 => n1085, C2 => n99, ZN => n1573);
   U255 : OAI221_X1 port map( B1 => n1109, B2 => n1569, C1 => n510, C2 => n1103
                           , A => n1570, ZN => n796);
   U256 : AOI222_X1 port map( A1 => n1097, A2 => n34, B1 => n1091, B2 => n1571,
                           C1 => n1085, C2 => n98, ZN => n1570);
   U257 : OAI221_X1 port map( B1 => n1109, B2 => n1566, C1 => n511, C2 => n1103
                           , A => n1567, ZN => n798);
   U258 : AOI222_X1 port map( A1 => n1097, A2 => n33, B1 => n1091, B2 => n1568,
                           C1 => n1085, C2 => n97, ZN => n1567);
   U259 : OAI221_X1 port map( B1 => n1109, B2 => n1563, C1 => n512, C2 => n1103
                           , A => n1564, ZN => n800);
   U260 : AOI222_X1 port map( A1 => n1097, A2 => n32, B1 => n1091, B2 => n1565,
                           C1 => n1085, C2 => n96, ZN => n1564);
   U261 : OAI221_X1 port map( B1 => n1109, B2 => n1560, C1 => n513, C2 => n1103
                           , A => n1561, ZN => n802);
   U262 : AOI222_X1 port map( A1 => n1097, A2 => n31, B1 => n1091, B2 => n1562,
                           C1 => n1085, C2 => n95, ZN => n1561);
   U263 : OAI221_X1 port map( B1 => n1109, B2 => n1557, C1 => n514, C2 => n1103
                           , A => n1558, ZN => n804);
   U264 : AOI222_X1 port map( A1 => n1097, A2 => n30, B1 => n1091, B2 => n1559,
                           C1 => n1085, C2 => n94, ZN => n1558);
   U265 : OAI221_X1 port map( B1 => n1109, B2 => n1554, C1 => n515, C2 => n1103
                           , A => n1555, ZN => n806);
   U266 : AOI222_X1 port map( A1 => n1097, A2 => n29, B1 => n1091, B2 => n1556,
                           C1 => n1085, C2 => n93, ZN => n1555);
   U267 : OAI221_X1 port map( B1 => n1687, B2 => n1077, C1 => n416, C2 => n1076
                           , A => n1762, ZN => n672);
   U268 : AOI222_X1 port map( A1 => n1065, A2 => n64, B1 => n1059, B2 => n1690,
                           C1 => n605, C2 => n1691, ZN => n1762);
   U269 : OAI221_X1 port map( B1 => n1683, B2 => n1077, C1 => n417, C2 => n1076
                           , A => n1761, ZN => n673);
   U270 : AOI222_X1 port map( A1 => n1065, A2 => n63, B1 => n1059, B2 => n1685,
                           C1 => n605, C2 => n1686, ZN => n1761);
   U271 : OAI221_X1 port map( B1 => n1679, B2 => n1077, C1 => n418, C2 => n1076
                           , A => n1760, ZN => n674);
   U272 : AOI222_X1 port map( A1 => n1065, A2 => n62, B1 => n1059, B2 => n1681,
                           C1 => n605, C2 => n1682, ZN => n1760);
   U273 : OAI221_X1 port map( B1 => n1675, B2 => n1077, C1 => n419, C2 => n1075
                           , A => n1759, ZN => n675);
   U274 : AOI222_X1 port map( A1 => n1065, A2 => n61, B1 => n1059, B2 => n1677,
                           C1 => n605, C2 => n1678, ZN => n1759);
   U275 : OAI221_X1 port map( B1 => n1671, B2 => n1077, C1 => n420, C2 => n1076
                           , A => n1758, ZN => n676);
   U276 : AOI222_X1 port map( A1 => n1065, A2 => n60, B1 => n1059, B2 => n1673,
                           C1 => n605, C2 => n1674, ZN => n1758);
   U277 : OAI221_X1 port map( B1 => n1667, B2 => n1077, C1 => n421, C2 => n1075
                           , A => n1757, ZN => n677);
   U278 : AOI222_X1 port map( A1 => n1065, A2 => n59, B1 => n1059, B2 => n1669,
                           C1 => n605, C2 => n1670, ZN => n1757);
   U279 : OAI221_X1 port map( B1 => n1663, B2 => n1077, C1 => n422, C2 => n1075
                           , A => n1756, ZN => n678);
   U280 : AOI222_X1 port map( A1 => n1065, A2 => n58, B1 => n1059, B2 => n1665,
                           C1 => n605, C2 => n1666, ZN => n1756);
   U281 : OAI221_X1 port map( B1 => n1659, B2 => n1077, C1 => n423, C2 => n1075
                           , A => n1755, ZN => n679);
   U282 : AOI222_X1 port map( A1 => n1065, A2 => n57, B1 => n1059, B2 => n1661,
                           C1 => n605, C2 => n1662, ZN => n1755);
   U283 : OAI221_X1 port map( B1 => n1655, B2 => n1077, C1 => n424, C2 => n1075
                           , A => n1754, ZN => n680);
   U284 : AOI222_X1 port map( A1 => n1065, A2 => n56, B1 => n1059, B2 => n1657,
                           C1 => n605, C2 => n1658, ZN => n1754);
   U285 : OAI221_X1 port map( B1 => n1651, B2 => n1077, C1 => n425, C2 => n1075
                           , A => n1753, ZN => n681);
   U286 : AOI222_X1 port map( A1 => n1065, A2 => n55, B1 => n1059, B2 => n1653,
                           C1 => n605, C2 => n1654, ZN => n1753);
   U287 : OAI221_X1 port map( B1 => n1647, B2 => n1077, C1 => n426, C2 => n1075
                           , A => n1752, ZN => n682);
   U288 : AOI222_X1 port map( A1 => n1065, A2 => n54, B1 => n1059, B2 => n1649,
                           C1 => n605, C2 => n1650, ZN => n1752);
   U289 : OAI221_X1 port map( B1 => n1643, B2 => n1077, C1 => n427, C2 => n1075
                           , A => n1751, ZN => n683);
   U290 : AOI222_X1 port map( A1 => n1065, A2 => n53, B1 => n1059, B2 => n1645,
                           C1 => n605, C2 => n1646, ZN => n1751);
   U291 : OAI221_X1 port map( B1 => n1639, B2 => n1078, C1 => n428, C2 => n1075
                           , A => n1750, ZN => n684);
   U292 : AOI222_X1 port map( A1 => n1066, A2 => n52, B1 => n1060, B2 => n1641,
                           C1 => n606, C2 => n1642, ZN => n1750);
   U293 : OAI221_X1 port map( B1 => n1635, B2 => n1078, C1 => n429, C2 => n1075
                           , A => n1749, ZN => n685);
   U294 : AOI222_X1 port map( A1 => n1066, A2 => n51, B1 => n1060, B2 => n1637,
                           C1 => n606, C2 => n1638, ZN => n1749);
   U295 : OAI221_X1 port map( B1 => n1631, B2 => n1078, C1 => n430, C2 => n1075
                           , A => n1748, ZN => n686);
   U296 : AOI222_X1 port map( A1 => n1066, A2 => n50, B1 => n1060, B2 => n1633,
                           C1 => n606, C2 => n1634, ZN => n1748);
   U297 : OAI221_X1 port map( B1 => n1627, B2 => n1078, C1 => n431, C2 => n1075
                           , A => n1747, ZN => n687);
   U298 : AOI222_X1 port map( A1 => n1066, A2 => n49, B1 => n1060, B2 => n1629,
                           C1 => n606, C2 => n1630, ZN => n1747);
   U299 : OAI221_X1 port map( B1 => n1623, B2 => n1078, C1 => n432, C2 => n1074
                           , A => n1746, ZN => n688);
   U300 : AOI222_X1 port map( A1 => n1066, A2 => n48, B1 => n1060, B2 => n1625,
                           C1 => n606, C2 => n1626, ZN => n1746);
   U301 : OAI221_X1 port map( B1 => n1619, B2 => n1078, C1 => n433, C2 => n1074
                           , A => n1745, ZN => n689);
   U302 : AOI222_X1 port map( A1 => n1066, A2 => n47, B1 => n1060, B2 => n1621,
                           C1 => n606, C2 => n1622, ZN => n1745);
   U303 : OAI221_X1 port map( B1 => n1615, B2 => n1078, C1 => n434, C2 => n1074
                           , A => n1744, ZN => n690);
   U304 : AOI222_X1 port map( A1 => n1066, A2 => n46, B1 => n1060, B2 => n1617,
                           C1 => n606, C2 => n1618, ZN => n1744);
   U305 : OAI221_X1 port map( B1 => n1611, B2 => n1078, C1 => n435, C2 => n1074
                           , A => n1743, ZN => n691);
   U306 : AOI222_X1 port map( A1 => n1066, A2 => n45, B1 => n1060, B2 => n1613,
                           C1 => n606, C2 => n1614, ZN => n1743);
   U307 : OAI221_X1 port map( B1 => n1607, B2 => n1078, C1 => n436, C2 => n1074
                           , A => n1742, ZN => n692);
   U308 : AOI222_X1 port map( A1 => n1066, A2 => n44, B1 => n1060, B2 => n1609,
                           C1 => n606, C2 => n1610, ZN => n1742);
   U309 : OAI221_X1 port map( B1 => n1603, B2 => n1078, C1 => n437, C2 => n1074
                           , A => n1741, ZN => n693);
   U310 : AOI222_X1 port map( A1 => n1066, A2 => n43, B1 => n1060, B2 => n1605,
                           C1 => n606, C2 => n1606, ZN => n1741);
   U311 : OAI221_X1 port map( B1 => n1599, B2 => n1078, C1 => n438, C2 => n1074
                           , A => n1740, ZN => n694);
   U312 : AOI222_X1 port map( A1 => n1066, A2 => n42, B1 => n1060, B2 => n1601,
                           C1 => n606, C2 => n1602, ZN => n1740);
   U313 : OAI221_X1 port map( B1 => n1595, B2 => n1078, C1 => n439, C2 => n1074
                           , A => n1739, ZN => n695);
   U314 : AOI222_X1 port map( A1 => n1066, A2 => n41, B1 => n1060, B2 => n1597,
                           C1 => n606, C2 => n1598, ZN => n1739);
   U315 : OAI221_X1 port map( B1 => n1591, B2 => n1079, C1 => n440, C2 => n1074
                           , A => n1738, ZN => n696);
   U316 : AOI222_X1 port map( A1 => n1067, A2 => n40, B1 => n1061, B2 => n1593,
                           C1 => n607, C2 => n1594, ZN => n1738);
   U317 : OAI221_X1 port map( B1 => n1587, B2 => n1079, C1 => n441, C2 => n1074
                           , A => n1737, ZN => n697);
   U318 : AOI222_X1 port map( A1 => n1067, A2 => n39, B1 => n1061, B2 => n1589,
                           C1 => n607, C2 => n1590, ZN => n1737);
   U319 : OAI221_X1 port map( B1 => n1583, B2 => n1079, C1 => n442, C2 => n1074
                           , A => n1736, ZN => n698);
   U320 : AOI222_X1 port map( A1 => n1067, A2 => n38, B1 => n1061, B2 => n1585,
                           C1 => n607, C2 => n1586, ZN => n1736);
   U321 : OAI221_X1 port map( B1 => n1579, B2 => n1079, C1 => n443, C2 => n1074
                           , A => n1735, ZN => n699);
   U322 : AOI222_X1 port map( A1 => n1067, A2 => n37, B1 => n1061, B2 => n1581,
                           C1 => n607, C2 => n1582, ZN => n1735);
   U323 : OAI221_X1 port map( B1 => n1575, B2 => n1079, C1 => n444, C2 => n1073
                           , A => n1734, ZN => n700);
   U324 : AOI222_X1 port map( A1 => n1067, A2 => n36, B1 => n1061, B2 => n1577,
                           C1 => n607, C2 => n1578, ZN => n1734);
   U325 : OAI221_X1 port map( B1 => n1572, B2 => n1079, C1 => n445, C2 => n1073
                           , A => n1733, ZN => n701);
   U326 : AOI222_X1 port map( A1 => n1067, A2 => n35, B1 => n1061, B2 => n1574,
                           C1 => n607, C2 => n99, ZN => n1733);
   U327 : OAI221_X1 port map( B1 => n1569, B2 => n1079, C1 => n446, C2 => n1073
                           , A => n1732, ZN => n702);
   U328 : AOI222_X1 port map( A1 => n1067, A2 => n34, B1 => n1061, B2 => n1571,
                           C1 => n607, C2 => n98, ZN => n1732);
   U329 : OAI221_X1 port map( B1 => n1566, B2 => n1079, C1 => n447, C2 => n1073
                           , A => n1731, ZN => n703);
   U330 : AOI222_X1 port map( A1 => n1067, A2 => n33, B1 => n1061, B2 => n1568,
                           C1 => n607, C2 => n97, ZN => n1731);
   U331 : OAI221_X1 port map( B1 => n1563, B2 => n1079, C1 => n448, C2 => n1073
                           , A => n1730, ZN => n704);
   U332 : AOI222_X1 port map( A1 => n1067, A2 => n32, B1 => n1061, B2 => n1565,
                           C1 => n607, C2 => n96, ZN => n1730);
   U333 : OAI221_X1 port map( B1 => n1560, B2 => n1079, C1 => n449, C2 => n1073
                           , A => n1729, ZN => n705);
   U334 : AOI222_X1 port map( A1 => n1067, A2 => n31, B1 => n1061, B2 => n1562,
                           C1 => n607, C2 => n95, ZN => n1729);
   U335 : OAI221_X1 port map( B1 => n1557, B2 => n1079, C1 => n450, C2 => n1073
                           , A => n1728, ZN => n706);
   U336 : AOI222_X1 port map( A1 => n1067, A2 => n30, B1 => n1061, B2 => n1559,
                           C1 => n607, C2 => n94, ZN => n1728);
   U337 : OAI221_X1 port map( B1 => n1554, B2 => n1079, C1 => n451, C2 => n1073
                           , A => n1727, ZN => n707);
   U338 : AOI222_X1 port map( A1 => n1067, A2 => n29, B1 => n1061, B2 => n1556,
                           C1 => n607, C2 => n93, ZN => n1727);
   U339 : OAI221_X1 port map( B1 => n1551, B2 => n1080, C1 => n452, C2 => n1073
                           , A => n1726, ZN => n708);
   U340 : AOI222_X1 port map( A1 => n1068, A2 => n28, B1 => n1062, B2 => n1553,
                           C1 => n1056, C2 => n92, ZN => n1726);
   U341 : OAI221_X1 port map( B1 => n1548, B2 => n1080, C1 => n453, C2 => n1073
                           , A => n1725, ZN => n709);
   U342 : AOI222_X1 port map( A1 => n1068, A2 => n27, B1 => n1062, B2 => n1550,
                           C1 => n1056, C2 => n91, ZN => n1725);
   U343 : OAI221_X1 port map( B1 => n1545, B2 => n1080, C1 => n454, C2 => n1073
                           , A => n1724, ZN => n710);
   U344 : AOI222_X1 port map( A1 => n1068, A2 => n26, B1 => n1062, B2 => n1547,
                           C1 => n1056, C2 => n90, ZN => n1724);
   U345 : OAI221_X1 port map( B1 => n1542, B2 => n1080, C1 => n455, C2 => n1072
                           , A => n1723, ZN => n711);
   U346 : AOI222_X1 port map( A1 => n1068, A2 => n25, B1 => n1062, B2 => n1544,
                           C1 => n1056, C2 => n89, ZN => n1723);
   U347 : OAI221_X1 port map( B1 => n1539, B2 => n1080, C1 => n456, C2 => n1072
                           , A => n1722, ZN => n712);
   U348 : AOI222_X1 port map( A1 => n1068, A2 => n24, B1 => n1062, B2 => n1541,
                           C1 => n1056, C2 => n88, ZN => n1722);
   U349 : OAI221_X1 port map( B1 => n1536, B2 => n1080, C1 => n457, C2 => n1072
                           , A => n1721, ZN => n713);
   U350 : AOI222_X1 port map( A1 => n1068, A2 => n23, B1 => n1062, B2 => n1538,
                           C1 => n1056, C2 => n87, ZN => n1721);
   U351 : OAI221_X1 port map( B1 => n1533, B2 => n1080, C1 => n458, C2 => n1072
                           , A => n1720, ZN => n714);
   U352 : AOI222_X1 port map( A1 => n1068, A2 => n22, B1 => n1062, B2 => n1535,
                           C1 => n1056, C2 => n86, ZN => n1720);
   U353 : OAI221_X1 port map( B1 => n1530, B2 => n1080, C1 => n459, C2 => n1072
                           , A => n1719, ZN => n715);
   U354 : AOI222_X1 port map( A1 => n1068, A2 => n21, B1 => n1062, B2 => n1532,
                           C1 => n1056, C2 => n85, ZN => n1719);
   U355 : OAI221_X1 port map( B1 => n1527, B2 => n1080, C1 => n460, C2 => n1072
                           , A => n1718, ZN => n716);
   U356 : AOI222_X1 port map( A1 => n1068, A2 => n20, B1 => n1062, B2 => n1529,
                           C1 => n1056, C2 => n84, ZN => n1718);
   U357 : OAI221_X1 port map( B1 => n1524, B2 => n1080, C1 => n461, C2 => n1072
                           , A => n1717, ZN => n717);
   U358 : AOI222_X1 port map( A1 => n1068, A2 => n19, B1 => n1062, B2 => n1526,
                           C1 => n1056, C2 => n83, ZN => n1717);
   U359 : OAI221_X1 port map( B1 => n1521, B2 => n1080, C1 => n462, C2 => n1072
                           , A => n1716, ZN => n718);
   U360 : AOI222_X1 port map( A1 => n1068, A2 => n18, B1 => n1062, B2 => n1523,
                           C1 => n1056, C2 => n82, ZN => n1716);
   U361 : OAI221_X1 port map( B1 => n1518, B2 => n1080, C1 => n463, C2 => n1072
                           , A => n1715, ZN => n719);
   U362 : AOI222_X1 port map( A1 => n1068, A2 => n17, B1 => n1062, B2 => n1520,
                           C1 => n1056, C2 => n81, ZN => n1715);
   U363 : OAI221_X1 port map( B1 => n1515, B2 => n1081, C1 => n464, C2 => n1073
                           , A => n1714, ZN => n720);
   U364 : AOI222_X1 port map( A1 => n1069, A2 => n16, B1 => n1063, B2 => n1517,
                           C1 => n1057, C2 => n80, ZN => n1714);
   U365 : OAI221_X1 port map( B1 => n1512, B2 => n1081, C1 => n465, C2 => n1072
                           , A => n1713, ZN => n721);
   U366 : AOI222_X1 port map( A1 => n1069, A2 => n15, B1 => n1063, B2 => n1514,
                           C1 => n1057, C2 => n79, ZN => n1713);
   U367 : OAI221_X1 port map( B1 => n1509, B2 => n1081, C1 => n466, C2 => n1072
                           , A => n1712, ZN => n722);
   U368 : AOI222_X1 port map( A1 => n1069, A2 => n14, B1 => n1063, B2 => n1511,
                           C1 => n1057, C2 => n78, ZN => n1712);
   U369 : OAI221_X1 port map( B1 => n1506, B2 => n1081, C1 => n467, C2 => n1072
                           , A => n1711, ZN => n723);
   U370 : AOI222_X1 port map( A1 => n1069, A2 => n13, B1 => n1063, B2 => n1508,
                           C1 => n1057, C2 => n77, ZN => n1711);
   U371 : OAI221_X1 port map( B1 => n1503, B2 => n1081, C1 => n468, C2 => n1071
                           , A => n1710, ZN => n724);
   U372 : AOI222_X1 port map( A1 => n1069, A2 => n12, B1 => n1063, B2 => n1505,
                           C1 => n1057, C2 => n76, ZN => n1710);
   U373 : OAI221_X1 port map( B1 => n1499, B2 => n1081, C1 => n469, C2 => n1071
                           , A => n1709, ZN => n725);
   U374 : AOI222_X1 port map( A1 => n1069, A2 => n1501, B1 => n1063, B2 => 
                           n1502, C1 => n1057, C2 => n75, ZN => n1709);
   U375 : OAI221_X1 port map( B1 => n1495, B2 => n1081, C1 => n470, C2 => n1071
                           , A => n1708, ZN => n726);
   U376 : AOI222_X1 port map( A1 => n1069, A2 => n1497, B1 => n1063, B2 => 
                           n1498, C1 => n1057, C2 => n74, ZN => n1708);
   U377 : OAI221_X1 port map( B1 => n1492, B2 => n1081, C1 => n471, C2 => n1071
                           , A => n1707, ZN => n727);
   U378 : AOI222_X1 port map( A1 => n1069, A2 => n9, B1 => n1063, B2 => n1494, 
                           C1 => n1057, C2 => n73, ZN => n1707);
   U379 : OAI221_X1 port map( B1 => n1489, B2 => n1081, C1 => n472, C2 => n1071
                           , A => n1706, ZN => n728);
   U380 : AOI222_X1 port map( A1 => n1069, A2 => n8, B1 => n1063, B2 => n1491, 
                           C1 => n1057, C2 => n72, ZN => n1706);
   U381 : OAI221_X1 port map( B1 => n1486, B2 => n1081, C1 => n473, C2 => n1071
                           , A => n1705, ZN => n729);
   U382 : AOI222_X1 port map( A1 => n1069, A2 => n7, B1 => n1063, B2 => n1488, 
                           C1 => n1057, C2 => n71, ZN => n1705);
   U383 : OAI221_X1 port map( B1 => n1483, B2 => n1081, C1 => n474, C2 => n1071
                           , A => n1704, ZN => n730);
   U384 : AOI222_X1 port map( A1 => n1069, A2 => n6, B1 => n1063, B2 => n1485, 
                           C1 => n1057, C2 => n70, ZN => n1704);
   U385 : OAI221_X1 port map( B1 => n1480, B2 => n1081, C1 => n475, C2 => n1071
                           , A => n1703, ZN => n731);
   U386 : AOI222_X1 port map( A1 => n1069, A2 => n5, B1 => n1063, B2 => n1482, 
                           C1 => n1057, C2 => n69, ZN => n1703);
   U387 : OAI221_X1 port map( B1 => n1110, B2 => n1551, C1 => n516, C2 => n1103
                           , A => n1552, ZN => n808);
   U388 : AOI222_X1 port map( A1 => n1098, A2 => n28, B1 => n1092, B2 => n1553,
                           C1 => n1086, C2 => n92, ZN => n1552);
   U389 : OAI221_X1 port map( B1 => n1110, B2 => n1548, C1 => n517, C2 => n1103
                           , A => n1549, ZN => n810);
   U390 : AOI222_X1 port map( A1 => n1098, A2 => n27, B1 => n1092, B2 => n1550,
                           C1 => n1086, C2 => n91, ZN => n1549);
   U391 : OAI221_X1 port map( B1 => n1110, B2 => n1545, C1 => n518, C2 => n1103
                           , A => n1546, ZN => n812);
   U392 : AOI222_X1 port map( A1 => n1098, A2 => n26, B1 => n1092, B2 => n1547,
                           C1 => n1086, C2 => n90, ZN => n1546);
   U393 : OAI221_X1 port map( B1 => n1110, B2 => n1542, C1 => n519, C2 => n1102
                           , A => n1543, ZN => n814);
   U394 : AOI222_X1 port map( A1 => n1098, A2 => n25, B1 => n1092, B2 => n1544,
                           C1 => n1086, C2 => n89, ZN => n1543);
   U395 : OAI221_X1 port map( B1 => n1110, B2 => n1539, C1 => n520, C2 => n1102
                           , A => n1540, ZN => n816);
   U396 : AOI222_X1 port map( A1 => n1098, A2 => n24, B1 => n1092, B2 => n1541,
                           C1 => n1086, C2 => n88, ZN => n1540);
   U397 : OAI221_X1 port map( B1 => n1110, B2 => n1536, C1 => n521, C2 => n1102
                           , A => n1537, ZN => n818);
   U398 : AOI222_X1 port map( A1 => n1098, A2 => n23, B1 => n1092, B2 => n1538,
                           C1 => n1086, C2 => n87, ZN => n1537);
   U399 : OAI221_X1 port map( B1 => n1110, B2 => n1533, C1 => n522, C2 => n1102
                           , A => n1534, ZN => n820);
   U400 : AOI222_X1 port map( A1 => n1098, A2 => n22, B1 => n1092, B2 => n1535,
                           C1 => n1086, C2 => n86, ZN => n1534);
   U401 : OAI221_X1 port map( B1 => n1110, B2 => n1530, C1 => n523, C2 => n1102
                           , A => n1531, ZN => n822);
   U402 : AOI222_X1 port map( A1 => n1098, A2 => n21, B1 => n1092, B2 => n1532,
                           C1 => n1086, C2 => n85, ZN => n1531);
   U403 : OAI221_X1 port map( B1 => n1110, B2 => n1527, C1 => n524, C2 => n1102
                           , A => n1528, ZN => n824);
   U404 : AOI222_X1 port map( A1 => n1098, A2 => n20, B1 => n1092, B2 => n1529,
                           C1 => n1086, C2 => n84, ZN => n1528);
   U405 : OAI221_X1 port map( B1 => n1110, B2 => n1524, C1 => n525, C2 => n1102
                           , A => n1525, ZN => n826);
   U406 : AOI222_X1 port map( A1 => n1098, A2 => n19, B1 => n1092, B2 => n1526,
                           C1 => n1086, C2 => n83, ZN => n1525);
   U407 : OAI221_X1 port map( B1 => n1110, B2 => n1521, C1 => n526, C2 => n1102
                           , A => n1522, ZN => n828);
   U408 : AOI222_X1 port map( A1 => n1098, A2 => n18, B1 => n1092, B2 => n1523,
                           C1 => n1086, C2 => n82, ZN => n1522);
   U409 : OAI221_X1 port map( B1 => n1110, B2 => n1518, C1 => n527, C2 => n1102
                           , A => n1519, ZN => n830);
   U410 : AOI222_X1 port map( A1 => n1098, A2 => n17, B1 => n1092, B2 => n1520,
                           C1 => n1086, C2 => n81, ZN => n1519);
   U411 : OAI221_X1 port map( B1 => n1111, B2 => n1515, C1 => n528, C2 => n1103
                           , A => n1516, ZN => n832);
   U412 : AOI222_X1 port map( A1 => n1099, A2 => n16, B1 => n1093, B2 => n1517,
                           C1 => n1087, C2 => n80, ZN => n1516);
   U413 : OAI221_X1 port map( B1 => n1111, B2 => n1512, C1 => n529, C2 => n1102
                           , A => n1513, ZN => n834);
   U414 : AOI222_X1 port map( A1 => n1099, A2 => n15, B1 => n1093, B2 => n1514,
                           C1 => n1087, C2 => n79, ZN => n1513);
   U415 : OAI221_X1 port map( B1 => n1111, B2 => n1509, C1 => n530, C2 => n1102
                           , A => n1510, ZN => n836);
   U416 : AOI222_X1 port map( A1 => n1099, A2 => n14, B1 => n1093, B2 => n1511,
                           C1 => n1087, C2 => n78, ZN => n1510);
   U417 : OAI221_X1 port map( B1 => n1111, B2 => n1506, C1 => n531, C2 => n1102
                           , A => n1507, ZN => n838);
   U418 : AOI222_X1 port map( A1 => n1099, A2 => n13, B1 => n1093, B2 => n1508,
                           C1 => n1087, C2 => n77, ZN => n1507);
   U419 : OAI221_X1 port map( B1 => n1111, B2 => n1503, C1 => n532, C2 => n1101
                           , A => n1504, ZN => n840);
   U420 : AOI222_X1 port map( A1 => n1099, A2 => n12, B1 => n1093, B2 => n1505,
                           C1 => n1087, C2 => n76, ZN => n1504);
   U421 : OAI221_X1 port map( B1 => n1111, B2 => n1499, C1 => n533, C2 => n1101
                           , A => n1500, ZN => n842);
   U422 : AOI222_X1 port map( A1 => n1099, A2 => n1501, B1 => n1093, B2 => 
                           n1502, C1 => n1087, C2 => n75, ZN => n1500);
   U423 : OAI221_X1 port map( B1 => n1111, B2 => n1495, C1 => n534, C2 => n1101
                           , A => n1496, ZN => n844);
   U424 : AOI222_X1 port map( A1 => n1099, A2 => n1497, B1 => n1093, B2 => 
                           n1498, C1 => n1087, C2 => n74, ZN => n1496);
   U425 : OAI221_X1 port map( B1 => n1111, B2 => n1492, C1 => n535, C2 => n1101
                           , A => n1493, ZN => n846);
   U426 : AOI222_X1 port map( A1 => n1099, A2 => n9, B1 => n1093, B2 => n1494, 
                           C1 => n1087, C2 => n73, ZN => n1493);
   U427 : OAI221_X1 port map( B1 => n1111, B2 => n1489, C1 => n536, C2 => n1101
                           , A => n1490, ZN => n848);
   U428 : AOI222_X1 port map( A1 => n1099, A2 => n8, B1 => n1093, B2 => n1491, 
                           C1 => n1087, C2 => n72, ZN => n1490);
   U429 : OAI221_X1 port map( B1 => n1111, B2 => n1486, C1 => n537, C2 => n1101
                           , A => n1487, ZN => n850);
   U430 : AOI222_X1 port map( A1 => n1099, A2 => n7, B1 => n1093, B2 => n1488, 
                           C1 => n1087, C2 => n71, ZN => n1487);
   U431 : OAI221_X1 port map( B1 => n1111, B2 => n1483, C1 => n538, C2 => n1101
                           , A => n1484, ZN => n852);
   U432 : AOI222_X1 port map( A1 => n1099, A2 => n6, B1 => n1093, B2 => n1485, 
                           C1 => n1087, C2 => n70, ZN => n1484);
   U433 : OAI221_X1 port map( B1 => n1111, B2 => n1480, C1 => n539, C2 => n1101
                           , A => n1481, ZN => n854);
   U434 : AOI222_X1 port map( A1 => n1099, A2 => n5, B1 => n1093, B2 => n1482, 
                           C1 => n1087, C2 => n69, ZN => n1481);
   U435 : OAI22_X1 port map( A1 => n608, A2 => n1162, B1 => n1156, B2 => n1297,
                           ZN => n992);
   U436 : OAI22_X1 port map( A1 => n609, A2 => n1162, B1 => n1156, B2 => n1296,
                           ZN => n993);
   U437 : OAI22_X1 port map( A1 => n610, A2 => n1162, B1 => n1156, B2 => n1295,
                           ZN => n994);
   U438 : OAI22_X1 port map( A1 => n611, A2 => n1164, B1 => n1156, B2 => n1294,
                           ZN => n995);
   U439 : OAI22_X1 port map( A1 => n628, A2 => n1159, B1 => n1153, B2 => n1378,
                           ZN => n1012);
   U440 : OAI22_X1 port map( A1 => n629, A2 => n1159, B1 => n1153, B2 => n1377,
                           ZN => n1013);
   U441 : OAI22_X1 port map( A1 => n630, A2 => n1159, B1 => n1153, B2 => n1376,
                           ZN => n1014);
   U442 : OAI22_X1 port map( A1 => n631, A2 => n1159, B1 => n1153, B2 => n1375,
                           ZN => n1015);
   U443 : OAI22_X1 port map( A1 => n632, A2 => n1159, B1 => n1153, B2 => n1374,
                           ZN => n1016);
   U444 : OAI22_X1 port map( A1 => n633, A2 => n1159, B1 => n1153, B2 => n1373,
                           ZN => n1017);
   U445 : OAI22_X1 port map( A1 => n634, A2 => n1159, B1 => n1153, B2 => n1372,
                           ZN => n1018);
   U446 : OAI22_X1 port map( A1 => n635, A2 => n1159, B1 => n1153, B2 => n1371,
                           ZN => n1019);
   U447 : OAI22_X1 port map( A1 => n636, A2 => n1159, B1 => n1153, B2 => n1370,
                           ZN => n1020);
   U448 : OAI22_X1 port map( A1 => n637, A2 => n1159, B1 => n1153, B2 => n1369,
                           ZN => n1021);
   U449 : OAI22_X1 port map( A1 => n638, A2 => n1159, B1 => n1153, B2 => n1367,
                           ZN => n1022);
   U450 : OAI22_X1 port map( A1 => n639, A2 => n1160, B1 => n1153, B2 => n1365,
                           ZN => n1023);
   U451 : OAI22_X1 port map( A1 => n640, A2 => n1160, B1 => n1154, B2 => n1363,
                           ZN => n1024);
   U452 : OAI22_X1 port map( A1 => n641, A2 => n1160, B1 => n1154, B2 => n1361,
                           ZN => n1025);
   U453 : OAI22_X1 port map( A1 => n642, A2 => n1160, B1 => n1154, B2 => n1359,
                           ZN => n1026);
   U454 : OAI22_X1 port map( A1 => n643, A2 => n1160, B1 => n1154, B2 => n1357,
                           ZN => n1027);
   U455 : OAI22_X1 port map( A1 => n644, A2 => n1160, B1 => n1154, B2 => n1355,
                           ZN => n1028);
   U456 : OAI22_X1 port map( A1 => n645, A2 => n1160, B1 => n1154, B2 => n1353,
                           ZN => n1029);
   U457 : OAI22_X1 port map( A1 => n646, A2 => n1160, B1 => n1154, B2 => n1351,
                           ZN => n1030);
   U458 : OAI22_X1 port map( A1 => n647, A2 => n1160, B1 => n1154, B2 => n1349,
                           ZN => n1031);
   U459 : OAI22_X1 port map( A1 => n648, A2 => n1160, B1 => n1154, B2 => n1347,
                           ZN => n1032);
   U460 : OAI22_X1 port map( A1 => n649, A2 => n1160, B1 => n1154, B2 => n1345,
                           ZN => n1033);
   U461 : OAI22_X1 port map( A1 => n650, A2 => n1160, B1 => n1154, B2 => n1343,
                           ZN => n1034);
   U462 : OAI22_X1 port map( A1 => n651, A2 => n1161, B1 => n1154, B2 => n1341,
                           ZN => n1035);
   U463 : OAI22_X1 port map( A1 => n652, A2 => n1161, B1 => n1155, B2 => n1339,
                           ZN => n1036);
   U464 : OAI22_X1 port map( A1 => n653, A2 => n1161, B1 => n1155, B2 => n1337,
                           ZN => n1037);
   U465 : OAI22_X1 port map( A1 => n654, A2 => n1161, B1 => n1155, B2 => n1335,
                           ZN => n1038);
   U466 : OAI22_X1 port map( A1 => n655, A2 => n1161, B1 => n1155, B2 => n1333,
                           ZN => n1039);
   U467 : OAI22_X1 port map( A1 => n656, A2 => n1161, B1 => n1155, B2 => n1331,
                           ZN => n1040);
   U468 : OAI22_X1 port map( A1 => n657, A2 => n1161, B1 => n1155, B2 => n1329,
                           ZN => n1041);
   U469 : OAI22_X1 port map( A1 => n658, A2 => n1161, B1 => n1155, B2 => n1327,
                           ZN => n1042);
   U470 : OAI22_X1 port map( A1 => n659, A2 => n1161, B1 => n1155, B2 => n1325,
                           ZN => n1043);
   U471 : OAI22_X1 port map( A1 => n660, A2 => n1161, B1 => n1155, B2 => n1323,
                           ZN => n1044);
   U472 : OAI22_X1 port map( A1 => n661, A2 => n1161, B1 => n1155, B2 => n1321,
                           ZN => n1045);
   U473 : OAI22_X1 port map( A1 => n662, A2 => n1161, B1 => n1155, B2 => n1319,
                           ZN => n1046);
   U474 : OAI22_X1 port map( A1 => n663, A2 => n1162, B1 => n1155, B2 => n1317,
                           ZN => n1047);
   U475 : OAI22_X1 port map( A1 => n664, A2 => n1162, B1 => n1156, B2 => n1315,
                           ZN => n1048);
   U476 : OAI22_X1 port map( A1 => n665, A2 => n1162, B1 => n1156, B2 => n1313,
                           ZN => n1049);
   U477 : OAI22_X1 port map( A1 => n666, A2 => n1162, B1 => n1156, B2 => n1311,
                           ZN => n1050);
   U478 : OAI22_X1 port map( A1 => n667, A2 => n1162, B1 => n1156, B2 => n1309,
                           ZN => n1051);
   U479 : OAI22_X1 port map( A1 => n668, A2 => n1162, B1 => n1156, B2 => n1307,
                           ZN => n1052);
   U480 : OAI22_X1 port map( A1 => n669, A2 => n1162, B1 => n1156, B2 => n1305,
                           ZN => n1053);
   U481 : OAI22_X1 port map( A1 => n670, A2 => n1162, B1 => n1156, B2 => n1303,
                           ZN => n1054);
   U482 : OAI22_X1 port map( A1 => n671, A2 => n1162, B1 => n1156, B2 => n1301,
                           ZN => n1055);
   U483 : OAI22_X1 port map( A1 => n612, A2 => n1164, B1 => n1157, B2 => n1293,
                           ZN => n996);
   U484 : OAI22_X1 port map( A1 => n613, A2 => n1164, B1 => n1157, B2 => n1292,
                           ZN => n997);
   U485 : OAI22_X1 port map( A1 => n614, A2 => n1164, B1 => n1157, B2 => n1291,
                           ZN => n998);
   U486 : OAI22_X1 port map( A1 => n615, A2 => n1164, B1 => n1157, B2 => n1290,
                           ZN => n999);
   U487 : OAI22_X1 port map( A1 => n1134, A2 => n1399, B1 => n1307, B2 => n1131
                           , ZN => n924);
   U488 : OAI22_X1 port map( A1 => n1134, A2 => n1398, B1 => n1305, B2 => n1131
                           , ZN => n925);
   U489 : OAI22_X1 port map( A1 => n1134, A2 => n1397, B1 => n1303, B2 => n1131
                           , ZN => n926);
   U490 : OAI22_X1 port map( A1 => n1183, A2 => n1134, B1 => n1301, B2 => n1131
                           , ZN => n927);
   U491 : OAI22_X1 port map( A1 => n1134, A2 => n1457, B1 => n1297, B2 => n1126
                           , ZN => n864);
   U492 : OAI22_X1 port map( A1 => n1138, A2 => n1456, B1 => n1296, B2 => n1126
                           , ZN => n865);
   U493 : OAI22_X1 port map( A1 => n1138, A2 => n1455, B1 => n1295, B2 => n1126
                           , ZN => n866);
   U494 : OAI22_X1 port map( A1 => n1138, A2 => n1454, B1 => n1294, B2 => n1126
                           , ZN => n867);
   U495 : OAI22_X1 port map( A1 => n1138, A2 => n1453, B1 => n1293, B2 => n1126
                           , ZN => n868);
   U496 : OAI22_X1 port map( A1 => n1138, A2 => n1452, B1 => n1292, B2 => n1126
                           , ZN => n869);
   U497 : OAI22_X1 port map( A1 => n1138, A2 => n1451, B1 => n1291, B2 => n1126
                           , ZN => n870);
   U498 : OAI22_X1 port map( A1 => n1138, A2 => n1450, B1 => n1290, B2 => n1126
                           , ZN => n871);
   U499 : OAI22_X1 port map( A1 => n1138, A2 => n1449, B1 => n1390, B2 => n1126
                           , ZN => n872);
   U500 : OAI22_X1 port map( A1 => n1138, A2 => n1448, B1 => n1389, B2 => n1126
                           , ZN => n873);
   U501 : OAI22_X1 port map( A1 => n1138, A2 => n1447, B1 => n1388, B2 => n1126
                           , ZN => n874);
   U502 : OAI22_X1 port map( A1 => n1138, A2 => n1446, B1 => n1387, B2 => n1126
                           , ZN => n875);
   U503 : OAI22_X1 port map( A1 => n1138, A2 => n1445, B1 => n1386, B2 => n1127
                           , ZN => n876);
   U504 : OAI22_X1 port map( A1 => n1138, A2 => n1444, B1 => n1385, B2 => n1127
                           , ZN => n877);
   U505 : OAI22_X1 port map( A1 => n1137, A2 => n1443, B1 => n1384, B2 => n1127
                           , ZN => n878);
   U506 : OAI22_X1 port map( A1 => n1137, A2 => n1442, B1 => n1383, B2 => n1127
                           , ZN => n879);
   U507 : OAI22_X1 port map( A1 => n1137, A2 => n1441, B1 => n1382, B2 => n1127
                           , ZN => n880);
   U508 : OAI22_X1 port map( A1 => n1137, A2 => n1440, B1 => n1381, B2 => n1127
                           , ZN => n881);
   U509 : OAI22_X1 port map( A1 => n1137, A2 => n1439, B1 => n1380, B2 => n1127
                           , ZN => n882);
   U510 : OAI22_X1 port map( A1 => n1137, A2 => n1438, B1 => n1379, B2 => n1127
                           , ZN => n883);
   U511 : OAI22_X1 port map( A1 => n1137, A2 => n1437, B1 => n1378, B2 => n1127
                           , ZN => n884);
   U512 : OAI22_X1 port map( A1 => n1137, A2 => n1436, B1 => n1377, B2 => n1127
                           , ZN => n885);
   U513 : OAI22_X1 port map( A1 => n1137, A2 => n1435, B1 => n1376, B2 => n1127
                           , ZN => n886);
   U514 : OAI22_X1 port map( A1 => n1137, A2 => n1434, B1 => n1375, B2 => n1127
                           , ZN => n887);
   U515 : OAI22_X1 port map( A1 => n1137, A2 => n1433, B1 => n1374, B2 => n1128
                           , ZN => n888);
   U516 : OAI22_X1 port map( A1 => n1137, A2 => n1432, B1 => n1373, B2 => n1128
                           , ZN => n889);
   U517 : OAI22_X1 port map( A1 => n1137, A2 => n1431, B1 => n1372, B2 => n1128
                           , ZN => n890);
   U518 : OAI22_X1 port map( A1 => n1136, A2 => n1430, B1 => n1371, B2 => n1128
                           , ZN => n891);
   U519 : OAI22_X1 port map( A1 => n1136, A2 => n1429, B1 => n1370, B2 => n1128
                           , ZN => n892);
   U520 : OAI22_X1 port map( A1 => n1136, A2 => n1428, B1 => n1369, B2 => n1128
                           , ZN => n893);
   U521 : OAI22_X1 port map( A1 => n1136, A2 => n1427, B1 => n1367, B2 => n1128
                           , ZN => n894);
   U522 : OAI22_X1 port map( A1 => n1136, A2 => n1426, B1 => n1365, B2 => n1128
                           , ZN => n895);
   U523 : OAI22_X1 port map( A1 => n1136, A2 => n1425, B1 => n1363, B2 => n1128
                           , ZN => n896);
   U524 : OAI22_X1 port map( A1 => n1136, A2 => n1424, B1 => n1361, B2 => n1128
                           , ZN => n897);
   U525 : OAI22_X1 port map( A1 => n1136, A2 => n1423, B1 => n1359, B2 => n1128
                           , ZN => n898);
   U526 : OAI22_X1 port map( A1 => n1136, A2 => n1422, B1 => n1357, B2 => n1128
                           , ZN => n899);
   U527 : OAI22_X1 port map( A1 => n1136, A2 => n1421, B1 => n1355, B2 => n1129
                           , ZN => n900);
   U528 : OAI22_X1 port map( A1 => n1136, A2 => n1420, B1 => n1353, B2 => n1129
                           , ZN => n901);
   U529 : OAI22_X1 port map( A1 => n1136, A2 => n1419, B1 => n1351, B2 => n1129
                           , ZN => n902);
   U530 : OAI22_X1 port map( A1 => n1135, A2 => n1418, B1 => n1349, B2 => n1129
                           , ZN => n903);
   U531 : OAI22_X1 port map( A1 => n1135, A2 => n1417, B1 => n1347, B2 => n1129
                           , ZN => n904);
   U532 : OAI22_X1 port map( A1 => n1135, A2 => n1416, B1 => n1345, B2 => n1129
                           , ZN => n905);
   U533 : OAI22_X1 port map( A1 => n1135, A2 => n1415, B1 => n1343, B2 => n1129
                           , ZN => n906);
   U534 : OAI22_X1 port map( A1 => n1135, A2 => n1414, B1 => n1341, B2 => n1129
                           , ZN => n907);
   U535 : OAI22_X1 port map( A1 => n1135, A2 => n1413, B1 => n1339, B2 => n1129
                           , ZN => n908);
   U536 : OAI22_X1 port map( A1 => n1135, A2 => n1412, B1 => n1337, B2 => n1129
                           , ZN => n909);
   U537 : OAI22_X1 port map( A1 => n1135, A2 => n1411, B1 => n1335, B2 => n1129
                           , ZN => n910);
   U538 : OAI22_X1 port map( A1 => n1136, A2 => n1410, B1 => n1333, B2 => n1129
                           , ZN => n911);
   U539 : OAI22_X1 port map( A1 => n1135, A2 => n1409, B1 => n1331, B2 => n1130
                           , ZN => n912);
   U540 : OAI22_X1 port map( A1 => n1135, A2 => n1408, B1 => n1329, B2 => n1130
                           , ZN => n913);
   U541 : OAI22_X1 port map( A1 => n1135, A2 => n1407, B1 => n1327, B2 => n1130
                           , ZN => n914);
   U542 : OAI22_X1 port map( A1 => n1135, A2 => n1406, B1 => n1325, B2 => n1130
                           , ZN => n915);
   U543 : OAI22_X1 port map( A1 => n1135, A2 => n1405, B1 => n1323, B2 => n1130
                           , ZN => n916);
   U544 : OAI22_X1 port map( A1 => n1163, A2 => n1134, B1 => n1321, B2 => n1130
                           , ZN => n917);
   U545 : OAI22_X1 port map( A1 => n1165, A2 => n1134, B1 => n1319, B2 => n1130
                           , ZN => n918);
   U546 : OAI22_X1 port map( A1 => n1134, A2 => n1404, B1 => n1317, B2 => n1130
                           , ZN => n919);
   U547 : OAI22_X1 port map( A1 => n1134, A2 => n1403, B1 => n1315, B2 => n1130
                           , ZN => n920);
   U548 : OAI22_X1 port map( A1 => n1134, A2 => n1402, B1 => n1313, B2 => n1130
                           , ZN => n921);
   U549 : OAI22_X1 port map( A1 => n1134, A2 => n1401, B1 => n1311, B2 => n1130
                           , ZN => n922);
   U550 : OAI22_X1 port map( A1 => n1134, A2 => n1400, B1 => n1309, B2 => n1130
                           , ZN => n923);
   U551 : OAI22_X1 port map( A1 => n544, A2 => n1146, B1 => n1297, B2 => n1141,
                           ZN => n928);
   U552 : OAI22_X1 port map( A1 => n545, A2 => n1146, B1 => n1296, B2 => n1141,
                           ZN => n929);
   U553 : OAI22_X1 port map( A1 => n546, A2 => n1146, B1 => n1295, B2 => n1141,
                           ZN => n930);
   U554 : OAI22_X1 port map( A1 => n547, A2 => n1146, B1 => n1294, B2 => n1141,
                           ZN => n931);
   U555 : OAI22_X1 port map( A1 => n548, A2 => n1146, B1 => n1293, B2 => n1141,
                           ZN => n932);
   U556 : OAI22_X1 port map( A1 => n549, A2 => n1146, B1 => n1292, B2 => n1141,
                           ZN => n933);
   U557 : OAI22_X1 port map( A1 => n550, A2 => n1146, B1 => n1291, B2 => n1141,
                           ZN => n934);
   U558 : OAI22_X1 port map( A1 => n551, A2 => n1146, B1 => n1290, B2 => n1141,
                           ZN => n935);
   U559 : OAI22_X1 port map( A1 => n552, A2 => n1146, B1 => n1141, B2 => n1390,
                           ZN => n936);
   U560 : OAI22_X1 port map( A1 => n553, A2 => n1146, B1 => n1141, B2 => n1389,
                           ZN => n937);
   U561 : OAI22_X1 port map( A1 => n554, A2 => n1146, B1 => n1141, B2 => n1388,
                           ZN => n938);
   U562 : OAI22_X1 port map( A1 => n555, A2 => n1147, B1 => n1141, B2 => n1387,
                           ZN => n939);
   U563 : OAI22_X1 port map( A1 => n556, A2 => n1147, B1 => n1142, B2 => n1386,
                           ZN => n940);
   U564 : OAI22_X1 port map( A1 => n557, A2 => n1147, B1 => n1142, B2 => n1385,
                           ZN => n941);
   U565 : OAI22_X1 port map( A1 => n558, A2 => n1147, B1 => n1142, B2 => n1384,
                           ZN => n942);
   U566 : OAI22_X1 port map( A1 => n559, A2 => n1147, B1 => n1142, B2 => n1383,
                           ZN => n943);
   U567 : OAI22_X1 port map( A1 => n560, A2 => n1147, B1 => n1142, B2 => n1382,
                           ZN => n944);
   U568 : OAI22_X1 port map( A1 => n561, A2 => n1147, B1 => n1142, B2 => n1381,
                           ZN => n945);
   U569 : OAI22_X1 port map( A1 => n562, A2 => n1147, B1 => n1142, B2 => n1380,
                           ZN => n946);
   U570 : OAI22_X1 port map( A1 => n563, A2 => n1147, B1 => n1142, B2 => n1379,
                           ZN => n947);
   U571 : OAI22_X1 port map( A1 => n564, A2 => n1147, B1 => n1142, B2 => n1378,
                           ZN => n948);
   U572 : OAI22_X1 port map( A1 => n565, A2 => n1147, B1 => n1142, B2 => n1377,
                           ZN => n949);
   U573 : OAI22_X1 port map( A1 => n566, A2 => n1147, B1 => n1142, B2 => n1376,
                           ZN => n950);
   U574 : OAI22_X1 port map( A1 => n567, A2 => n1148, B1 => n1142, B2 => n1375,
                           ZN => n951);
   U575 : OAI22_X1 port map( A1 => n568, A2 => n1148, B1 => n1142, B2 => n1374,
                           ZN => n952);
   U576 : OAI22_X1 port map( A1 => n569, A2 => n1148, B1 => n1143, B2 => n1373,
                           ZN => n953);
   U577 : OAI22_X1 port map( A1 => n570, A2 => n1148, B1 => n1143, B2 => n1372,
                           ZN => n954);
   U578 : OAI22_X1 port map( A1 => n571, A2 => n1148, B1 => n1143, B2 => n1371,
                           ZN => n955);
   U579 : OAI22_X1 port map( A1 => n572, A2 => n1148, B1 => n1143, B2 => n1370,
                           ZN => n956);
   U580 : OAI22_X1 port map( A1 => n1148, A2 => n1368, B1 => n1143, B2 => n1369
                           , ZN => n957);
   U581 : OAI22_X1 port map( A1 => n1148, A2 => n1366, B1 => n1143, B2 => n1367
                           , ZN => n958);
   U582 : OAI22_X1 port map( A1 => n1148, A2 => n1364, B1 => n1143, B2 => n1365
                           , ZN => n959);
   U583 : OAI22_X1 port map( A1 => n1148, A2 => n1362, B1 => n1143, B2 => n1363
                           , ZN => n960);
   U584 : OAI22_X1 port map( A1 => n1148, A2 => n1360, B1 => n1143, B2 => n1361
                           , ZN => n961);
   U585 : OAI22_X1 port map( A1 => n1148, A2 => n1358, B1 => n1143, B2 => n1359
                           , ZN => n962);
   U586 : OAI22_X1 port map( A1 => n1148, A2 => n1356, B1 => n1143, B2 => n1357
                           , ZN => n963);
   U587 : OAI22_X1 port map( A1 => n1149, A2 => n1354, B1 => n1143, B2 => n1355
                           , ZN => n964);
   U588 : OAI22_X1 port map( A1 => n1149, A2 => n1352, B1 => n1143, B2 => n1353
                           , ZN => n965);
   U589 : OAI22_X1 port map( A1 => n1149, A2 => n1350, B1 => n1144, B2 => n1351
                           , ZN => n966);
   U590 : OAI22_X1 port map( A1 => n1149, A2 => n1348, B1 => n1144, B2 => n1349
                           , ZN => n967);
   U591 : OAI22_X1 port map( A1 => n1149, A2 => n1346, B1 => n1144, B2 => n1347
                           , ZN => n968);
   U592 : OAI22_X1 port map( A1 => n1149, A2 => n1344, B1 => n1144, B2 => n1345
                           , ZN => n969);
   U593 : OAI22_X1 port map( A1 => n1149, A2 => n1342, B1 => n1144, B2 => n1343
                           , ZN => n970);
   U594 : OAI22_X1 port map( A1 => n1149, A2 => n1340, B1 => n1144, B2 => n1341
                           , ZN => n971);
   U595 : OAI22_X1 port map( A1 => n1149, A2 => n1338, B1 => n1144, B2 => n1339
                           , ZN => n972);
   U596 : OAI22_X1 port map( A1 => n1149, A2 => n1336, B1 => n1144, B2 => n1337
                           , ZN => n973);
   U597 : OAI22_X1 port map( A1 => n1149, A2 => n1334, B1 => n1144, B2 => n1335
                           , ZN => n974);
   U598 : OAI22_X1 port map( A1 => n1149, A2 => n1332, B1 => n1144, B2 => n1333
                           , ZN => n975);
   U599 : OAI22_X1 port map( A1 => n1149, A2 => n1330, B1 => n1144, B2 => n1331
                           , ZN => n976);
   U600 : OAI22_X1 port map( A1 => n1150, A2 => n1328, B1 => n1144, B2 => n1329
                           , ZN => n977);
   U601 : OAI22_X1 port map( A1 => n1150, A2 => n1326, B1 => n1144, B2 => n1327
                           , ZN => n978);
   U602 : OAI22_X1 port map( A1 => n1150, A2 => n1324, B1 => n1145, B2 => n1325
                           , ZN => n979);
   U603 : OAI22_X1 port map( A1 => n1150, A2 => n1322, B1 => n1145, B2 => n1323
                           , ZN => n980);
   U604 : OAI22_X1 port map( A1 => n1150, A2 => n1320, B1 => n1145, B2 => n1321
                           , ZN => n981);
   U605 : OAI22_X1 port map( A1 => n1150, A2 => n1318, B1 => n1145, B2 => n1319
                           , ZN => n982);
   U606 : OAI22_X1 port map( A1 => n1150, A2 => n1316, B1 => n1145, B2 => n1317
                           , ZN => n983);
   U607 : OAI22_X1 port map( A1 => n1150, A2 => n1314, B1 => n1145, B2 => n1315
                           , ZN => n984);
   U608 : OAI22_X1 port map( A1 => n1150, A2 => n1312, B1 => n1145, B2 => n1313
                           , ZN => n985);
   U609 : OAI22_X1 port map( A1 => n1150, A2 => n1310, B1 => n1145, B2 => n1311
                           , ZN => n986);
   U610 : OAI22_X1 port map( A1 => n1150, A2 => n1308, B1 => n1145, B2 => n1309
                           , ZN => n987);
   U611 : OAI22_X1 port map( A1 => n1150, A2 => n1306, B1 => n1145, B2 => n1307
                           , ZN => n988);
   U612 : OAI22_X1 port map( A1 => n1150, A2 => n1304, B1 => n1145, B2 => n1305
                           , ZN => n989);
   U613 : OAI22_X1 port map( A1 => n1151, A2 => n1302, B1 => n1145, B2 => n1303
                           , ZN => n990);
   U614 : OAI22_X1 port map( A1 => n1151, A2 => n1299, B1 => n1145, B2 => n1301
                           , ZN => n991);
   U615 : OAI22_X1 port map( A1 => n616, A2 => n1158, B1 => n1152, B2 => n1390,
                           ZN => n1000);
   U616 : OAI22_X1 port map( A1 => n617, A2 => n1158, B1 => n1152, B2 => n1389,
                           ZN => n1001);
   U617 : OAI22_X1 port map( A1 => n618, A2 => n1158, B1 => n1152, B2 => n1388,
                           ZN => n1002);
   U618 : OAI22_X1 port map( A1 => n619, A2 => n1158, B1 => n1152, B2 => n1387,
                           ZN => n1003);
   U619 : OAI22_X1 port map( A1 => n620, A2 => n1158, B1 => n1152, B2 => n1386,
                           ZN => n1004);
   U620 : OAI22_X1 port map( A1 => n621, A2 => n1158, B1 => n1152, B2 => n1385,
                           ZN => n1005);
   U621 : OAI22_X1 port map( A1 => n622, A2 => n1158, B1 => n1152, B2 => n1384,
                           ZN => n1006);
   U622 : OAI22_X1 port map( A1 => n623, A2 => n1158, B1 => n1152, B2 => n1383,
                           ZN => n1007);
   U623 : OAI22_X1 port map( A1 => n624, A2 => n1158, B1 => n1152, B2 => n1382,
                           ZN => n1008);
   U624 : OAI22_X1 port map( A1 => n625, A2 => n1158, B1 => n1152, B2 => n1381,
                           ZN => n1009);
   U625 : OAI22_X1 port map( A1 => n626, A2 => n1158, B1 => n1152, B2 => n1380,
                           ZN => n1010);
   U626 : OAI22_X1 port map( A1 => n627, A2 => n1159, B1 => n1152, B2 => n1379,
                           ZN => n1011);
   U627 : INV_X1 port map( A => DATAIN(8), ZN => n1390);
   U628 : INV_X1 port map( A => DATAIN(9), ZN => n1389);
   U629 : INV_X1 port map( A => DATAIN(10), ZN => n1388);
   U630 : INV_X1 port map( A => DATAIN(11), ZN => n1387);
   U631 : INV_X1 port map( A => DATAIN(12), ZN => n1386);
   U632 : INV_X1 port map( A => DATAIN(13), ZN => n1385);
   U633 : INV_X1 port map( A => DATAIN(14), ZN => n1384);
   U634 : INV_X1 port map( A => DATAIN(15), ZN => n1383);
   U635 : INV_X1 port map( A => DATAIN(16), ZN => n1382);
   U636 : INV_X1 port map( A => DATAIN(17), ZN => n1381);
   U637 : INV_X1 port map( A => DATAIN(18), ZN => n1380);
   U638 : INV_X1 port map( A => DATAIN(19), ZN => n1379);
   U639 : INV_X1 port map( A => DATAIN(20), ZN => n1378);
   U640 : INV_X1 port map( A => DATAIN(21), ZN => n1377);
   U641 : INV_X1 port map( A => DATAIN(22), ZN => n1376);
   U642 : INV_X1 port map( A => DATAIN(23), ZN => n1375);
   U643 : INV_X1 port map( A => DATAIN(24), ZN => n1374);
   U644 : INV_X1 port map( A => DATAIN(25), ZN => n1373);
   U645 : INV_X1 port map( A => DATAIN(26), ZN => n1372);
   U646 : INV_X1 port map( A => DATAIN(27), ZN => n1371);
   U647 : INV_X1 port map( A => DATAIN(28), ZN => n1370);
   U648 : INV_X1 port map( A => DATAIN(29), ZN => n1369);
   U649 : INV_X1 port map( A => DATAIN(30), ZN => n1367);
   U650 : INV_X1 port map( A => DATAIN(31), ZN => n1365);
   U651 : INV_X1 port map( A => DATAIN(32), ZN => n1363);
   U652 : INV_X1 port map( A => DATAIN(33), ZN => n1361);
   U653 : INV_X1 port map( A => DATAIN(34), ZN => n1359);
   U654 : INV_X1 port map( A => DATAIN(35), ZN => n1357);
   U655 : INV_X1 port map( A => DATAIN(36), ZN => n1355);
   U656 : INV_X1 port map( A => DATAIN(37), ZN => n1353);
   U657 : INV_X1 port map( A => DATAIN(38), ZN => n1351);
   U658 : INV_X1 port map( A => DATAIN(39), ZN => n1349);
   U659 : INV_X1 port map( A => DATAIN(40), ZN => n1347);
   U660 : INV_X1 port map( A => DATAIN(41), ZN => n1345);
   U661 : INV_X1 port map( A => DATAIN(42), ZN => n1343);
   U662 : INV_X1 port map( A => DATAIN(43), ZN => n1341);
   U663 : INV_X1 port map( A => DATAIN(44), ZN => n1339);
   U664 : INV_X1 port map( A => DATAIN(45), ZN => n1337);
   U665 : INV_X1 port map( A => DATAIN(46), ZN => n1335);
   U666 : INV_X1 port map( A => DATAIN(47), ZN => n1333);
   U667 : INV_X1 port map( A => DATAIN(48), ZN => n1331);
   U668 : INV_X1 port map( A => DATAIN(49), ZN => n1329);
   U669 : INV_X1 port map( A => DATAIN(50), ZN => n1327);
   U670 : INV_X1 port map( A => DATAIN(51), ZN => n1325);
   U671 : INV_X1 port map( A => DATAIN(52), ZN => n1323);
   U672 : INV_X1 port map( A => DATAIN(53), ZN => n1321);
   U673 : INV_X1 port map( A => DATAIN(54), ZN => n1319);
   U674 : INV_X1 port map( A => DATAIN(55), ZN => n1317);
   U675 : INV_X1 port map( A => DATAIN(56), ZN => n1315);
   U676 : INV_X1 port map( A => DATAIN(57), ZN => n1313);
   U677 : INV_X1 port map( A => DATAIN(58), ZN => n1311);
   U678 : INV_X1 port map( A => DATAIN(59), ZN => n1309);
   U679 : INV_X1 port map( A => DATAIN(60), ZN => n1307);
   U680 : INV_X1 port map( A => DATAIN(61), ZN => n1305);
   U681 : INV_X1 port map( A => DATAIN(62), ZN => n1303);
   U682 : INV_X1 port map( A => DATAIN(63), ZN => n1301);
   U683 : INV_X1 port map( A => DATAIN(0), ZN => n1297);
   U684 : INV_X1 port map( A => DATAIN(1), ZN => n1296);
   U685 : INV_X1 port map( A => DATAIN(2), ZN => n1295);
   U686 : INV_X1 port map( A => DATAIN(3), ZN => n1294);
   U687 : INV_X1 port map( A => DATAIN(4), ZN => n1293);
   U688 : INV_X1 port map( A => DATAIN(5), ZN => n1292);
   U689 : INV_X1 port map( A => DATAIN(6), ZN => n1291);
   U690 : INV_X1 port map( A => DATAIN(7), ZN => n1290);
   U691 : AND2_X1 port map( A1 => RD2, A2 => n1391, ZN => n1464);
   U692 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n1393);
   U693 : CLKBUF_X1 port map( A => n1699, Z => n1058);
   U694 : CLKBUF_X1 port map( A => n1698, Z => n1064);
   U695 : CLKBUF_X1 port map( A => n1697, Z => n1070);
   U696 : CLKBUF_X1 port map( A => n1695, Z => n1076);
   U697 : CLKBUF_X1 port map( A => n1694, Z => n1082);
   U698 : CLKBUF_X1 port map( A => n1470, Z => n1088);
   U699 : CLKBUF_X1 port map( A => n1468, Z => n1094);
   U700 : CLKBUF_X1 port map( A => n1466, Z => n1100);
   U701 : CLKBUF_X1 port map( A => n1464, Z => n1106);
   U702 : CLKBUF_X1 port map( A => n1463, Z => n1112);
   U703 : CLKBUF_X1 port map( A => n1462, Z => n1118);
   U704 : CLKBUF_X1 port map( A => n1396, Z => n1131);
   U705 : CLKBUF_X1 port map( A => n1298, Z => n1151);
   U706 : CLKBUF_X1 port map( A => n1289, Z => n1157);
   U707 : CLKBUF_X1 port map( A => n1288, Z => n1164);
   U708 : INV_X1 port map( A => ADD_RD2(0), ZN => n1166);
   U709 : INV_X1 port map( A => ADD_RD2(1), ZN => n1167);
   U710 : INV_X1 port map( A => ADD_RD1(0), ZN => n1168);
   U711 : INV_X1 port map( A => ADD_RD1(1), ZN => n1169);
   U712 : INV_X1 port map( A => ADD_WR(0), ZN => n1170);
   U713 : INV_X1 port map( A => ADD_WR(1), ZN => n1171);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_windowed_register_file_reg_size64_M4_N4_F4.all;

entity windowed_register_file_reg_size64_M4_N4_F4 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR, CALL, RETN : in std_logic;  SPILL, 
         FILL : out std_logic;  ADD_WR, ADD_RD1, ADD_RD2 : in std_logic_vector 
         (3 downto 0);  DATAIN : in std_logic_vector (63 downto 0);  OUT1, OUT2
         : out std_logic_vector (63 downto 0));

end windowed_register_file_reg_size64_M4_N4_F4;

architecture SYN_BEHAVIORAL of windowed_register_file_reg_size64_M4_N4_F4 is

   component CLKBUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XNOR2_X1
      port( A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   component register_file_reg_size64_file_size4_1
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component register_file_reg_size64_file_size4_2
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component register_file_reg_size64_file_size4_3
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component register_file_reg_size64_file_size4_4
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component register_file_reg_size64_file_size4_5
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component register_file_reg_size64_file_size4_6
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component register_file_reg_size64_file_size4_7
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component register_file_reg_size64_file_size4_8
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   component register_file_reg_size64_file_size4_0
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (1 downto 0);  DATAIN : in 
            std_logic_vector (63 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (63 downto 0));
   end component;
   
   signal global_read1, global_read2, global_write, global_out1_63_port, 
      global_out1_62_port, global_out1_61_port, global_out1_60_port, 
      global_out1_59_port, global_out1_58_port, global_out1_57_port, 
      global_out1_56_port, global_out1_55_port, global_out1_54_port, 
      global_out1_53_port, global_out1_52_port, global_out1_51_port, 
      global_out1_50_port, global_out1_49_port, global_out1_48_port, 
      global_out1_47_port, global_out1_46_port, global_out1_45_port, 
      global_out1_44_port, global_out1_43_port, global_out1_42_port, 
      global_out1_41_port, global_out1_40_port, global_out1_39_port, 
      global_out1_38_port, global_out1_37_port, global_out1_36_port, 
      global_out1_35_port, global_out1_34_port, global_out1_33_port, 
      global_out1_32_port, global_out1_31_port, global_out1_30_port, 
      global_out1_29_port, global_out1_28_port, global_out1_27_port, 
      global_out1_26_port, global_out1_25_port, global_out1_24_port, 
      global_out1_23_port, global_out1_22_port, global_out1_21_port, 
      global_out1_20_port, global_out1_19_port, global_out1_18_port, 
      global_out1_17_port, global_out1_16_port, global_out1_15_port, 
      global_out1_14_port, global_out1_13_port, global_out1_12_port, 
      global_out1_11_port, global_out1_10_port, global_out1_9_port, 
      global_out1_8_port, global_out1_7_port, global_out1_6_port, 
      global_out1_5_port, global_out1_4_port, global_out1_3_port, 
      global_out1_2_port, global_out1_1_port, global_out1_0_port, 
      io_out2_3_63_port, io_out2_3_62_port, io_out2_3_61_port, 
      io_out2_3_60_port, io_out2_3_59_port, io_out2_3_58_port, 
      io_out2_3_57_port, io_out2_3_56_port, io_out2_3_55_port, 
      io_out2_3_54_port, io_out2_3_53_port, io_out2_3_52_port, 
      io_out2_3_51_port, io_out2_3_50_port, io_out2_3_49_port, 
      io_out2_3_48_port, io_out2_3_47_port, io_out2_3_46_port, 
      io_out2_3_45_port, io_out2_3_44_port, io_out2_3_43_port, 
      io_out2_3_42_port, io_out2_3_41_port, io_out2_3_40_port, 
      io_out2_3_39_port, io_out2_3_38_port, io_out2_3_37_port, 
      io_out2_3_36_port, io_out2_3_35_port, io_out2_3_34_port, 
      io_out2_3_33_port, io_out2_3_32_port, io_out2_3_31_port, 
      io_out2_3_30_port, io_out2_3_29_port, io_out2_3_28_port, 
      io_out2_3_27_port, io_out2_3_26_port, io_out2_3_25_port, 
      io_out2_3_24_port, io_out2_3_23_port, io_out2_3_22_port, 
      io_out2_3_21_port, io_out2_3_20_port, io_out2_3_19_port, 
      io_out2_3_18_port, io_out2_3_17_port, io_out2_3_16_port, 
      io_out2_3_15_port, io_out2_3_14_port, io_out2_3_13_port, 
      io_out2_3_12_port, io_out2_3_11_port, io_out2_3_10_port, io_out2_3_9_port
      , io_out2_3_8_port, io_out2_3_7_port, io_out2_3_6_port, io_out2_3_5_port,
      io_out2_3_4_port, io_out2_3_3_port, io_out2_3_2_port, io_out2_3_1_port, 
      io_out2_3_0_port, io_out2_2_63_port, io_out2_2_62_port, io_out2_2_61_port
      , io_out2_2_60_port, io_out2_2_59_port, io_out2_2_58_port, 
      io_out2_2_57_port, io_out2_2_56_port, io_out2_2_55_port, 
      io_out2_2_54_port, io_out2_2_53_port, io_out2_2_52_port, 
      io_out2_2_51_port, io_out2_2_50_port, io_out2_2_49_port, 
      io_out2_2_48_port, io_out2_2_47_port, io_out2_2_46_port, 
      io_out2_2_45_port, io_out2_2_44_port, io_out2_2_43_port, 
      io_out2_2_42_port, io_out2_2_41_port, io_out2_2_40_port, 
      io_out2_2_39_port, io_out2_2_38_port, io_out2_2_37_port, 
      io_out2_2_36_port, io_out2_2_35_port, io_out2_2_34_port, 
      io_out2_2_33_port, io_out2_2_32_port, io_out2_2_31_port, 
      io_out2_2_30_port, io_out2_2_29_port, io_out2_2_28_port, 
      io_out2_2_27_port, io_out2_2_26_port, io_out2_2_25_port, 
      io_out2_2_24_port, io_out2_2_23_port, io_out2_2_22_port, 
      io_out2_2_21_port, io_out2_2_20_port, io_out2_2_19_port, 
      io_out2_2_18_port, io_out2_2_17_port, io_out2_2_16_port, 
      io_out2_2_15_port, io_out2_2_14_port, io_out2_2_13_port, 
      io_out2_2_12_port, io_out2_2_11_port, io_out2_2_10_port, io_out2_2_9_port
      , io_out2_2_8_port, io_out2_2_7_port, io_out2_2_6_port, io_out2_2_5_port,
      io_out2_2_4_port, io_out2_2_3_port, io_out2_2_2_port, io_out2_2_1_port, 
      io_out2_2_0_port, io_out2_1_63_port, io_out2_1_62_port, io_out2_1_61_port
      , io_out2_1_60_port, io_out2_1_59_port, io_out2_1_58_port, 
      io_out2_1_57_port, io_out2_1_56_port, io_out2_1_55_port, 
      io_out2_1_54_port, io_out2_1_53_port, io_out2_1_52_port, 
      io_out2_1_51_port, io_out2_1_50_port, io_out2_1_49_port, 
      io_out2_1_48_port, io_out2_1_47_port, io_out2_1_46_port, 
      io_out2_1_45_port, io_out2_1_44_port, io_out2_1_43_port, 
      io_out2_1_42_port, io_out2_1_41_port, io_out2_1_40_port, 
      io_out2_1_39_port, io_out2_1_38_port, io_out2_1_37_port, 
      io_out2_1_36_port, io_out2_1_35_port, io_out2_1_34_port, 
      io_out2_1_33_port, io_out2_1_32_port, io_out2_1_31_port, 
      io_out2_1_30_port, io_out2_1_29_port, io_out2_1_28_port, 
      io_out2_1_27_port, io_out2_1_26_port, io_out2_1_25_port, 
      io_out2_1_24_port, io_out2_1_23_port, io_out2_1_22_port, 
      io_out2_1_21_port, io_out2_1_20_port, io_out2_1_19_port, 
      io_out2_1_18_port, io_out2_1_17_port, io_out2_1_16_port, 
      io_out2_1_15_port, io_out2_1_14_port, io_out2_1_13_port, 
      io_out2_1_12_port, io_out2_1_11_port, io_out2_1_10_port, io_out2_1_9_port
      , io_out2_1_8_port, io_out2_1_7_port, io_out2_1_6_port, io_out2_1_5_port,
      io_out2_1_4_port, io_out2_1_3_port, io_out2_1_2_port, io_out2_1_1_port, 
      io_out2_1_0_port, io_out2_0_63_port, io_out2_0_62_port, io_out2_0_61_port
      , io_out2_0_60_port, io_out2_0_59_port, io_out2_0_58_port, 
      io_out2_0_57_port, io_out2_0_56_port, io_out2_0_55_port, 
      io_out2_0_54_port, io_out2_0_53_port, io_out2_0_52_port, 
      io_out2_0_51_port, io_out2_0_50_port, io_out2_0_49_port, 
      io_out2_0_48_port, io_out2_0_47_port, io_out2_0_46_port, 
      io_out2_0_45_port, io_out2_0_44_port, io_out2_0_43_port, 
      io_out2_0_42_port, io_out2_0_41_port, io_out2_0_40_port, 
      io_out2_0_39_port, io_out2_0_38_port, io_out2_0_37_port, 
      io_out2_0_36_port, io_out2_0_35_port, io_out2_0_34_port, 
      io_out2_0_33_port, io_out2_0_32_port, io_out2_0_31_port, 
      io_out2_0_30_port, io_out2_0_29_port, io_out2_0_28_port, 
      io_out2_0_27_port, io_out2_0_26_port, io_out2_0_25_port, 
      io_out2_0_24_port, io_out2_0_23_port, io_out2_0_22_port, 
      io_out2_0_21_port, io_out2_0_20_port, io_out2_0_19_port, 
      io_out2_0_18_port, io_out2_0_17_port, io_out2_0_16_port, 
      io_out2_0_15_port, io_out2_0_14_port, io_out2_0_13_port, 
      io_out2_0_12_port, io_out2_0_11_port, io_out2_0_10_port, io_out2_0_9_port
      , io_out2_0_8_port, io_out2_0_7_port, io_out2_0_6_port, io_out2_0_5_port,
      io_out2_0_4_port, io_out2_0_3_port, io_out2_0_2_port, io_out2_0_1_port, 
      io_out2_0_0_port, io_out1_3_63_port, io_out1_3_62_port, io_out1_3_61_port
      , io_out1_3_60_port, io_out1_3_59_port, io_out1_3_58_port, 
      io_out1_3_57_port, io_out1_3_56_port, io_out1_3_55_port, 
      io_out1_3_54_port, io_out1_3_53_port, io_out1_3_52_port, 
      io_out1_3_51_port, io_out1_3_50_port, io_out1_3_49_port, 
      io_out1_3_48_port, io_out1_3_47_port, io_out1_3_46_port, 
      io_out1_3_45_port, io_out1_3_44_port, io_out1_3_43_port, 
      io_out1_3_42_port, io_out1_3_41_port, io_out1_3_40_port, 
      io_out1_3_39_port, io_out1_3_38_port, io_out1_3_37_port, 
      io_out1_3_36_port, io_out1_3_35_port, io_out1_3_34_port, 
      io_out1_3_33_port, io_out1_3_32_port, io_out1_3_31_port, 
      io_out1_3_30_port, io_out1_3_29_port, io_out1_3_28_port, 
      io_out1_3_27_port, io_out1_3_26_port, io_out1_3_25_port, 
      io_out1_3_24_port, io_out1_3_23_port, io_out1_3_22_port, 
      io_out1_3_21_port, io_out1_3_20_port, io_out1_3_19_port, 
      io_out1_3_18_port, io_out1_3_17_port, io_out1_3_16_port, 
      io_out1_3_15_port, io_out1_3_14_port, io_out1_3_13_port, 
      io_out1_3_12_port, io_out1_3_11_port, io_out1_3_10_port, io_out1_3_9_port
      , io_out1_3_8_port, io_out1_3_7_port, io_out1_3_6_port, io_out1_3_5_port,
      io_out1_3_4_port, io_out1_3_3_port, io_out1_3_2_port, io_out1_3_1_port, 
      io_out1_3_0_port, io_out1_2_63_port, io_out1_2_62_port, io_out1_2_61_port
      , io_out1_2_60_port, io_out1_2_59_port, io_out1_2_58_port, 
      io_out1_2_57_port, io_out1_2_56_port, io_out1_2_55_port, 
      io_out1_2_54_port, io_out1_2_53_port, io_out1_2_52_port, 
      io_out1_2_51_port, io_out1_2_50_port, io_out1_2_49_port, 
      io_out1_2_48_port, io_out1_2_47_port, io_out1_2_46_port, 
      io_out1_2_45_port, io_out1_2_44_port, io_out1_2_43_port, 
      io_out1_2_42_port, io_out1_2_41_port, io_out1_2_40_port, 
      io_out1_2_39_port, io_out1_2_38_port, io_out1_2_37_port, 
      io_out1_2_36_port, io_out1_2_35_port, io_out1_2_34_port, 
      io_out1_2_33_port, io_out1_2_32_port, io_out1_2_31_port, 
      io_out1_2_30_port, io_out1_2_29_port, io_out1_2_28_port, 
      io_out1_2_27_port, io_out1_2_26_port, io_out1_2_25_port, 
      io_out1_2_24_port, io_out1_2_23_port, io_out1_2_22_port, 
      io_out1_2_21_port, io_out1_2_20_port, io_out1_2_19_port, 
      io_out1_2_18_port, io_out1_2_17_port, io_out1_2_16_port, 
      io_out1_2_15_port, io_out1_2_14_port, io_out1_2_13_port, 
      io_out1_2_12_port, io_out1_2_11_port, io_out1_2_10_port, io_out1_2_9_port
      , io_out1_2_8_port, io_out1_2_7_port, io_out1_2_6_port, io_out1_2_5_port,
      io_out1_2_4_port, io_out1_2_3_port, io_out1_2_2_port, io_out1_2_1_port, 
      io_out1_2_0_port, io_out1_1_63_port, io_out1_1_62_port, io_out1_1_61_port
      , io_out1_1_60_port, io_out1_1_59_port, io_out1_1_58_port, 
      io_out1_1_57_port, io_out1_1_56_port, io_out1_1_55_port, 
      io_out1_1_54_port, io_out1_1_53_port, io_out1_1_52_port, 
      io_out1_1_51_port, io_out1_1_50_port, io_out1_1_49_port, 
      io_out1_1_48_port, io_out1_1_47_port, io_out1_1_46_port, 
      io_out1_1_45_port, io_out1_1_44_port, io_out1_1_43_port, 
      io_out1_1_42_port, io_out1_1_41_port, io_out1_1_40_port, 
      io_out1_1_39_port, io_out1_1_38_port, io_out1_1_37_port, 
      io_out1_1_36_port, io_out1_1_35_port, io_out1_1_34_port, 
      io_out1_1_33_port, io_out1_1_32_port, io_out1_1_31_port, 
      io_out1_1_30_port, io_out1_1_29_port, io_out1_1_28_port, 
      io_out1_1_27_port, io_out1_1_26_port, io_out1_1_25_port, 
      io_out1_1_24_port, io_out1_1_23_port, io_out1_1_22_port, 
      io_out1_1_21_port, io_out1_1_20_port, io_out1_1_19_port, 
      io_out1_1_18_port, io_out1_1_17_port, io_out1_1_16_port, 
      io_out1_1_15_port, io_out1_1_14_port, io_out1_1_13_port, 
      io_out1_1_12_port, io_out1_1_11_port, io_out1_1_10_port, io_out1_1_9_port
      , io_out1_1_8_port, io_out1_1_7_port, io_out1_1_6_port, io_out1_1_5_port,
      io_out1_1_4_port, io_out1_1_3_port, io_out1_1_2_port, io_out1_1_1_port, 
      io_out1_1_0_port, io_out1_0_63_port, io_out1_0_62_port, io_out1_0_61_port
      , io_out1_0_60_port, io_out1_0_59_port, io_out1_0_58_port, 
      io_out1_0_57_port, io_out1_0_56_port, io_out1_0_55_port, 
      io_out1_0_54_port, io_out1_0_53_port, io_out1_0_52_port, 
      io_out1_0_51_port, io_out1_0_50_port, io_out1_0_49_port, 
      io_out1_0_48_port, io_out1_0_47_port, io_out1_0_46_port, 
      io_out1_0_45_port, io_out1_0_44_port, io_out1_0_43_port, 
      io_out1_0_42_port, io_out1_0_41_port, io_out1_0_40_port, 
      io_out1_0_39_port, io_out1_0_38_port, io_out1_0_37_port, 
      io_out1_0_36_port, io_out1_0_35_port, io_out1_0_34_port, 
      io_out1_0_33_port, io_out1_0_32_port, io_out1_0_31_port, 
      io_out1_0_30_port, io_out1_0_29_port, io_out1_0_28_port, 
      io_out1_0_27_port, io_out1_0_26_port, io_out1_0_25_port, 
      io_out1_0_24_port, io_out1_0_23_port, io_out1_0_22_port, 
      io_out1_0_21_port, io_out1_0_20_port, io_out1_0_19_port, 
      io_out1_0_18_port, io_out1_0_17_port, io_out1_0_16_port, 
      io_out1_0_15_port, io_out1_0_14_port, io_out1_0_13_port, 
      io_out1_0_12_port, io_out1_0_11_port, io_out1_0_10_port, io_out1_0_9_port
      , io_out1_0_8_port, io_out1_0_7_port, io_out1_0_6_port, io_out1_0_5_port,
      io_out1_0_4_port, io_out1_0_3_port, io_out1_0_2_port, io_out1_0_1_port, 
      io_out1_0_0_port, io_write_3_port, io_read2_3_port, io_read1_3_port, 
      enable_io_3_port, enable_io_2_port, enable_io_1_port, enable_io_0_port, 
      loc_out2_3_63_port, loc_out2_3_62_port, loc_out2_3_61_port, 
      loc_out2_3_60_port, loc_out2_3_59_port, loc_out2_3_58_port, 
      loc_out2_3_57_port, loc_out2_3_56_port, loc_out2_3_55_port, 
      loc_out2_3_54_port, loc_out2_3_53_port, loc_out2_3_52_port, 
      loc_out2_3_51_port, loc_out2_3_50_port, loc_out2_3_49_port, 
      loc_out2_3_48_port, loc_out2_3_47_port, loc_out2_3_46_port, 
      loc_out2_3_45_port, loc_out2_3_44_port, loc_out2_3_43_port, 
      loc_out2_3_42_port, loc_out2_3_41_port, loc_out2_3_40_port, 
      loc_out2_3_39_port, loc_out2_3_38_port, loc_out2_3_37_port, 
      loc_out2_3_36_port, loc_out2_3_35_port, loc_out2_3_34_port, 
      loc_out2_3_33_port, loc_out2_3_32_port, loc_out2_3_31_port, 
      loc_out2_3_30_port, loc_out2_3_29_port, loc_out2_3_28_port, 
      loc_out2_3_27_port, loc_out2_3_26_port, loc_out2_3_25_port, 
      loc_out2_3_24_port, loc_out2_3_23_port, loc_out2_3_22_port, 
      loc_out2_3_21_port, loc_out2_3_20_port, loc_out2_3_19_port, 
      loc_out2_3_18_port, loc_out2_3_17_port, loc_out2_3_16_port, 
      loc_out2_3_15_port, loc_out2_3_14_port, loc_out2_3_13_port, 
      loc_out2_3_12_port, loc_out2_3_11_port, loc_out2_3_10_port, 
      loc_out2_3_9_port, loc_out2_3_8_port, loc_out2_3_7_port, 
      loc_out2_3_6_port, loc_out2_3_5_port, loc_out2_3_4_port, 
      loc_out2_3_3_port, loc_out2_3_2_port, loc_out2_3_1_port, 
      loc_out2_3_0_port, loc_out2_2_63_port, loc_out2_2_62_port, 
      loc_out2_2_61_port, loc_out2_2_60_port, loc_out2_2_59_port, 
      loc_out2_2_58_port, loc_out2_2_57_port, loc_out2_2_56_port, 
      loc_out2_2_55_port, loc_out2_2_54_port, loc_out2_2_53_port, 
      loc_out2_2_52_port, loc_out2_2_51_port, loc_out2_2_50_port, 
      loc_out2_2_49_port, loc_out2_2_48_port, loc_out2_2_47_port, 
      loc_out2_2_46_port, loc_out2_2_45_port, loc_out2_2_44_port, 
      loc_out2_2_43_port, loc_out2_2_42_port, loc_out2_2_41_port, 
      loc_out2_2_40_port, loc_out2_2_39_port, loc_out2_2_38_port, 
      loc_out2_2_37_port, loc_out2_2_36_port, loc_out2_2_35_port, 
      loc_out2_2_34_port, loc_out2_2_33_port, loc_out2_2_32_port, 
      loc_out2_2_31_port, loc_out2_2_30_port, loc_out2_2_29_port, 
      loc_out2_2_28_port, loc_out2_2_27_port, loc_out2_2_26_port, 
      loc_out2_2_25_port, loc_out2_2_24_port, loc_out2_2_23_port, 
      loc_out2_2_22_port, loc_out2_2_21_port, loc_out2_2_20_port, 
      loc_out2_2_19_port, loc_out2_2_18_port, loc_out2_2_17_port, 
      loc_out2_2_16_port, loc_out2_2_15_port, loc_out2_2_14_port, 
      loc_out2_2_13_port, loc_out2_2_12_port, loc_out2_2_11_port, 
      loc_out2_2_10_port, loc_out2_2_9_port, loc_out2_2_8_port, 
      loc_out2_2_7_port, loc_out2_2_6_port, loc_out2_2_5_port, 
      loc_out2_2_4_port, loc_out2_2_3_port, loc_out2_2_2_port, 
      loc_out2_2_1_port, loc_out2_2_0_port, loc_out2_1_63_port, 
      loc_out2_1_62_port, loc_out2_1_61_port, loc_out2_1_60_port, 
      loc_out2_1_59_port, loc_out2_1_58_port, loc_out2_1_57_port, 
      loc_out2_1_56_port, loc_out2_1_55_port, loc_out2_1_54_port, 
      loc_out2_1_53_port, loc_out2_1_52_port, loc_out2_1_51_port, 
      loc_out2_1_50_port, loc_out2_1_49_port, loc_out2_1_48_port, 
      loc_out2_1_47_port, loc_out2_1_46_port, loc_out2_1_45_port, 
      loc_out2_1_44_port, loc_out2_1_43_port, loc_out2_1_42_port, 
      loc_out2_1_41_port, loc_out2_1_40_port, loc_out2_1_39_port, 
      loc_out2_1_38_port, loc_out2_1_37_port, loc_out2_1_36_port, 
      loc_out2_1_35_port, loc_out2_1_34_port, loc_out2_1_33_port, 
      loc_out2_1_32_port, loc_out2_1_31_port, loc_out2_1_30_port, 
      loc_out2_1_29_port, loc_out2_1_28_port, loc_out2_1_27_port, 
      loc_out2_1_26_port, loc_out2_1_25_port, loc_out2_1_24_port, 
      loc_out2_1_23_port, loc_out2_1_22_port, loc_out2_1_21_port, 
      loc_out2_1_20_port, loc_out2_1_19_port, loc_out2_1_18_port, 
      loc_out2_1_17_port, loc_out2_1_16_port, loc_out2_1_15_port, 
      loc_out2_1_14_port, loc_out2_1_13_port, loc_out2_1_12_port, 
      loc_out2_1_11_port, loc_out2_1_10_port, loc_out2_1_9_port, 
      loc_out2_1_8_port, loc_out2_1_7_port, loc_out2_1_6_port, 
      loc_out2_1_5_port, loc_out2_1_4_port, loc_out2_1_3_port, 
      loc_out2_1_2_port, loc_out2_1_1_port, loc_out2_1_0_port, 
      loc_out2_0_63_port, loc_out2_0_62_port, loc_out2_0_61_port, 
      loc_out2_0_60_port, loc_out2_0_59_port, loc_out2_0_58_port, 
      loc_out2_0_57_port, loc_out2_0_56_port, loc_out2_0_55_port, 
      loc_out2_0_54_port, loc_out2_0_53_port, loc_out2_0_52_port, 
      loc_out2_0_51_port, loc_out2_0_50_port, loc_out2_0_49_port, 
      loc_out2_0_48_port, loc_out2_0_47_port, loc_out2_0_46_port, 
      loc_out2_0_45_port, loc_out2_0_44_port, loc_out2_0_43_port, 
      loc_out2_0_42_port, loc_out2_0_41_port, loc_out2_0_40_port, 
      loc_out2_0_39_port, loc_out2_0_38_port, loc_out2_0_37_port, 
      loc_out2_0_36_port, loc_out2_0_35_port, loc_out2_0_34_port, 
      loc_out2_0_33_port, loc_out2_0_32_port, loc_out2_0_31_port, 
      loc_out2_0_30_port, loc_out2_0_29_port, loc_out2_0_28_port, 
      loc_out2_0_27_port, loc_out2_0_26_port, loc_out2_0_25_port, 
      loc_out2_0_24_port, loc_out2_0_23_port, loc_out2_0_22_port, 
      loc_out2_0_21_port, loc_out2_0_20_port, loc_out2_0_19_port, 
      loc_out2_0_18_port, loc_out2_0_17_port, loc_out2_0_16_port, 
      loc_out2_0_15_port, loc_out2_0_14_port, loc_out2_0_13_port, 
      loc_out2_0_12_port, loc_out2_0_11_port, loc_out2_0_10_port, 
      loc_out2_0_9_port, loc_out2_0_8_port, loc_out2_0_7_port, 
      loc_out2_0_6_port, loc_out2_0_5_port, loc_out2_0_4_port, 
      loc_out2_0_3_port, loc_out2_0_2_port, loc_out2_0_1_port, 
      loc_out2_0_0_port, loc_out1_3_63_port, loc_out1_3_62_port, 
      loc_out1_3_61_port, loc_out1_3_60_port, loc_out1_3_59_port, 
      loc_out1_3_58_port, loc_out1_3_57_port, loc_out1_3_56_port, 
      loc_out1_3_55_port, loc_out1_3_54_port, loc_out1_3_53_port, 
      loc_out1_3_52_port, loc_out1_3_51_port, loc_out1_3_50_port, 
      loc_out1_3_49_port, loc_out1_3_48_port, loc_out1_3_47_port, 
      loc_out1_3_46_port, loc_out1_3_45_port, loc_out1_3_44_port, 
      loc_out1_3_43_port, loc_out1_3_42_port, loc_out1_3_41_port, 
      loc_out1_3_40_port, loc_out1_3_39_port, loc_out1_3_38_port, 
      loc_out1_3_37_port, loc_out1_3_36_port, loc_out1_3_35_port, 
      loc_out1_3_34_port, loc_out1_3_33_port, loc_out1_3_32_port, 
      loc_out1_3_31_port, loc_out1_3_30_port, loc_out1_3_29_port, 
      loc_out1_3_28_port, loc_out1_3_27_port, loc_out1_3_26_port, 
      loc_out1_3_25_port, loc_out1_3_24_port, loc_out1_3_23_port, 
      loc_out1_3_22_port, loc_out1_3_21_port, loc_out1_3_20_port, 
      loc_out1_3_19_port, loc_out1_3_18_port, loc_out1_3_17_port, 
      loc_out1_3_16_port, loc_out1_3_15_port, loc_out1_3_14_port, 
      loc_out1_3_13_port, loc_out1_3_12_port, loc_out1_3_11_port, 
      loc_out1_3_10_port, loc_out1_3_9_port, loc_out1_3_8_port, 
      loc_out1_3_7_port, loc_out1_3_6_port, loc_out1_3_5_port, 
      loc_out1_3_4_port, loc_out1_3_3_port, loc_out1_3_2_port, 
      loc_out1_3_1_port, loc_out1_3_0_port, loc_out1_2_63_port, 
      loc_out1_2_62_port, loc_out1_2_61_port, loc_out1_2_60_port, 
      loc_out1_2_59_port, loc_out1_2_58_port, loc_out1_2_57_port, 
      loc_out1_2_56_port, loc_out1_2_55_port, loc_out1_2_54_port, 
      loc_out1_2_53_port, loc_out1_2_52_port, loc_out1_2_51_port, 
      loc_out1_2_50_port, loc_out1_2_49_port, loc_out1_2_48_port, 
      loc_out1_2_47_port, loc_out1_2_46_port, loc_out1_2_45_port, 
      loc_out1_2_44_port, loc_out1_2_43_port, loc_out1_2_42_port, 
      loc_out1_2_41_port, loc_out1_2_40_port, loc_out1_2_39_port, 
      loc_out1_2_38_port, loc_out1_2_37_port, loc_out1_2_36_port, 
      loc_out1_2_35_port, loc_out1_2_34_port, loc_out1_2_33_port, 
      loc_out1_2_32_port, loc_out1_2_31_port, loc_out1_2_30_port, 
      loc_out1_2_29_port, loc_out1_2_28_port, loc_out1_2_27_port, 
      loc_out1_2_26_port, loc_out1_2_25_port, loc_out1_2_24_port, 
      loc_out1_2_23_port, loc_out1_2_22_port, loc_out1_2_21_port, 
      loc_out1_2_20_port, loc_out1_2_19_port, loc_out1_2_18_port, 
      loc_out1_2_17_port, loc_out1_2_16_port, loc_out1_2_15_port, 
      loc_out1_2_14_port, loc_out1_2_13_port, loc_out1_2_12_port, 
      loc_out1_2_11_port, loc_out1_2_10_port, loc_out1_2_9_port, 
      loc_out1_2_8_port, loc_out1_2_7_port, loc_out1_2_6_port, 
      loc_out1_2_5_port, loc_out1_2_4_port, loc_out1_2_3_port, 
      loc_out1_2_2_port, loc_out1_2_1_port, loc_out1_2_0_port, 
      loc_out1_1_63_port, loc_out1_1_62_port, loc_out1_1_61_port, 
      loc_out1_1_60_port, loc_out1_1_59_port, loc_out1_1_58_port, 
      loc_out1_1_57_port, loc_out1_1_56_port, loc_out1_1_55_port, 
      loc_out1_1_54_port, loc_out1_1_53_port, loc_out1_1_52_port, 
      loc_out1_1_51_port, loc_out1_1_50_port, loc_out1_1_49_port, 
      loc_out1_1_48_port, loc_out1_1_47_port, loc_out1_1_46_port, 
      loc_out1_1_45_port, loc_out1_1_44_port, loc_out1_1_43_port, 
      loc_out1_1_42_port, loc_out1_1_41_port, loc_out1_1_40_port, 
      loc_out1_1_39_port, loc_out1_1_38_port, loc_out1_1_37_port, 
      loc_out1_1_36_port, loc_out1_1_35_port, loc_out1_1_34_port, 
      loc_out1_1_33_port, loc_out1_1_32_port, loc_out1_1_31_port, 
      loc_out1_1_30_port, loc_out1_1_29_port, loc_out1_1_28_port, 
      loc_out1_1_27_port, loc_out1_1_26_port, loc_out1_1_25_port, 
      loc_out1_1_24_port, loc_out1_1_23_port, loc_out1_1_22_port, 
      loc_out1_1_21_port, loc_out1_1_20_port, loc_out1_1_19_port, 
      loc_out1_1_18_port, loc_out1_1_17_port, loc_out1_1_16_port, 
      loc_out1_1_15_port, loc_out1_1_14_port, loc_out1_1_13_port, 
      loc_out1_1_12_port, loc_out1_1_11_port, loc_out1_1_10_port, 
      loc_out1_1_9_port, loc_out1_1_8_port, loc_out1_1_7_port, 
      loc_out1_1_6_port, loc_out1_1_5_port, loc_out1_1_4_port, 
      loc_out1_1_3_port, loc_out1_1_2_port, loc_out1_1_1_port, 
      loc_out1_1_0_port, loc_out1_0_63_port, loc_out1_0_62_port, 
      loc_out1_0_61_port, loc_out1_0_60_port, loc_out1_0_59_port, 
      loc_out1_0_58_port, loc_out1_0_57_port, loc_out1_0_56_port, 
      loc_out1_0_55_port, loc_out1_0_54_port, loc_out1_0_53_port, 
      loc_out1_0_52_port, loc_out1_0_51_port, loc_out1_0_50_port, 
      loc_out1_0_49_port, loc_out1_0_48_port, loc_out1_0_47_port, 
      loc_out1_0_46_port, loc_out1_0_45_port, loc_out1_0_44_port, 
      loc_out1_0_43_port, loc_out1_0_42_port, loc_out1_0_41_port, 
      loc_out1_0_40_port, loc_out1_0_39_port, loc_out1_0_38_port, 
      loc_out1_0_37_port, loc_out1_0_36_port, loc_out1_0_35_port, 
      loc_out1_0_34_port, loc_out1_0_33_port, loc_out1_0_32_port, 
      loc_out1_0_31_port, loc_out1_0_30_port, loc_out1_0_29_port, 
      loc_out1_0_28_port, loc_out1_0_27_port, loc_out1_0_26_port, 
      loc_out1_0_25_port, loc_out1_0_24_port, loc_out1_0_23_port, 
      loc_out1_0_22_port, loc_out1_0_21_port, loc_out1_0_20_port, 
      loc_out1_0_19_port, loc_out1_0_18_port, loc_out1_0_17_port, 
      loc_out1_0_16_port, loc_out1_0_15_port, loc_out1_0_14_port, 
      loc_out1_0_13_port, loc_out1_0_12_port, loc_out1_0_11_port, 
      loc_out1_0_10_port, loc_out1_0_9_port, loc_out1_0_8_port, 
      loc_out1_0_7_port, loc_out1_0_6_port, loc_out1_0_5_port, 
      loc_out1_0_4_port, loc_out1_0_3_port, loc_out1_0_2_port, 
      loc_out1_0_1_port, loc_out1_0_0_port, loc_write_3_port, loc_read2_3_port,
      loc_read1_3_port, enable_loc_3_port, enable_loc_2_port, enable_loc_1_port
      , enable_loc_0_port, N1132, N1133, N1134, N1135, N1136, N1137, N1138, 
      N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148, 
      N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158, 
      N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168, 
      N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177, N1178, 
      N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187, N1188, 
      N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1235, net320, net321, 
      net322, net323, net324, net325, net326, net327, net328, net329, net330, 
      net331, net332, net333, net334, net335, net336, net337, net338, net339, 
      net340, net341, net342, net343, net344, net345, net346, net347, net348, 
      net349, net350, net351, net352, net353, net354, net355, net356, net357, 
      net358, net359, net360, net361, net362, net363, net364, net365, net366, 
      net367, net368, net369, net370, net371, net372, net373, net374, net375, 
      net376, net377, net378, net379, net380, net381, net382, net383, n1035, 
      n1036, n1038, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, 
      n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, 
      n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, 
      n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, 
      n2140, n2141, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, 
      n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, 
      n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, 
      n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, 
      n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, 
      n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, 
      n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, 
      n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, 
      n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, 
      n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, 
      n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, 
      n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, 
      n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, 
      n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, 
      n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, 
      n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, 
      n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, 
      n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, 
      n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, 
      n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, 
      n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, 
      n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, 
      n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, 
      n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, 
      n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, 
      n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, 
      n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, 
      n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, 
      n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, 
      n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, 
      n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, 
      n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, 
      n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, 
      n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, 
      n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, 
      n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, 
      n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, 
      n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, 
      n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, 
      n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, 
      n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, 
      n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, 
      n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, 
      n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, 
      n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, 
      n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, 
      n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, 
      n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, 
      n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, 
      n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, 
      n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, 
      n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, 
      n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, 
      n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, 
      n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, 
      n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, 
      n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, 
      n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, 
      n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, 
      n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, 
      n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, 
      n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, 
      n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, 
      n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, 
      n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, 
      n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, 
      n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, 
      n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, 
      n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, 
      n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, 
      n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, 
      n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, 
      n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, 
      n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, 
      n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, 
      n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, 
      n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, 
      n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, 
      n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, 
      n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, 
      n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, 
      n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, 
      n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, 
      n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, 
      n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, 
      n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, 
      n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, 
      n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, 
      n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, 
      n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, 
      n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, 
      n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, 
      n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, 
      n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080 : 
      std_logic;

begin
   
   global_rf : register_file_reg_size64_file_size4_0 port map( CLK => CLK, 
                           RESET => RESET, ENABLE => ENABLE, RD1 => 
                           global_read1, RD2 => global_read2, WR => 
                           global_write, ADD_WR(1) => ADD_WR(1), ADD_WR(0) => 
                           ADD_WR(0), ADD_RD1(1) => ADD_RD1(1), ADD_RD1(0) => 
                           ADD_RD1(0), ADD_RD2(1) => ADD_RD2(1), ADD_RD2(0) => 
                           ADD_RD2(0), DATAIN(63) => DATAIN(63), DATAIN(62) => 
                           DATAIN(62), DATAIN(61) => DATAIN(61), DATAIN(60) => 
                           DATAIN(60), DATAIN(59) => DATAIN(59), DATAIN(58) => 
                           DATAIN(58), DATAIN(57) => DATAIN(57), DATAIN(56) => 
                           DATAIN(56), DATAIN(55) => DATAIN(55), DATAIN(54) => 
                           DATAIN(54), DATAIN(53) => DATAIN(53), DATAIN(52) => 
                           DATAIN(52), DATAIN(51) => DATAIN(51), DATAIN(50) => 
                           DATAIN(50), DATAIN(49) => DATAIN(49), DATAIN(48) => 
                           DATAIN(48), DATAIN(47) => DATAIN(47), DATAIN(46) => 
                           DATAIN(46), DATAIN(45) => DATAIN(45), DATAIN(44) => 
                           DATAIN(44), DATAIN(43) => DATAIN(43), DATAIN(42) => 
                           DATAIN(42), DATAIN(41) => DATAIN(41), DATAIN(40) => 
                           DATAIN(40), DATAIN(39) => DATAIN(39), DATAIN(38) => 
                           DATAIN(38), DATAIN(37) => DATAIN(37), DATAIN(36) => 
                           DATAIN(36), DATAIN(35) => DATAIN(35), DATAIN(34) => 
                           DATAIN(34), DATAIN(33) => DATAIN(33), DATAIN(32) => 
                           DATAIN(32), DATAIN(31) => DATAIN(31), DATAIN(30) => 
                           DATAIN(30), DATAIN(29) => DATAIN(29), DATAIN(28) => 
                           DATAIN(28), DATAIN(27) => DATAIN(27), DATAIN(26) => 
                           DATAIN(26), DATAIN(25) => DATAIN(25), DATAIN(24) => 
                           DATAIN(24), DATAIN(23) => DATAIN(23), DATAIN(22) => 
                           DATAIN(22), DATAIN(21) => DATAIN(21), DATAIN(20) => 
                           DATAIN(20), DATAIN(19) => DATAIN(19), DATAIN(18) => 
                           DATAIN(18), DATAIN(17) => DATAIN(17), DATAIN(16) => 
                           DATAIN(16), DATAIN(15) => DATAIN(15), DATAIN(14) => 
                           DATAIN(14), DATAIN(13) => DATAIN(13), DATAIN(12) => 
                           DATAIN(12), DATAIN(11) => DATAIN(11), DATAIN(10) => 
                           DATAIN(10), DATAIN(9) => DATAIN(9), DATAIN(8) => 
                           DATAIN(8), DATAIN(7) => DATAIN(7), DATAIN(6) => 
                           DATAIN(6), DATAIN(5) => DATAIN(5), DATAIN(4) => 
                           DATAIN(4), DATAIN(3) => DATAIN(3), DATAIN(2) => 
                           DATAIN(2), DATAIN(1) => DATAIN(1), DATAIN(0) => 
                           DATAIN(0), OUT1(63) => global_out1_63_port, OUT1(62)
                           => global_out1_62_port, OUT1(61) => 
                           global_out1_61_port, OUT1(60) => global_out1_60_port
                           , OUT1(59) => global_out1_59_port, OUT1(58) => 
                           global_out1_58_port, OUT1(57) => global_out1_57_port
                           , OUT1(56) => global_out1_56_port, OUT1(55) => 
                           global_out1_55_port, OUT1(54) => global_out1_54_port
                           , OUT1(53) => global_out1_53_port, OUT1(52) => 
                           global_out1_52_port, OUT1(51) => global_out1_51_port
                           , OUT1(50) => global_out1_50_port, OUT1(49) => 
                           global_out1_49_port, OUT1(48) => global_out1_48_port
                           , OUT1(47) => global_out1_47_port, OUT1(46) => 
                           global_out1_46_port, OUT1(45) => global_out1_45_port
                           , OUT1(44) => global_out1_44_port, OUT1(43) => 
                           global_out1_43_port, OUT1(42) => global_out1_42_port
                           , OUT1(41) => global_out1_41_port, OUT1(40) => 
                           global_out1_40_port, OUT1(39) => global_out1_39_port
                           , OUT1(38) => global_out1_38_port, OUT1(37) => 
                           global_out1_37_port, OUT1(36) => global_out1_36_port
                           , OUT1(35) => global_out1_35_port, OUT1(34) => 
                           global_out1_34_port, OUT1(33) => global_out1_33_port
                           , OUT1(32) => global_out1_32_port, OUT1(31) => 
                           global_out1_31_port, OUT1(30) => global_out1_30_port
                           , OUT1(29) => global_out1_29_port, OUT1(28) => 
                           global_out1_28_port, OUT1(27) => global_out1_27_port
                           , OUT1(26) => global_out1_26_port, OUT1(25) => 
                           global_out1_25_port, OUT1(24) => global_out1_24_port
                           , OUT1(23) => global_out1_23_port, OUT1(22) => 
                           global_out1_22_port, OUT1(21) => global_out1_21_port
                           , OUT1(20) => global_out1_20_port, OUT1(19) => 
                           global_out1_19_port, OUT1(18) => global_out1_18_port
                           , OUT1(17) => global_out1_17_port, OUT1(16) => 
                           global_out1_16_port, OUT1(15) => global_out1_15_port
                           , OUT1(14) => global_out1_14_port, OUT1(13) => 
                           global_out1_13_port, OUT1(12) => global_out1_12_port
                           , OUT1(11) => global_out1_11_port, OUT1(10) => 
                           global_out1_10_port, OUT1(9) => global_out1_9_port, 
                           OUT1(8) => global_out1_8_port, OUT1(7) => 
                           global_out1_7_port, OUT1(6) => global_out1_6_port, 
                           OUT1(5) => global_out1_5_port, OUT1(4) => 
                           global_out1_4_port, OUT1(3) => global_out1_3_port, 
                           OUT1(2) => global_out1_2_port, OUT1(1) => 
                           global_out1_1_port, OUT1(0) => global_out1_0_port, 
                           OUT2(63) => net320, OUT2(62) => net321, OUT2(61) => 
                           net322, OUT2(60) => net323, OUT2(59) => net324, 
                           OUT2(58) => net325, OUT2(57) => net326, OUT2(56) => 
                           net327, OUT2(55) => net328, OUT2(54) => net329, 
                           OUT2(53) => net330, OUT2(52) => net331, OUT2(51) => 
                           net332, OUT2(50) => net333, OUT2(49) => net334, 
                           OUT2(48) => net335, OUT2(47) => net336, OUT2(46) => 
                           net337, OUT2(45) => net338, OUT2(44) => net339, 
                           OUT2(43) => net340, OUT2(42) => net341, OUT2(41) => 
                           net342, OUT2(40) => net343, OUT2(39) => net344, 
                           OUT2(38) => net345, OUT2(37) => net346, OUT2(36) => 
                           net347, OUT2(35) => net348, OUT2(34) => net349, 
                           OUT2(33) => net350, OUT2(32) => net351, OUT2(31) => 
                           net352, OUT2(30) => net353, OUT2(29) => net354, 
                           OUT2(28) => net355, OUT2(27) => net356, OUT2(26) => 
                           net357, OUT2(25) => net358, OUT2(24) => net359, 
                           OUT2(23) => net360, OUT2(22) => net361, OUT2(21) => 
                           net362, OUT2(20) => net363, OUT2(19) => net364, 
                           OUT2(18) => net365, OUT2(17) => net366, OUT2(16) => 
                           net367, OUT2(15) => net368, OUT2(14) => net369, 
                           OUT2(13) => net370, OUT2(12) => net371, OUT2(11) => 
                           net372, OUT2(10) => net373, OUT2(9) => net374, 
                           OUT2(8) => net375, OUT2(7) => net376, OUT2(6) => 
                           net377, OUT2(5) => net378, OUT2(4) => net379, 
                           OUT2(3) => net380, OUT2(2) => net381, OUT2(1) => 
                           net382, OUT2(0) => net383);
   io_rf_0 : register_file_reg_size64_file_size4_8 port map( CLK => CLK, RESET 
                           => RESET, ENABLE => enable_io_0_port, RD1 => 
                           io_read1_3_port, RD2 => io_read2_3_port, WR => 
                           io_write_3_port, ADD_WR(1) => ADD_WR(1), ADD_WR(0) 
                           => ADD_WR(0), ADD_RD1(1) => ADD_RD1(1), ADD_RD1(0) 
                           => ADD_RD1(0), ADD_RD2(1) => ADD_RD2(1), ADD_RD2(0) 
                           => ADD_RD2(0), DATAIN(63) => DATAIN(63), DATAIN(62) 
                           => DATAIN(62), DATAIN(61) => DATAIN(61), DATAIN(60) 
                           => DATAIN(60), DATAIN(59) => DATAIN(59), DATAIN(58) 
                           => DATAIN(58), DATAIN(57) => DATAIN(57), DATAIN(56) 
                           => DATAIN(56), DATAIN(55) => DATAIN(55), DATAIN(54) 
                           => DATAIN(54), DATAIN(53) => DATAIN(53), DATAIN(52) 
                           => DATAIN(52), DATAIN(51) => DATAIN(51), DATAIN(50) 
                           => DATAIN(50), DATAIN(49) => DATAIN(49), DATAIN(48) 
                           => DATAIN(48), DATAIN(47) => DATAIN(47), DATAIN(46) 
                           => DATAIN(46), DATAIN(45) => DATAIN(45), DATAIN(44) 
                           => DATAIN(44), DATAIN(43) => DATAIN(43), DATAIN(42) 
                           => DATAIN(42), DATAIN(41) => DATAIN(41), DATAIN(40) 
                           => DATAIN(40), DATAIN(39) => DATAIN(39), DATAIN(38) 
                           => DATAIN(38), DATAIN(37) => DATAIN(37), DATAIN(36) 
                           => DATAIN(36), DATAIN(35) => DATAIN(35), DATAIN(34) 
                           => DATAIN(34), DATAIN(33) => DATAIN(33), DATAIN(32) 
                           => DATAIN(32), DATAIN(31) => DATAIN(31), DATAIN(30) 
                           => DATAIN(30), DATAIN(29) => DATAIN(29), DATAIN(28) 
                           => DATAIN(28), DATAIN(27) => DATAIN(27), DATAIN(26) 
                           => DATAIN(26), DATAIN(25) => DATAIN(25), DATAIN(24) 
                           => DATAIN(24), DATAIN(23) => DATAIN(23), DATAIN(22) 
                           => DATAIN(22), DATAIN(21) => DATAIN(21), DATAIN(20) 
                           => DATAIN(20), DATAIN(19) => DATAIN(19), DATAIN(18) 
                           => DATAIN(18), DATAIN(17) => DATAIN(17), DATAIN(16) 
                           => DATAIN(16), DATAIN(15) => DATAIN(15), DATAIN(14) 
                           => DATAIN(14), DATAIN(13) => DATAIN(13), DATAIN(12) 
                           => DATAIN(12), DATAIN(11) => DATAIN(11), DATAIN(10) 
                           => DATAIN(10), DATAIN(9) => DATAIN(9), DATAIN(8) => 
                           DATAIN(8), DATAIN(7) => DATAIN(7), DATAIN(6) => 
                           DATAIN(6), DATAIN(5) => DATAIN(5), DATAIN(4) => 
                           DATAIN(4), DATAIN(3) => DATAIN(3), DATAIN(2) => 
                           DATAIN(2), DATAIN(1) => DATAIN(1), DATAIN(0) => 
                           DATAIN(0), OUT1(63) => io_out1_0_63_port, OUT1(62) 
                           => io_out1_0_62_port, OUT1(61) => io_out1_0_61_port,
                           OUT1(60) => io_out1_0_60_port, OUT1(59) => 
                           io_out1_0_59_port, OUT1(58) => io_out1_0_58_port, 
                           OUT1(57) => io_out1_0_57_port, OUT1(56) => 
                           io_out1_0_56_port, OUT1(55) => io_out1_0_55_port, 
                           OUT1(54) => io_out1_0_54_port, OUT1(53) => 
                           io_out1_0_53_port, OUT1(52) => io_out1_0_52_port, 
                           OUT1(51) => io_out1_0_51_port, OUT1(50) => 
                           io_out1_0_50_port, OUT1(49) => io_out1_0_49_port, 
                           OUT1(48) => io_out1_0_48_port, OUT1(47) => 
                           io_out1_0_47_port, OUT1(46) => io_out1_0_46_port, 
                           OUT1(45) => io_out1_0_45_port, OUT1(44) => 
                           io_out1_0_44_port, OUT1(43) => io_out1_0_43_port, 
                           OUT1(42) => io_out1_0_42_port, OUT1(41) => 
                           io_out1_0_41_port, OUT1(40) => io_out1_0_40_port, 
                           OUT1(39) => io_out1_0_39_port, OUT1(38) => 
                           io_out1_0_38_port, OUT1(37) => io_out1_0_37_port, 
                           OUT1(36) => io_out1_0_36_port, OUT1(35) => 
                           io_out1_0_35_port, OUT1(34) => io_out1_0_34_port, 
                           OUT1(33) => io_out1_0_33_port, OUT1(32) => 
                           io_out1_0_32_port, OUT1(31) => io_out1_0_31_port, 
                           OUT1(30) => io_out1_0_30_port, OUT1(29) => 
                           io_out1_0_29_port, OUT1(28) => io_out1_0_28_port, 
                           OUT1(27) => io_out1_0_27_port, OUT1(26) => 
                           io_out1_0_26_port, OUT1(25) => io_out1_0_25_port, 
                           OUT1(24) => io_out1_0_24_port, OUT1(23) => 
                           io_out1_0_23_port, OUT1(22) => io_out1_0_22_port, 
                           OUT1(21) => io_out1_0_21_port, OUT1(20) => 
                           io_out1_0_20_port, OUT1(19) => io_out1_0_19_port, 
                           OUT1(18) => io_out1_0_18_port, OUT1(17) => 
                           io_out1_0_17_port, OUT1(16) => io_out1_0_16_port, 
                           OUT1(15) => io_out1_0_15_port, OUT1(14) => 
                           io_out1_0_14_port, OUT1(13) => io_out1_0_13_port, 
                           OUT1(12) => io_out1_0_12_port, OUT1(11) => 
                           io_out1_0_11_port, OUT1(10) => io_out1_0_10_port, 
                           OUT1(9) => io_out1_0_9_port, OUT1(8) => 
                           io_out1_0_8_port, OUT1(7) => io_out1_0_7_port, 
                           OUT1(6) => io_out1_0_6_port, OUT1(5) => 
                           io_out1_0_5_port, OUT1(4) => io_out1_0_4_port, 
                           OUT1(3) => io_out1_0_3_port, OUT1(2) => 
                           io_out1_0_2_port, OUT1(1) => io_out1_0_1_port, 
                           OUT1(0) => io_out1_0_0_port, OUT2(63) => 
                           io_out2_0_63_port, OUT2(62) => io_out2_0_62_port, 
                           OUT2(61) => io_out2_0_61_port, OUT2(60) => 
                           io_out2_0_60_port, OUT2(59) => io_out2_0_59_port, 
                           OUT2(58) => io_out2_0_58_port, OUT2(57) => 
                           io_out2_0_57_port, OUT2(56) => io_out2_0_56_port, 
                           OUT2(55) => io_out2_0_55_port, OUT2(54) => 
                           io_out2_0_54_port, OUT2(53) => io_out2_0_53_port, 
                           OUT2(52) => io_out2_0_52_port, OUT2(51) => 
                           io_out2_0_51_port, OUT2(50) => io_out2_0_50_port, 
                           OUT2(49) => io_out2_0_49_port, OUT2(48) => 
                           io_out2_0_48_port, OUT2(47) => io_out2_0_47_port, 
                           OUT2(46) => io_out2_0_46_port, OUT2(45) => 
                           io_out2_0_45_port, OUT2(44) => io_out2_0_44_port, 
                           OUT2(43) => io_out2_0_43_port, OUT2(42) => 
                           io_out2_0_42_port, OUT2(41) => io_out2_0_41_port, 
                           OUT2(40) => io_out2_0_40_port, OUT2(39) => 
                           io_out2_0_39_port, OUT2(38) => io_out2_0_38_port, 
                           OUT2(37) => io_out2_0_37_port, OUT2(36) => 
                           io_out2_0_36_port, OUT2(35) => io_out2_0_35_port, 
                           OUT2(34) => io_out2_0_34_port, OUT2(33) => 
                           io_out2_0_33_port, OUT2(32) => io_out2_0_32_port, 
                           OUT2(31) => io_out2_0_31_port, OUT2(30) => 
                           io_out2_0_30_port, OUT2(29) => io_out2_0_29_port, 
                           OUT2(28) => io_out2_0_28_port, OUT2(27) => 
                           io_out2_0_27_port, OUT2(26) => io_out2_0_26_port, 
                           OUT2(25) => io_out2_0_25_port, OUT2(24) => 
                           io_out2_0_24_port, OUT2(23) => io_out2_0_23_port, 
                           OUT2(22) => io_out2_0_22_port, OUT2(21) => 
                           io_out2_0_21_port, OUT2(20) => io_out2_0_20_port, 
                           OUT2(19) => io_out2_0_19_port, OUT2(18) => 
                           io_out2_0_18_port, OUT2(17) => io_out2_0_17_port, 
                           OUT2(16) => io_out2_0_16_port, OUT2(15) => 
                           io_out2_0_15_port, OUT2(14) => io_out2_0_14_port, 
                           OUT2(13) => io_out2_0_13_port, OUT2(12) => 
                           io_out2_0_12_port, OUT2(11) => io_out2_0_11_port, 
                           OUT2(10) => io_out2_0_10_port, OUT2(9) => 
                           io_out2_0_9_port, OUT2(8) => io_out2_0_8_port, 
                           OUT2(7) => io_out2_0_7_port, OUT2(6) => 
                           io_out2_0_6_port, OUT2(5) => io_out2_0_5_port, 
                           OUT2(4) => io_out2_0_4_port, OUT2(3) => 
                           io_out2_0_3_port, OUT2(2) => io_out2_0_2_port, 
                           OUT2(1) => io_out2_0_1_port, OUT2(0) => 
                           io_out2_0_0_port);
   loc_rf_0 : register_file_reg_size64_file_size4_7 port map( CLK => CLK, RESET
                           => RESET, ENABLE => enable_loc_0_port, RD1 => 
                           loc_read1_3_port, RD2 => loc_read2_3_port, WR => 
                           loc_write_3_port, ADD_WR(1) => ADD_WR(1), ADD_WR(0) 
                           => ADD_WR(0), ADD_RD1(1) => ADD_RD1(1), ADD_RD1(0) 
                           => ADD_RD1(0), ADD_RD2(1) => ADD_RD2(1), ADD_RD2(0) 
                           => ADD_RD2(0), DATAIN(63) => DATAIN(63), DATAIN(62) 
                           => DATAIN(62), DATAIN(61) => DATAIN(61), DATAIN(60) 
                           => DATAIN(60), DATAIN(59) => DATAIN(59), DATAIN(58) 
                           => DATAIN(58), DATAIN(57) => DATAIN(57), DATAIN(56) 
                           => DATAIN(56), DATAIN(55) => DATAIN(55), DATAIN(54) 
                           => DATAIN(54), DATAIN(53) => DATAIN(53), DATAIN(52) 
                           => DATAIN(52), DATAIN(51) => DATAIN(51), DATAIN(50) 
                           => DATAIN(50), DATAIN(49) => DATAIN(49), DATAIN(48) 
                           => DATAIN(48), DATAIN(47) => DATAIN(47), DATAIN(46) 
                           => DATAIN(46), DATAIN(45) => DATAIN(45), DATAIN(44) 
                           => DATAIN(44), DATAIN(43) => DATAIN(43), DATAIN(42) 
                           => DATAIN(42), DATAIN(41) => DATAIN(41), DATAIN(40) 
                           => DATAIN(40), DATAIN(39) => DATAIN(39), DATAIN(38) 
                           => DATAIN(38), DATAIN(37) => DATAIN(37), DATAIN(36) 
                           => DATAIN(36), DATAIN(35) => DATAIN(35), DATAIN(34) 
                           => DATAIN(34), DATAIN(33) => DATAIN(33), DATAIN(32) 
                           => DATAIN(32), DATAIN(31) => DATAIN(31), DATAIN(30) 
                           => DATAIN(30), DATAIN(29) => DATAIN(29), DATAIN(28) 
                           => DATAIN(28), DATAIN(27) => DATAIN(27), DATAIN(26) 
                           => DATAIN(26), DATAIN(25) => DATAIN(25), DATAIN(24) 
                           => DATAIN(24), DATAIN(23) => DATAIN(23), DATAIN(22) 
                           => DATAIN(22), DATAIN(21) => DATAIN(21), DATAIN(20) 
                           => DATAIN(20), DATAIN(19) => DATAIN(19), DATAIN(18) 
                           => DATAIN(18), DATAIN(17) => DATAIN(17), DATAIN(16) 
                           => DATAIN(16), DATAIN(15) => DATAIN(15), DATAIN(14) 
                           => DATAIN(14), DATAIN(13) => DATAIN(13), DATAIN(12) 
                           => DATAIN(12), DATAIN(11) => DATAIN(11), DATAIN(10) 
                           => DATAIN(10), DATAIN(9) => DATAIN(9), DATAIN(8) => 
                           DATAIN(8), DATAIN(7) => DATAIN(7), DATAIN(6) => 
                           DATAIN(6), DATAIN(5) => DATAIN(5), DATAIN(4) => 
                           DATAIN(4), DATAIN(3) => DATAIN(3), DATAIN(2) => 
                           DATAIN(2), DATAIN(1) => DATAIN(1), DATAIN(0) => 
                           DATAIN(0), OUT1(63) => loc_out1_0_63_port, OUT1(62) 
                           => loc_out1_0_62_port, OUT1(61) => 
                           loc_out1_0_61_port, OUT1(60) => loc_out1_0_60_port, 
                           OUT1(59) => loc_out1_0_59_port, OUT1(58) => 
                           loc_out1_0_58_port, OUT1(57) => loc_out1_0_57_port, 
                           OUT1(56) => loc_out1_0_56_port, OUT1(55) => 
                           loc_out1_0_55_port, OUT1(54) => loc_out1_0_54_port, 
                           OUT1(53) => loc_out1_0_53_port, OUT1(52) => 
                           loc_out1_0_52_port, OUT1(51) => loc_out1_0_51_port, 
                           OUT1(50) => loc_out1_0_50_port, OUT1(49) => 
                           loc_out1_0_49_port, OUT1(48) => loc_out1_0_48_port, 
                           OUT1(47) => loc_out1_0_47_port, OUT1(46) => 
                           loc_out1_0_46_port, OUT1(45) => loc_out1_0_45_port, 
                           OUT1(44) => loc_out1_0_44_port, OUT1(43) => 
                           loc_out1_0_43_port, OUT1(42) => loc_out1_0_42_port, 
                           OUT1(41) => loc_out1_0_41_port, OUT1(40) => 
                           loc_out1_0_40_port, OUT1(39) => loc_out1_0_39_port, 
                           OUT1(38) => loc_out1_0_38_port, OUT1(37) => 
                           loc_out1_0_37_port, OUT1(36) => loc_out1_0_36_port, 
                           OUT1(35) => loc_out1_0_35_port, OUT1(34) => 
                           loc_out1_0_34_port, OUT1(33) => loc_out1_0_33_port, 
                           OUT1(32) => loc_out1_0_32_port, OUT1(31) => 
                           loc_out1_0_31_port, OUT1(30) => loc_out1_0_30_port, 
                           OUT1(29) => loc_out1_0_29_port, OUT1(28) => 
                           loc_out1_0_28_port, OUT1(27) => loc_out1_0_27_port, 
                           OUT1(26) => loc_out1_0_26_port, OUT1(25) => 
                           loc_out1_0_25_port, OUT1(24) => loc_out1_0_24_port, 
                           OUT1(23) => loc_out1_0_23_port, OUT1(22) => 
                           loc_out1_0_22_port, OUT1(21) => loc_out1_0_21_port, 
                           OUT1(20) => loc_out1_0_20_port, OUT1(19) => 
                           loc_out1_0_19_port, OUT1(18) => loc_out1_0_18_port, 
                           OUT1(17) => loc_out1_0_17_port, OUT1(16) => 
                           loc_out1_0_16_port, OUT1(15) => loc_out1_0_15_port, 
                           OUT1(14) => loc_out1_0_14_port, OUT1(13) => 
                           loc_out1_0_13_port, OUT1(12) => loc_out1_0_12_port, 
                           OUT1(11) => loc_out1_0_11_port, OUT1(10) => 
                           loc_out1_0_10_port, OUT1(9) => loc_out1_0_9_port, 
                           OUT1(8) => loc_out1_0_8_port, OUT1(7) => 
                           loc_out1_0_7_port, OUT1(6) => loc_out1_0_6_port, 
                           OUT1(5) => loc_out1_0_5_port, OUT1(4) => 
                           loc_out1_0_4_port, OUT1(3) => loc_out1_0_3_port, 
                           OUT1(2) => loc_out1_0_2_port, OUT1(1) => 
                           loc_out1_0_1_port, OUT1(0) => loc_out1_0_0_port, 
                           OUT2(63) => loc_out2_0_63_port, OUT2(62) => 
                           loc_out2_0_62_port, OUT2(61) => loc_out2_0_61_port, 
                           OUT2(60) => loc_out2_0_60_port, OUT2(59) => 
                           loc_out2_0_59_port, OUT2(58) => loc_out2_0_58_port, 
                           OUT2(57) => loc_out2_0_57_port, OUT2(56) => 
                           loc_out2_0_56_port, OUT2(55) => loc_out2_0_55_port, 
                           OUT2(54) => loc_out2_0_54_port, OUT2(53) => 
                           loc_out2_0_53_port, OUT2(52) => loc_out2_0_52_port, 
                           OUT2(51) => loc_out2_0_51_port, OUT2(50) => 
                           loc_out2_0_50_port, OUT2(49) => loc_out2_0_49_port, 
                           OUT2(48) => loc_out2_0_48_port, OUT2(47) => 
                           loc_out2_0_47_port, OUT2(46) => loc_out2_0_46_port, 
                           OUT2(45) => loc_out2_0_45_port, OUT2(44) => 
                           loc_out2_0_44_port, OUT2(43) => loc_out2_0_43_port, 
                           OUT2(42) => loc_out2_0_42_port, OUT2(41) => 
                           loc_out2_0_41_port, OUT2(40) => loc_out2_0_40_port, 
                           OUT2(39) => loc_out2_0_39_port, OUT2(38) => 
                           loc_out2_0_38_port, OUT2(37) => loc_out2_0_37_port, 
                           OUT2(36) => loc_out2_0_36_port, OUT2(35) => 
                           loc_out2_0_35_port, OUT2(34) => loc_out2_0_34_port, 
                           OUT2(33) => loc_out2_0_33_port, OUT2(32) => 
                           loc_out2_0_32_port, OUT2(31) => loc_out2_0_31_port, 
                           OUT2(30) => loc_out2_0_30_port, OUT2(29) => 
                           loc_out2_0_29_port, OUT2(28) => loc_out2_0_28_port, 
                           OUT2(27) => loc_out2_0_27_port, OUT2(26) => 
                           loc_out2_0_26_port, OUT2(25) => loc_out2_0_25_port, 
                           OUT2(24) => loc_out2_0_24_port, OUT2(23) => 
                           loc_out2_0_23_port, OUT2(22) => loc_out2_0_22_port, 
                           OUT2(21) => loc_out2_0_21_port, OUT2(20) => 
                           loc_out2_0_20_port, OUT2(19) => loc_out2_0_19_port, 
                           OUT2(18) => loc_out2_0_18_port, OUT2(17) => 
                           loc_out2_0_17_port, OUT2(16) => loc_out2_0_16_port, 
                           OUT2(15) => loc_out2_0_15_port, OUT2(14) => 
                           loc_out2_0_14_port, OUT2(13) => loc_out2_0_13_port, 
                           OUT2(12) => loc_out2_0_12_port, OUT2(11) => 
                           loc_out2_0_11_port, OUT2(10) => loc_out2_0_10_port, 
                           OUT2(9) => loc_out2_0_9_port, OUT2(8) => 
                           loc_out2_0_8_port, OUT2(7) => loc_out2_0_7_port, 
                           OUT2(6) => loc_out2_0_6_port, OUT2(5) => 
                           loc_out2_0_5_port, OUT2(4) => loc_out2_0_4_port, 
                           OUT2(3) => loc_out2_0_3_port, OUT2(2) => 
                           loc_out2_0_2_port, OUT2(1) => loc_out2_0_1_port, 
                           OUT2(0) => loc_out2_0_0_port);
   io_rf_1 : register_file_reg_size64_file_size4_6 port map( CLK => CLK, RESET 
                           => RESET, ENABLE => enable_io_1_port, RD1 => 
                           io_read1_3_port, RD2 => io_read2_3_port, WR => 
                           io_write_3_port, ADD_WR(1) => ADD_WR(1), ADD_WR(0) 
                           => ADD_WR(0), ADD_RD1(1) => ADD_RD1(1), ADD_RD1(0) 
                           => ADD_RD1(0), ADD_RD2(1) => ADD_RD2(1), ADD_RD2(0) 
                           => ADD_RD2(0), DATAIN(63) => DATAIN(63), DATAIN(62) 
                           => DATAIN(62), DATAIN(61) => DATAIN(61), DATAIN(60) 
                           => DATAIN(60), DATAIN(59) => DATAIN(59), DATAIN(58) 
                           => DATAIN(58), DATAIN(57) => DATAIN(57), DATAIN(56) 
                           => DATAIN(56), DATAIN(55) => DATAIN(55), DATAIN(54) 
                           => DATAIN(54), DATAIN(53) => DATAIN(53), DATAIN(52) 
                           => DATAIN(52), DATAIN(51) => DATAIN(51), DATAIN(50) 
                           => DATAIN(50), DATAIN(49) => DATAIN(49), DATAIN(48) 
                           => DATAIN(48), DATAIN(47) => DATAIN(47), DATAIN(46) 
                           => DATAIN(46), DATAIN(45) => DATAIN(45), DATAIN(44) 
                           => DATAIN(44), DATAIN(43) => DATAIN(43), DATAIN(42) 
                           => DATAIN(42), DATAIN(41) => DATAIN(41), DATAIN(40) 
                           => DATAIN(40), DATAIN(39) => DATAIN(39), DATAIN(38) 
                           => DATAIN(38), DATAIN(37) => DATAIN(37), DATAIN(36) 
                           => DATAIN(36), DATAIN(35) => DATAIN(35), DATAIN(34) 
                           => DATAIN(34), DATAIN(33) => DATAIN(33), DATAIN(32) 
                           => DATAIN(32), DATAIN(31) => DATAIN(31), DATAIN(30) 
                           => DATAIN(30), DATAIN(29) => DATAIN(29), DATAIN(28) 
                           => DATAIN(28), DATAIN(27) => DATAIN(27), DATAIN(26) 
                           => DATAIN(26), DATAIN(25) => DATAIN(25), DATAIN(24) 
                           => DATAIN(24), DATAIN(23) => DATAIN(23), DATAIN(22) 
                           => DATAIN(22), DATAIN(21) => DATAIN(21), DATAIN(20) 
                           => DATAIN(20), DATAIN(19) => DATAIN(19), DATAIN(18) 
                           => DATAIN(18), DATAIN(17) => DATAIN(17), DATAIN(16) 
                           => DATAIN(16), DATAIN(15) => DATAIN(15), DATAIN(14) 
                           => DATAIN(14), DATAIN(13) => DATAIN(13), DATAIN(12) 
                           => DATAIN(12), DATAIN(11) => DATAIN(11), DATAIN(10) 
                           => DATAIN(10), DATAIN(9) => DATAIN(9), DATAIN(8) => 
                           DATAIN(8), DATAIN(7) => DATAIN(7), DATAIN(6) => 
                           DATAIN(6), DATAIN(5) => DATAIN(5), DATAIN(4) => 
                           DATAIN(4), DATAIN(3) => DATAIN(3), DATAIN(2) => 
                           DATAIN(2), DATAIN(1) => DATAIN(1), DATAIN(0) => 
                           DATAIN(0), OUT1(63) => io_out1_1_63_port, OUT1(62) 
                           => io_out1_1_62_port, OUT1(61) => io_out1_1_61_port,
                           OUT1(60) => io_out1_1_60_port, OUT1(59) => 
                           io_out1_1_59_port, OUT1(58) => io_out1_1_58_port, 
                           OUT1(57) => io_out1_1_57_port, OUT1(56) => 
                           io_out1_1_56_port, OUT1(55) => io_out1_1_55_port, 
                           OUT1(54) => io_out1_1_54_port, OUT1(53) => 
                           io_out1_1_53_port, OUT1(52) => io_out1_1_52_port, 
                           OUT1(51) => io_out1_1_51_port, OUT1(50) => 
                           io_out1_1_50_port, OUT1(49) => io_out1_1_49_port, 
                           OUT1(48) => io_out1_1_48_port, OUT1(47) => 
                           io_out1_1_47_port, OUT1(46) => io_out1_1_46_port, 
                           OUT1(45) => io_out1_1_45_port, OUT1(44) => 
                           io_out1_1_44_port, OUT1(43) => io_out1_1_43_port, 
                           OUT1(42) => io_out1_1_42_port, OUT1(41) => 
                           io_out1_1_41_port, OUT1(40) => io_out1_1_40_port, 
                           OUT1(39) => io_out1_1_39_port, OUT1(38) => 
                           io_out1_1_38_port, OUT1(37) => io_out1_1_37_port, 
                           OUT1(36) => io_out1_1_36_port, OUT1(35) => 
                           io_out1_1_35_port, OUT1(34) => io_out1_1_34_port, 
                           OUT1(33) => io_out1_1_33_port, OUT1(32) => 
                           io_out1_1_32_port, OUT1(31) => io_out1_1_31_port, 
                           OUT1(30) => io_out1_1_30_port, OUT1(29) => 
                           io_out1_1_29_port, OUT1(28) => io_out1_1_28_port, 
                           OUT1(27) => io_out1_1_27_port, OUT1(26) => 
                           io_out1_1_26_port, OUT1(25) => io_out1_1_25_port, 
                           OUT1(24) => io_out1_1_24_port, OUT1(23) => 
                           io_out1_1_23_port, OUT1(22) => io_out1_1_22_port, 
                           OUT1(21) => io_out1_1_21_port, OUT1(20) => 
                           io_out1_1_20_port, OUT1(19) => io_out1_1_19_port, 
                           OUT1(18) => io_out1_1_18_port, OUT1(17) => 
                           io_out1_1_17_port, OUT1(16) => io_out1_1_16_port, 
                           OUT1(15) => io_out1_1_15_port, OUT1(14) => 
                           io_out1_1_14_port, OUT1(13) => io_out1_1_13_port, 
                           OUT1(12) => io_out1_1_12_port, OUT1(11) => 
                           io_out1_1_11_port, OUT1(10) => io_out1_1_10_port, 
                           OUT1(9) => io_out1_1_9_port, OUT1(8) => 
                           io_out1_1_8_port, OUT1(7) => io_out1_1_7_port, 
                           OUT1(6) => io_out1_1_6_port, OUT1(5) => 
                           io_out1_1_5_port, OUT1(4) => io_out1_1_4_port, 
                           OUT1(3) => io_out1_1_3_port, OUT1(2) => 
                           io_out1_1_2_port, OUT1(1) => io_out1_1_1_port, 
                           OUT1(0) => io_out1_1_0_port, OUT2(63) => 
                           io_out2_1_63_port, OUT2(62) => io_out2_1_62_port, 
                           OUT2(61) => io_out2_1_61_port, OUT2(60) => 
                           io_out2_1_60_port, OUT2(59) => io_out2_1_59_port, 
                           OUT2(58) => io_out2_1_58_port, OUT2(57) => 
                           io_out2_1_57_port, OUT2(56) => io_out2_1_56_port, 
                           OUT2(55) => io_out2_1_55_port, OUT2(54) => 
                           io_out2_1_54_port, OUT2(53) => io_out2_1_53_port, 
                           OUT2(52) => io_out2_1_52_port, OUT2(51) => 
                           io_out2_1_51_port, OUT2(50) => io_out2_1_50_port, 
                           OUT2(49) => io_out2_1_49_port, OUT2(48) => 
                           io_out2_1_48_port, OUT2(47) => io_out2_1_47_port, 
                           OUT2(46) => io_out2_1_46_port, OUT2(45) => 
                           io_out2_1_45_port, OUT2(44) => io_out2_1_44_port, 
                           OUT2(43) => io_out2_1_43_port, OUT2(42) => 
                           io_out2_1_42_port, OUT2(41) => io_out2_1_41_port, 
                           OUT2(40) => io_out2_1_40_port, OUT2(39) => 
                           io_out2_1_39_port, OUT2(38) => io_out2_1_38_port, 
                           OUT2(37) => io_out2_1_37_port, OUT2(36) => 
                           io_out2_1_36_port, OUT2(35) => io_out2_1_35_port, 
                           OUT2(34) => io_out2_1_34_port, OUT2(33) => 
                           io_out2_1_33_port, OUT2(32) => io_out2_1_32_port, 
                           OUT2(31) => io_out2_1_31_port, OUT2(30) => 
                           io_out2_1_30_port, OUT2(29) => io_out2_1_29_port, 
                           OUT2(28) => io_out2_1_28_port, OUT2(27) => 
                           io_out2_1_27_port, OUT2(26) => io_out2_1_26_port, 
                           OUT2(25) => io_out2_1_25_port, OUT2(24) => 
                           io_out2_1_24_port, OUT2(23) => io_out2_1_23_port, 
                           OUT2(22) => io_out2_1_22_port, OUT2(21) => 
                           io_out2_1_21_port, OUT2(20) => io_out2_1_20_port, 
                           OUT2(19) => io_out2_1_19_port, OUT2(18) => 
                           io_out2_1_18_port, OUT2(17) => io_out2_1_17_port, 
                           OUT2(16) => io_out2_1_16_port, OUT2(15) => 
                           io_out2_1_15_port, OUT2(14) => io_out2_1_14_port, 
                           OUT2(13) => io_out2_1_13_port, OUT2(12) => 
                           io_out2_1_12_port, OUT2(11) => io_out2_1_11_port, 
                           OUT2(10) => io_out2_1_10_port, OUT2(9) => 
                           io_out2_1_9_port, OUT2(8) => io_out2_1_8_port, 
                           OUT2(7) => io_out2_1_7_port, OUT2(6) => 
                           io_out2_1_6_port, OUT2(5) => io_out2_1_5_port, 
                           OUT2(4) => io_out2_1_4_port, OUT2(3) => 
                           io_out2_1_3_port, OUT2(2) => io_out2_1_2_port, 
                           OUT2(1) => io_out2_1_1_port, OUT2(0) => 
                           io_out2_1_0_port);
   loc_rf_1 : register_file_reg_size64_file_size4_5 port map( CLK => CLK, RESET
                           => RESET, ENABLE => enable_loc_1_port, RD1 => 
                           loc_read1_3_port, RD2 => loc_read2_3_port, WR => 
                           loc_write_3_port, ADD_WR(1) => ADD_WR(1), ADD_WR(0) 
                           => ADD_WR(0), ADD_RD1(1) => ADD_RD1(1), ADD_RD1(0) 
                           => ADD_RD1(0), ADD_RD2(1) => ADD_RD2(1), ADD_RD2(0) 
                           => ADD_RD2(0), DATAIN(63) => DATAIN(63), DATAIN(62) 
                           => DATAIN(62), DATAIN(61) => DATAIN(61), DATAIN(60) 
                           => DATAIN(60), DATAIN(59) => DATAIN(59), DATAIN(58) 
                           => DATAIN(58), DATAIN(57) => DATAIN(57), DATAIN(56) 
                           => DATAIN(56), DATAIN(55) => DATAIN(55), DATAIN(54) 
                           => DATAIN(54), DATAIN(53) => DATAIN(53), DATAIN(52) 
                           => DATAIN(52), DATAIN(51) => DATAIN(51), DATAIN(50) 
                           => DATAIN(50), DATAIN(49) => DATAIN(49), DATAIN(48) 
                           => DATAIN(48), DATAIN(47) => DATAIN(47), DATAIN(46) 
                           => DATAIN(46), DATAIN(45) => DATAIN(45), DATAIN(44) 
                           => DATAIN(44), DATAIN(43) => DATAIN(43), DATAIN(42) 
                           => DATAIN(42), DATAIN(41) => DATAIN(41), DATAIN(40) 
                           => DATAIN(40), DATAIN(39) => DATAIN(39), DATAIN(38) 
                           => DATAIN(38), DATAIN(37) => DATAIN(37), DATAIN(36) 
                           => DATAIN(36), DATAIN(35) => DATAIN(35), DATAIN(34) 
                           => DATAIN(34), DATAIN(33) => DATAIN(33), DATAIN(32) 
                           => DATAIN(32), DATAIN(31) => DATAIN(31), DATAIN(30) 
                           => DATAIN(30), DATAIN(29) => DATAIN(29), DATAIN(28) 
                           => DATAIN(28), DATAIN(27) => DATAIN(27), DATAIN(26) 
                           => DATAIN(26), DATAIN(25) => DATAIN(25), DATAIN(24) 
                           => DATAIN(24), DATAIN(23) => DATAIN(23), DATAIN(22) 
                           => DATAIN(22), DATAIN(21) => DATAIN(21), DATAIN(20) 
                           => DATAIN(20), DATAIN(19) => DATAIN(19), DATAIN(18) 
                           => DATAIN(18), DATAIN(17) => DATAIN(17), DATAIN(16) 
                           => DATAIN(16), DATAIN(15) => DATAIN(15), DATAIN(14) 
                           => DATAIN(14), DATAIN(13) => DATAIN(13), DATAIN(12) 
                           => DATAIN(12), DATAIN(11) => DATAIN(11), DATAIN(10) 
                           => DATAIN(10), DATAIN(9) => DATAIN(9), DATAIN(8) => 
                           DATAIN(8), DATAIN(7) => DATAIN(7), DATAIN(6) => 
                           DATAIN(6), DATAIN(5) => DATAIN(5), DATAIN(4) => 
                           DATAIN(4), DATAIN(3) => DATAIN(3), DATAIN(2) => 
                           DATAIN(2), DATAIN(1) => DATAIN(1), DATAIN(0) => 
                           DATAIN(0), OUT1(63) => loc_out1_1_63_port, OUT1(62) 
                           => loc_out1_1_62_port, OUT1(61) => 
                           loc_out1_1_61_port, OUT1(60) => loc_out1_1_60_port, 
                           OUT1(59) => loc_out1_1_59_port, OUT1(58) => 
                           loc_out1_1_58_port, OUT1(57) => loc_out1_1_57_port, 
                           OUT1(56) => loc_out1_1_56_port, OUT1(55) => 
                           loc_out1_1_55_port, OUT1(54) => loc_out1_1_54_port, 
                           OUT1(53) => loc_out1_1_53_port, OUT1(52) => 
                           loc_out1_1_52_port, OUT1(51) => loc_out1_1_51_port, 
                           OUT1(50) => loc_out1_1_50_port, OUT1(49) => 
                           loc_out1_1_49_port, OUT1(48) => loc_out1_1_48_port, 
                           OUT1(47) => loc_out1_1_47_port, OUT1(46) => 
                           loc_out1_1_46_port, OUT1(45) => loc_out1_1_45_port, 
                           OUT1(44) => loc_out1_1_44_port, OUT1(43) => 
                           loc_out1_1_43_port, OUT1(42) => loc_out1_1_42_port, 
                           OUT1(41) => loc_out1_1_41_port, OUT1(40) => 
                           loc_out1_1_40_port, OUT1(39) => loc_out1_1_39_port, 
                           OUT1(38) => loc_out1_1_38_port, OUT1(37) => 
                           loc_out1_1_37_port, OUT1(36) => loc_out1_1_36_port, 
                           OUT1(35) => loc_out1_1_35_port, OUT1(34) => 
                           loc_out1_1_34_port, OUT1(33) => loc_out1_1_33_port, 
                           OUT1(32) => loc_out1_1_32_port, OUT1(31) => 
                           loc_out1_1_31_port, OUT1(30) => loc_out1_1_30_port, 
                           OUT1(29) => loc_out1_1_29_port, OUT1(28) => 
                           loc_out1_1_28_port, OUT1(27) => loc_out1_1_27_port, 
                           OUT1(26) => loc_out1_1_26_port, OUT1(25) => 
                           loc_out1_1_25_port, OUT1(24) => loc_out1_1_24_port, 
                           OUT1(23) => loc_out1_1_23_port, OUT1(22) => 
                           loc_out1_1_22_port, OUT1(21) => loc_out1_1_21_port, 
                           OUT1(20) => loc_out1_1_20_port, OUT1(19) => 
                           loc_out1_1_19_port, OUT1(18) => loc_out1_1_18_port, 
                           OUT1(17) => loc_out1_1_17_port, OUT1(16) => 
                           loc_out1_1_16_port, OUT1(15) => loc_out1_1_15_port, 
                           OUT1(14) => loc_out1_1_14_port, OUT1(13) => 
                           loc_out1_1_13_port, OUT1(12) => loc_out1_1_12_port, 
                           OUT1(11) => loc_out1_1_11_port, OUT1(10) => 
                           loc_out1_1_10_port, OUT1(9) => loc_out1_1_9_port, 
                           OUT1(8) => loc_out1_1_8_port, OUT1(7) => 
                           loc_out1_1_7_port, OUT1(6) => loc_out1_1_6_port, 
                           OUT1(5) => loc_out1_1_5_port, OUT1(4) => 
                           loc_out1_1_4_port, OUT1(3) => loc_out1_1_3_port, 
                           OUT1(2) => loc_out1_1_2_port, OUT1(1) => 
                           loc_out1_1_1_port, OUT1(0) => loc_out1_1_0_port, 
                           OUT2(63) => loc_out2_1_63_port, OUT2(62) => 
                           loc_out2_1_62_port, OUT2(61) => loc_out2_1_61_port, 
                           OUT2(60) => loc_out2_1_60_port, OUT2(59) => 
                           loc_out2_1_59_port, OUT2(58) => loc_out2_1_58_port, 
                           OUT2(57) => loc_out2_1_57_port, OUT2(56) => 
                           loc_out2_1_56_port, OUT2(55) => loc_out2_1_55_port, 
                           OUT2(54) => loc_out2_1_54_port, OUT2(53) => 
                           loc_out2_1_53_port, OUT2(52) => loc_out2_1_52_port, 
                           OUT2(51) => loc_out2_1_51_port, OUT2(50) => 
                           loc_out2_1_50_port, OUT2(49) => loc_out2_1_49_port, 
                           OUT2(48) => loc_out2_1_48_port, OUT2(47) => 
                           loc_out2_1_47_port, OUT2(46) => loc_out2_1_46_port, 
                           OUT2(45) => loc_out2_1_45_port, OUT2(44) => 
                           loc_out2_1_44_port, OUT2(43) => loc_out2_1_43_port, 
                           OUT2(42) => loc_out2_1_42_port, OUT2(41) => 
                           loc_out2_1_41_port, OUT2(40) => loc_out2_1_40_port, 
                           OUT2(39) => loc_out2_1_39_port, OUT2(38) => 
                           loc_out2_1_38_port, OUT2(37) => loc_out2_1_37_port, 
                           OUT2(36) => loc_out2_1_36_port, OUT2(35) => 
                           loc_out2_1_35_port, OUT2(34) => loc_out2_1_34_port, 
                           OUT2(33) => loc_out2_1_33_port, OUT2(32) => 
                           loc_out2_1_32_port, OUT2(31) => loc_out2_1_31_port, 
                           OUT2(30) => loc_out2_1_30_port, OUT2(29) => 
                           loc_out2_1_29_port, OUT2(28) => loc_out2_1_28_port, 
                           OUT2(27) => loc_out2_1_27_port, OUT2(26) => 
                           loc_out2_1_26_port, OUT2(25) => loc_out2_1_25_port, 
                           OUT2(24) => loc_out2_1_24_port, OUT2(23) => 
                           loc_out2_1_23_port, OUT2(22) => loc_out2_1_22_port, 
                           OUT2(21) => loc_out2_1_21_port, OUT2(20) => 
                           loc_out2_1_20_port, OUT2(19) => loc_out2_1_19_port, 
                           OUT2(18) => loc_out2_1_18_port, OUT2(17) => 
                           loc_out2_1_17_port, OUT2(16) => loc_out2_1_16_port, 
                           OUT2(15) => loc_out2_1_15_port, OUT2(14) => 
                           loc_out2_1_14_port, OUT2(13) => loc_out2_1_13_port, 
                           OUT2(12) => loc_out2_1_12_port, OUT2(11) => 
                           loc_out2_1_11_port, OUT2(10) => loc_out2_1_10_port, 
                           OUT2(9) => loc_out2_1_9_port, OUT2(8) => 
                           loc_out2_1_8_port, OUT2(7) => loc_out2_1_7_port, 
                           OUT2(6) => loc_out2_1_6_port, OUT2(5) => 
                           loc_out2_1_5_port, OUT2(4) => loc_out2_1_4_port, 
                           OUT2(3) => loc_out2_1_3_port, OUT2(2) => 
                           loc_out2_1_2_port, OUT2(1) => loc_out2_1_1_port, 
                           OUT2(0) => loc_out2_1_0_port);
   io_rf_2 : register_file_reg_size64_file_size4_4 port map( CLK => CLK, RESET 
                           => RESET, ENABLE => enable_io_2_port, RD1 => 
                           io_read1_3_port, RD2 => io_read2_3_port, WR => 
                           io_write_3_port, ADD_WR(1) => ADD_WR(1), ADD_WR(0) 
                           => ADD_WR(0), ADD_RD1(1) => ADD_RD1(1), ADD_RD1(0) 
                           => ADD_RD1(0), ADD_RD2(1) => ADD_RD2(1), ADD_RD2(0) 
                           => ADD_RD2(0), DATAIN(63) => DATAIN(63), DATAIN(62) 
                           => DATAIN(62), DATAIN(61) => DATAIN(61), DATAIN(60) 
                           => DATAIN(60), DATAIN(59) => DATAIN(59), DATAIN(58) 
                           => DATAIN(58), DATAIN(57) => DATAIN(57), DATAIN(56) 
                           => DATAIN(56), DATAIN(55) => DATAIN(55), DATAIN(54) 
                           => DATAIN(54), DATAIN(53) => DATAIN(53), DATAIN(52) 
                           => DATAIN(52), DATAIN(51) => DATAIN(51), DATAIN(50) 
                           => DATAIN(50), DATAIN(49) => DATAIN(49), DATAIN(48) 
                           => DATAIN(48), DATAIN(47) => DATAIN(47), DATAIN(46) 
                           => DATAIN(46), DATAIN(45) => DATAIN(45), DATAIN(44) 
                           => DATAIN(44), DATAIN(43) => DATAIN(43), DATAIN(42) 
                           => DATAIN(42), DATAIN(41) => DATAIN(41), DATAIN(40) 
                           => DATAIN(40), DATAIN(39) => DATAIN(39), DATAIN(38) 
                           => DATAIN(38), DATAIN(37) => DATAIN(37), DATAIN(36) 
                           => DATAIN(36), DATAIN(35) => DATAIN(35), DATAIN(34) 
                           => DATAIN(34), DATAIN(33) => DATAIN(33), DATAIN(32) 
                           => DATAIN(32), DATAIN(31) => DATAIN(31), DATAIN(30) 
                           => DATAIN(30), DATAIN(29) => DATAIN(29), DATAIN(28) 
                           => DATAIN(28), DATAIN(27) => DATAIN(27), DATAIN(26) 
                           => DATAIN(26), DATAIN(25) => DATAIN(25), DATAIN(24) 
                           => DATAIN(24), DATAIN(23) => DATAIN(23), DATAIN(22) 
                           => DATAIN(22), DATAIN(21) => DATAIN(21), DATAIN(20) 
                           => DATAIN(20), DATAIN(19) => DATAIN(19), DATAIN(18) 
                           => DATAIN(18), DATAIN(17) => DATAIN(17), DATAIN(16) 
                           => DATAIN(16), DATAIN(15) => DATAIN(15), DATAIN(14) 
                           => DATAIN(14), DATAIN(13) => DATAIN(13), DATAIN(12) 
                           => DATAIN(12), DATAIN(11) => DATAIN(11), DATAIN(10) 
                           => DATAIN(10), DATAIN(9) => DATAIN(9), DATAIN(8) => 
                           DATAIN(8), DATAIN(7) => DATAIN(7), DATAIN(6) => 
                           DATAIN(6), DATAIN(5) => DATAIN(5), DATAIN(4) => 
                           DATAIN(4), DATAIN(3) => DATAIN(3), DATAIN(2) => 
                           DATAIN(2), DATAIN(1) => DATAIN(1), DATAIN(0) => 
                           DATAIN(0), OUT1(63) => io_out1_2_63_port, OUT1(62) 
                           => io_out1_2_62_port, OUT1(61) => io_out1_2_61_port,
                           OUT1(60) => io_out1_2_60_port, OUT1(59) => 
                           io_out1_2_59_port, OUT1(58) => io_out1_2_58_port, 
                           OUT1(57) => io_out1_2_57_port, OUT1(56) => 
                           io_out1_2_56_port, OUT1(55) => io_out1_2_55_port, 
                           OUT1(54) => io_out1_2_54_port, OUT1(53) => 
                           io_out1_2_53_port, OUT1(52) => io_out1_2_52_port, 
                           OUT1(51) => io_out1_2_51_port, OUT1(50) => 
                           io_out1_2_50_port, OUT1(49) => io_out1_2_49_port, 
                           OUT1(48) => io_out1_2_48_port, OUT1(47) => 
                           io_out1_2_47_port, OUT1(46) => io_out1_2_46_port, 
                           OUT1(45) => io_out1_2_45_port, OUT1(44) => 
                           io_out1_2_44_port, OUT1(43) => io_out1_2_43_port, 
                           OUT1(42) => io_out1_2_42_port, OUT1(41) => 
                           io_out1_2_41_port, OUT1(40) => io_out1_2_40_port, 
                           OUT1(39) => io_out1_2_39_port, OUT1(38) => 
                           io_out1_2_38_port, OUT1(37) => io_out1_2_37_port, 
                           OUT1(36) => io_out1_2_36_port, OUT1(35) => 
                           io_out1_2_35_port, OUT1(34) => io_out1_2_34_port, 
                           OUT1(33) => io_out1_2_33_port, OUT1(32) => 
                           io_out1_2_32_port, OUT1(31) => io_out1_2_31_port, 
                           OUT1(30) => io_out1_2_30_port, OUT1(29) => 
                           io_out1_2_29_port, OUT1(28) => io_out1_2_28_port, 
                           OUT1(27) => io_out1_2_27_port, OUT1(26) => 
                           io_out1_2_26_port, OUT1(25) => io_out1_2_25_port, 
                           OUT1(24) => io_out1_2_24_port, OUT1(23) => 
                           io_out1_2_23_port, OUT1(22) => io_out1_2_22_port, 
                           OUT1(21) => io_out1_2_21_port, OUT1(20) => 
                           io_out1_2_20_port, OUT1(19) => io_out1_2_19_port, 
                           OUT1(18) => io_out1_2_18_port, OUT1(17) => 
                           io_out1_2_17_port, OUT1(16) => io_out1_2_16_port, 
                           OUT1(15) => io_out1_2_15_port, OUT1(14) => 
                           io_out1_2_14_port, OUT1(13) => io_out1_2_13_port, 
                           OUT1(12) => io_out1_2_12_port, OUT1(11) => 
                           io_out1_2_11_port, OUT1(10) => io_out1_2_10_port, 
                           OUT1(9) => io_out1_2_9_port, OUT1(8) => 
                           io_out1_2_8_port, OUT1(7) => io_out1_2_7_port, 
                           OUT1(6) => io_out1_2_6_port, OUT1(5) => 
                           io_out1_2_5_port, OUT1(4) => io_out1_2_4_port, 
                           OUT1(3) => io_out1_2_3_port, OUT1(2) => 
                           io_out1_2_2_port, OUT1(1) => io_out1_2_1_port, 
                           OUT1(0) => io_out1_2_0_port, OUT2(63) => 
                           io_out2_2_63_port, OUT2(62) => io_out2_2_62_port, 
                           OUT2(61) => io_out2_2_61_port, OUT2(60) => 
                           io_out2_2_60_port, OUT2(59) => io_out2_2_59_port, 
                           OUT2(58) => io_out2_2_58_port, OUT2(57) => 
                           io_out2_2_57_port, OUT2(56) => io_out2_2_56_port, 
                           OUT2(55) => io_out2_2_55_port, OUT2(54) => 
                           io_out2_2_54_port, OUT2(53) => io_out2_2_53_port, 
                           OUT2(52) => io_out2_2_52_port, OUT2(51) => 
                           io_out2_2_51_port, OUT2(50) => io_out2_2_50_port, 
                           OUT2(49) => io_out2_2_49_port, OUT2(48) => 
                           io_out2_2_48_port, OUT2(47) => io_out2_2_47_port, 
                           OUT2(46) => io_out2_2_46_port, OUT2(45) => 
                           io_out2_2_45_port, OUT2(44) => io_out2_2_44_port, 
                           OUT2(43) => io_out2_2_43_port, OUT2(42) => 
                           io_out2_2_42_port, OUT2(41) => io_out2_2_41_port, 
                           OUT2(40) => io_out2_2_40_port, OUT2(39) => 
                           io_out2_2_39_port, OUT2(38) => io_out2_2_38_port, 
                           OUT2(37) => io_out2_2_37_port, OUT2(36) => 
                           io_out2_2_36_port, OUT2(35) => io_out2_2_35_port, 
                           OUT2(34) => io_out2_2_34_port, OUT2(33) => 
                           io_out2_2_33_port, OUT2(32) => io_out2_2_32_port, 
                           OUT2(31) => io_out2_2_31_port, OUT2(30) => 
                           io_out2_2_30_port, OUT2(29) => io_out2_2_29_port, 
                           OUT2(28) => io_out2_2_28_port, OUT2(27) => 
                           io_out2_2_27_port, OUT2(26) => io_out2_2_26_port, 
                           OUT2(25) => io_out2_2_25_port, OUT2(24) => 
                           io_out2_2_24_port, OUT2(23) => io_out2_2_23_port, 
                           OUT2(22) => io_out2_2_22_port, OUT2(21) => 
                           io_out2_2_21_port, OUT2(20) => io_out2_2_20_port, 
                           OUT2(19) => io_out2_2_19_port, OUT2(18) => 
                           io_out2_2_18_port, OUT2(17) => io_out2_2_17_port, 
                           OUT2(16) => io_out2_2_16_port, OUT2(15) => 
                           io_out2_2_15_port, OUT2(14) => io_out2_2_14_port, 
                           OUT2(13) => io_out2_2_13_port, OUT2(12) => 
                           io_out2_2_12_port, OUT2(11) => io_out2_2_11_port, 
                           OUT2(10) => io_out2_2_10_port, OUT2(9) => 
                           io_out2_2_9_port, OUT2(8) => io_out2_2_8_port, 
                           OUT2(7) => io_out2_2_7_port, OUT2(6) => 
                           io_out2_2_6_port, OUT2(5) => io_out2_2_5_port, 
                           OUT2(4) => io_out2_2_4_port, OUT2(3) => 
                           io_out2_2_3_port, OUT2(2) => io_out2_2_2_port, 
                           OUT2(1) => io_out2_2_1_port, OUT2(0) => 
                           io_out2_2_0_port);
   loc_rf_2 : register_file_reg_size64_file_size4_3 port map( CLK => CLK, RESET
                           => RESET, ENABLE => enable_loc_2_port, RD1 => 
                           loc_read1_3_port, RD2 => loc_read2_3_port, WR => 
                           loc_write_3_port, ADD_WR(1) => ADD_WR(1), ADD_WR(0) 
                           => ADD_WR(0), ADD_RD1(1) => ADD_RD1(1), ADD_RD1(0) 
                           => ADD_RD1(0), ADD_RD2(1) => ADD_RD2(1), ADD_RD2(0) 
                           => ADD_RD2(0), DATAIN(63) => DATAIN(63), DATAIN(62) 
                           => DATAIN(62), DATAIN(61) => DATAIN(61), DATAIN(60) 
                           => DATAIN(60), DATAIN(59) => DATAIN(59), DATAIN(58) 
                           => DATAIN(58), DATAIN(57) => DATAIN(57), DATAIN(56) 
                           => DATAIN(56), DATAIN(55) => DATAIN(55), DATAIN(54) 
                           => DATAIN(54), DATAIN(53) => DATAIN(53), DATAIN(52) 
                           => DATAIN(52), DATAIN(51) => DATAIN(51), DATAIN(50) 
                           => DATAIN(50), DATAIN(49) => DATAIN(49), DATAIN(48) 
                           => DATAIN(48), DATAIN(47) => DATAIN(47), DATAIN(46) 
                           => DATAIN(46), DATAIN(45) => DATAIN(45), DATAIN(44) 
                           => DATAIN(44), DATAIN(43) => DATAIN(43), DATAIN(42) 
                           => DATAIN(42), DATAIN(41) => DATAIN(41), DATAIN(40) 
                           => DATAIN(40), DATAIN(39) => DATAIN(39), DATAIN(38) 
                           => DATAIN(38), DATAIN(37) => DATAIN(37), DATAIN(36) 
                           => DATAIN(36), DATAIN(35) => DATAIN(35), DATAIN(34) 
                           => DATAIN(34), DATAIN(33) => DATAIN(33), DATAIN(32) 
                           => DATAIN(32), DATAIN(31) => DATAIN(31), DATAIN(30) 
                           => DATAIN(30), DATAIN(29) => DATAIN(29), DATAIN(28) 
                           => DATAIN(28), DATAIN(27) => DATAIN(27), DATAIN(26) 
                           => DATAIN(26), DATAIN(25) => DATAIN(25), DATAIN(24) 
                           => DATAIN(24), DATAIN(23) => DATAIN(23), DATAIN(22) 
                           => DATAIN(22), DATAIN(21) => DATAIN(21), DATAIN(20) 
                           => DATAIN(20), DATAIN(19) => DATAIN(19), DATAIN(18) 
                           => DATAIN(18), DATAIN(17) => DATAIN(17), DATAIN(16) 
                           => DATAIN(16), DATAIN(15) => DATAIN(15), DATAIN(14) 
                           => DATAIN(14), DATAIN(13) => DATAIN(13), DATAIN(12) 
                           => DATAIN(12), DATAIN(11) => DATAIN(11), DATAIN(10) 
                           => DATAIN(10), DATAIN(9) => DATAIN(9), DATAIN(8) => 
                           DATAIN(8), DATAIN(7) => DATAIN(7), DATAIN(6) => 
                           DATAIN(6), DATAIN(5) => DATAIN(5), DATAIN(4) => 
                           DATAIN(4), DATAIN(3) => DATAIN(3), DATAIN(2) => 
                           DATAIN(2), DATAIN(1) => DATAIN(1), DATAIN(0) => 
                           DATAIN(0), OUT1(63) => loc_out1_2_63_port, OUT1(62) 
                           => loc_out1_2_62_port, OUT1(61) => 
                           loc_out1_2_61_port, OUT1(60) => loc_out1_2_60_port, 
                           OUT1(59) => loc_out1_2_59_port, OUT1(58) => 
                           loc_out1_2_58_port, OUT1(57) => loc_out1_2_57_port, 
                           OUT1(56) => loc_out1_2_56_port, OUT1(55) => 
                           loc_out1_2_55_port, OUT1(54) => loc_out1_2_54_port, 
                           OUT1(53) => loc_out1_2_53_port, OUT1(52) => 
                           loc_out1_2_52_port, OUT1(51) => loc_out1_2_51_port, 
                           OUT1(50) => loc_out1_2_50_port, OUT1(49) => 
                           loc_out1_2_49_port, OUT1(48) => loc_out1_2_48_port, 
                           OUT1(47) => loc_out1_2_47_port, OUT1(46) => 
                           loc_out1_2_46_port, OUT1(45) => loc_out1_2_45_port, 
                           OUT1(44) => loc_out1_2_44_port, OUT1(43) => 
                           loc_out1_2_43_port, OUT1(42) => loc_out1_2_42_port, 
                           OUT1(41) => loc_out1_2_41_port, OUT1(40) => 
                           loc_out1_2_40_port, OUT1(39) => loc_out1_2_39_port, 
                           OUT1(38) => loc_out1_2_38_port, OUT1(37) => 
                           loc_out1_2_37_port, OUT1(36) => loc_out1_2_36_port, 
                           OUT1(35) => loc_out1_2_35_port, OUT1(34) => 
                           loc_out1_2_34_port, OUT1(33) => loc_out1_2_33_port, 
                           OUT1(32) => loc_out1_2_32_port, OUT1(31) => 
                           loc_out1_2_31_port, OUT1(30) => loc_out1_2_30_port, 
                           OUT1(29) => loc_out1_2_29_port, OUT1(28) => 
                           loc_out1_2_28_port, OUT1(27) => loc_out1_2_27_port, 
                           OUT1(26) => loc_out1_2_26_port, OUT1(25) => 
                           loc_out1_2_25_port, OUT1(24) => loc_out1_2_24_port, 
                           OUT1(23) => loc_out1_2_23_port, OUT1(22) => 
                           loc_out1_2_22_port, OUT1(21) => loc_out1_2_21_port, 
                           OUT1(20) => loc_out1_2_20_port, OUT1(19) => 
                           loc_out1_2_19_port, OUT1(18) => loc_out1_2_18_port, 
                           OUT1(17) => loc_out1_2_17_port, OUT1(16) => 
                           loc_out1_2_16_port, OUT1(15) => loc_out1_2_15_port, 
                           OUT1(14) => loc_out1_2_14_port, OUT1(13) => 
                           loc_out1_2_13_port, OUT1(12) => loc_out1_2_12_port, 
                           OUT1(11) => loc_out1_2_11_port, OUT1(10) => 
                           loc_out1_2_10_port, OUT1(9) => loc_out1_2_9_port, 
                           OUT1(8) => loc_out1_2_8_port, OUT1(7) => 
                           loc_out1_2_7_port, OUT1(6) => loc_out1_2_6_port, 
                           OUT1(5) => loc_out1_2_5_port, OUT1(4) => 
                           loc_out1_2_4_port, OUT1(3) => loc_out1_2_3_port, 
                           OUT1(2) => loc_out1_2_2_port, OUT1(1) => 
                           loc_out1_2_1_port, OUT1(0) => loc_out1_2_0_port, 
                           OUT2(63) => loc_out2_2_63_port, OUT2(62) => 
                           loc_out2_2_62_port, OUT2(61) => loc_out2_2_61_port, 
                           OUT2(60) => loc_out2_2_60_port, OUT2(59) => 
                           loc_out2_2_59_port, OUT2(58) => loc_out2_2_58_port, 
                           OUT2(57) => loc_out2_2_57_port, OUT2(56) => 
                           loc_out2_2_56_port, OUT2(55) => loc_out2_2_55_port, 
                           OUT2(54) => loc_out2_2_54_port, OUT2(53) => 
                           loc_out2_2_53_port, OUT2(52) => loc_out2_2_52_port, 
                           OUT2(51) => loc_out2_2_51_port, OUT2(50) => 
                           loc_out2_2_50_port, OUT2(49) => loc_out2_2_49_port, 
                           OUT2(48) => loc_out2_2_48_port, OUT2(47) => 
                           loc_out2_2_47_port, OUT2(46) => loc_out2_2_46_port, 
                           OUT2(45) => loc_out2_2_45_port, OUT2(44) => 
                           loc_out2_2_44_port, OUT2(43) => loc_out2_2_43_port, 
                           OUT2(42) => loc_out2_2_42_port, OUT2(41) => 
                           loc_out2_2_41_port, OUT2(40) => loc_out2_2_40_port, 
                           OUT2(39) => loc_out2_2_39_port, OUT2(38) => 
                           loc_out2_2_38_port, OUT2(37) => loc_out2_2_37_port, 
                           OUT2(36) => loc_out2_2_36_port, OUT2(35) => 
                           loc_out2_2_35_port, OUT2(34) => loc_out2_2_34_port, 
                           OUT2(33) => loc_out2_2_33_port, OUT2(32) => 
                           loc_out2_2_32_port, OUT2(31) => loc_out2_2_31_port, 
                           OUT2(30) => loc_out2_2_30_port, OUT2(29) => 
                           loc_out2_2_29_port, OUT2(28) => loc_out2_2_28_port, 
                           OUT2(27) => loc_out2_2_27_port, OUT2(26) => 
                           loc_out2_2_26_port, OUT2(25) => loc_out2_2_25_port, 
                           OUT2(24) => loc_out2_2_24_port, OUT2(23) => 
                           loc_out2_2_23_port, OUT2(22) => loc_out2_2_22_port, 
                           OUT2(21) => loc_out2_2_21_port, OUT2(20) => 
                           loc_out2_2_20_port, OUT2(19) => loc_out2_2_19_port, 
                           OUT2(18) => loc_out2_2_18_port, OUT2(17) => 
                           loc_out2_2_17_port, OUT2(16) => loc_out2_2_16_port, 
                           OUT2(15) => loc_out2_2_15_port, OUT2(14) => 
                           loc_out2_2_14_port, OUT2(13) => loc_out2_2_13_port, 
                           OUT2(12) => loc_out2_2_12_port, OUT2(11) => 
                           loc_out2_2_11_port, OUT2(10) => loc_out2_2_10_port, 
                           OUT2(9) => loc_out2_2_9_port, OUT2(8) => 
                           loc_out2_2_8_port, OUT2(7) => loc_out2_2_7_port, 
                           OUT2(6) => loc_out2_2_6_port, OUT2(5) => 
                           loc_out2_2_5_port, OUT2(4) => loc_out2_2_4_port, 
                           OUT2(3) => loc_out2_2_3_port, OUT2(2) => 
                           loc_out2_2_2_port, OUT2(1) => loc_out2_2_1_port, 
                           OUT2(0) => loc_out2_2_0_port);
   io_rf_3 : register_file_reg_size64_file_size4_2 port map( CLK => CLK, RESET 
                           => RESET, ENABLE => enable_io_3_port, RD1 => 
                           io_read1_3_port, RD2 => io_read2_3_port, WR => 
                           io_write_3_port, ADD_WR(1) => ADD_WR(1), ADD_WR(0) 
                           => ADD_WR(0), ADD_RD1(1) => ADD_RD1(1), ADD_RD1(0) 
                           => ADD_RD1(0), ADD_RD2(1) => ADD_RD2(1), ADD_RD2(0) 
                           => ADD_RD2(0), DATAIN(63) => DATAIN(63), DATAIN(62) 
                           => DATAIN(62), DATAIN(61) => DATAIN(61), DATAIN(60) 
                           => DATAIN(60), DATAIN(59) => DATAIN(59), DATAIN(58) 
                           => DATAIN(58), DATAIN(57) => DATAIN(57), DATAIN(56) 
                           => DATAIN(56), DATAIN(55) => DATAIN(55), DATAIN(54) 
                           => DATAIN(54), DATAIN(53) => DATAIN(53), DATAIN(52) 
                           => DATAIN(52), DATAIN(51) => DATAIN(51), DATAIN(50) 
                           => DATAIN(50), DATAIN(49) => DATAIN(49), DATAIN(48) 
                           => DATAIN(48), DATAIN(47) => DATAIN(47), DATAIN(46) 
                           => DATAIN(46), DATAIN(45) => DATAIN(45), DATAIN(44) 
                           => DATAIN(44), DATAIN(43) => DATAIN(43), DATAIN(42) 
                           => DATAIN(42), DATAIN(41) => DATAIN(41), DATAIN(40) 
                           => DATAIN(40), DATAIN(39) => DATAIN(39), DATAIN(38) 
                           => DATAIN(38), DATAIN(37) => DATAIN(37), DATAIN(36) 
                           => DATAIN(36), DATAIN(35) => DATAIN(35), DATAIN(34) 
                           => DATAIN(34), DATAIN(33) => DATAIN(33), DATAIN(32) 
                           => DATAIN(32), DATAIN(31) => DATAIN(31), DATAIN(30) 
                           => DATAIN(30), DATAIN(29) => DATAIN(29), DATAIN(28) 
                           => DATAIN(28), DATAIN(27) => DATAIN(27), DATAIN(26) 
                           => DATAIN(26), DATAIN(25) => DATAIN(25), DATAIN(24) 
                           => DATAIN(24), DATAIN(23) => DATAIN(23), DATAIN(22) 
                           => DATAIN(22), DATAIN(21) => DATAIN(21), DATAIN(20) 
                           => DATAIN(20), DATAIN(19) => DATAIN(19), DATAIN(18) 
                           => DATAIN(18), DATAIN(17) => DATAIN(17), DATAIN(16) 
                           => DATAIN(16), DATAIN(15) => DATAIN(15), DATAIN(14) 
                           => DATAIN(14), DATAIN(13) => DATAIN(13), DATAIN(12) 
                           => DATAIN(12), DATAIN(11) => DATAIN(11), DATAIN(10) 
                           => DATAIN(10), DATAIN(9) => DATAIN(9), DATAIN(8) => 
                           DATAIN(8), DATAIN(7) => DATAIN(7), DATAIN(6) => 
                           DATAIN(6), DATAIN(5) => DATAIN(5), DATAIN(4) => 
                           DATAIN(4), DATAIN(3) => DATAIN(3), DATAIN(2) => 
                           DATAIN(2), DATAIN(1) => DATAIN(1), DATAIN(0) => 
                           DATAIN(0), OUT1(63) => io_out1_3_63_port, OUT1(62) 
                           => io_out1_3_62_port, OUT1(61) => io_out1_3_61_port,
                           OUT1(60) => io_out1_3_60_port, OUT1(59) => 
                           io_out1_3_59_port, OUT1(58) => io_out1_3_58_port, 
                           OUT1(57) => io_out1_3_57_port, OUT1(56) => 
                           io_out1_3_56_port, OUT1(55) => io_out1_3_55_port, 
                           OUT1(54) => io_out1_3_54_port, OUT1(53) => 
                           io_out1_3_53_port, OUT1(52) => io_out1_3_52_port, 
                           OUT1(51) => io_out1_3_51_port, OUT1(50) => 
                           io_out1_3_50_port, OUT1(49) => io_out1_3_49_port, 
                           OUT1(48) => io_out1_3_48_port, OUT1(47) => 
                           io_out1_3_47_port, OUT1(46) => io_out1_3_46_port, 
                           OUT1(45) => io_out1_3_45_port, OUT1(44) => 
                           io_out1_3_44_port, OUT1(43) => io_out1_3_43_port, 
                           OUT1(42) => io_out1_3_42_port, OUT1(41) => 
                           io_out1_3_41_port, OUT1(40) => io_out1_3_40_port, 
                           OUT1(39) => io_out1_3_39_port, OUT1(38) => 
                           io_out1_3_38_port, OUT1(37) => io_out1_3_37_port, 
                           OUT1(36) => io_out1_3_36_port, OUT1(35) => 
                           io_out1_3_35_port, OUT1(34) => io_out1_3_34_port, 
                           OUT1(33) => io_out1_3_33_port, OUT1(32) => 
                           io_out1_3_32_port, OUT1(31) => io_out1_3_31_port, 
                           OUT1(30) => io_out1_3_30_port, OUT1(29) => 
                           io_out1_3_29_port, OUT1(28) => io_out1_3_28_port, 
                           OUT1(27) => io_out1_3_27_port, OUT1(26) => 
                           io_out1_3_26_port, OUT1(25) => io_out1_3_25_port, 
                           OUT1(24) => io_out1_3_24_port, OUT1(23) => 
                           io_out1_3_23_port, OUT1(22) => io_out1_3_22_port, 
                           OUT1(21) => io_out1_3_21_port, OUT1(20) => 
                           io_out1_3_20_port, OUT1(19) => io_out1_3_19_port, 
                           OUT1(18) => io_out1_3_18_port, OUT1(17) => 
                           io_out1_3_17_port, OUT1(16) => io_out1_3_16_port, 
                           OUT1(15) => io_out1_3_15_port, OUT1(14) => 
                           io_out1_3_14_port, OUT1(13) => io_out1_3_13_port, 
                           OUT1(12) => io_out1_3_12_port, OUT1(11) => 
                           io_out1_3_11_port, OUT1(10) => io_out1_3_10_port, 
                           OUT1(9) => io_out1_3_9_port, OUT1(8) => 
                           io_out1_3_8_port, OUT1(7) => io_out1_3_7_port, 
                           OUT1(6) => io_out1_3_6_port, OUT1(5) => 
                           io_out1_3_5_port, OUT1(4) => io_out1_3_4_port, 
                           OUT1(3) => io_out1_3_3_port, OUT1(2) => 
                           io_out1_3_2_port, OUT1(1) => io_out1_3_1_port, 
                           OUT1(0) => io_out1_3_0_port, OUT2(63) => 
                           io_out2_3_63_port, OUT2(62) => io_out2_3_62_port, 
                           OUT2(61) => io_out2_3_61_port, OUT2(60) => 
                           io_out2_3_60_port, OUT2(59) => io_out2_3_59_port, 
                           OUT2(58) => io_out2_3_58_port, OUT2(57) => 
                           io_out2_3_57_port, OUT2(56) => io_out2_3_56_port, 
                           OUT2(55) => io_out2_3_55_port, OUT2(54) => 
                           io_out2_3_54_port, OUT2(53) => io_out2_3_53_port, 
                           OUT2(52) => io_out2_3_52_port, OUT2(51) => 
                           io_out2_3_51_port, OUT2(50) => io_out2_3_50_port, 
                           OUT2(49) => io_out2_3_49_port, OUT2(48) => 
                           io_out2_3_48_port, OUT2(47) => io_out2_3_47_port, 
                           OUT2(46) => io_out2_3_46_port, OUT2(45) => 
                           io_out2_3_45_port, OUT2(44) => io_out2_3_44_port, 
                           OUT2(43) => io_out2_3_43_port, OUT2(42) => 
                           io_out2_3_42_port, OUT2(41) => io_out2_3_41_port, 
                           OUT2(40) => io_out2_3_40_port, OUT2(39) => 
                           io_out2_3_39_port, OUT2(38) => io_out2_3_38_port, 
                           OUT2(37) => io_out2_3_37_port, OUT2(36) => 
                           io_out2_3_36_port, OUT2(35) => io_out2_3_35_port, 
                           OUT2(34) => io_out2_3_34_port, OUT2(33) => 
                           io_out2_3_33_port, OUT2(32) => io_out2_3_32_port, 
                           OUT2(31) => io_out2_3_31_port, OUT2(30) => 
                           io_out2_3_30_port, OUT2(29) => io_out2_3_29_port, 
                           OUT2(28) => io_out2_3_28_port, OUT2(27) => 
                           io_out2_3_27_port, OUT2(26) => io_out2_3_26_port, 
                           OUT2(25) => io_out2_3_25_port, OUT2(24) => 
                           io_out2_3_24_port, OUT2(23) => io_out2_3_23_port, 
                           OUT2(22) => io_out2_3_22_port, OUT2(21) => 
                           io_out2_3_21_port, OUT2(20) => io_out2_3_20_port, 
                           OUT2(19) => io_out2_3_19_port, OUT2(18) => 
                           io_out2_3_18_port, OUT2(17) => io_out2_3_17_port, 
                           OUT2(16) => io_out2_3_16_port, OUT2(15) => 
                           io_out2_3_15_port, OUT2(14) => io_out2_3_14_port, 
                           OUT2(13) => io_out2_3_13_port, OUT2(12) => 
                           io_out2_3_12_port, OUT2(11) => io_out2_3_11_port, 
                           OUT2(10) => io_out2_3_10_port, OUT2(9) => 
                           io_out2_3_9_port, OUT2(8) => io_out2_3_8_port, 
                           OUT2(7) => io_out2_3_7_port, OUT2(6) => 
                           io_out2_3_6_port, OUT2(5) => io_out2_3_5_port, 
                           OUT2(4) => io_out2_3_4_port, OUT2(3) => 
                           io_out2_3_3_port, OUT2(2) => io_out2_3_2_port, 
                           OUT2(1) => io_out2_3_1_port, OUT2(0) => 
                           io_out2_3_0_port);
   loc_rf_3 : register_file_reg_size64_file_size4_1 port map( CLK => CLK, RESET
                           => RESET, ENABLE => enable_loc_3_port, RD1 => 
                           loc_read1_3_port, RD2 => loc_read2_3_port, WR => 
                           loc_write_3_port, ADD_WR(1) => ADD_WR(1), ADD_WR(0) 
                           => ADD_WR(0), ADD_RD1(1) => ADD_RD1(1), ADD_RD1(0) 
                           => ADD_RD1(0), ADD_RD2(1) => ADD_RD2(1), ADD_RD2(0) 
                           => ADD_RD2(0), DATAIN(63) => DATAIN(63), DATAIN(62) 
                           => DATAIN(62), DATAIN(61) => DATAIN(61), DATAIN(60) 
                           => DATAIN(60), DATAIN(59) => DATAIN(59), DATAIN(58) 
                           => DATAIN(58), DATAIN(57) => DATAIN(57), DATAIN(56) 
                           => DATAIN(56), DATAIN(55) => DATAIN(55), DATAIN(54) 
                           => DATAIN(54), DATAIN(53) => DATAIN(53), DATAIN(52) 
                           => DATAIN(52), DATAIN(51) => DATAIN(51), DATAIN(50) 
                           => DATAIN(50), DATAIN(49) => DATAIN(49), DATAIN(48) 
                           => DATAIN(48), DATAIN(47) => DATAIN(47), DATAIN(46) 
                           => DATAIN(46), DATAIN(45) => DATAIN(45), DATAIN(44) 
                           => DATAIN(44), DATAIN(43) => DATAIN(43), DATAIN(42) 
                           => DATAIN(42), DATAIN(41) => DATAIN(41), DATAIN(40) 
                           => DATAIN(40), DATAIN(39) => DATAIN(39), DATAIN(38) 
                           => DATAIN(38), DATAIN(37) => DATAIN(37), DATAIN(36) 
                           => DATAIN(36), DATAIN(35) => DATAIN(35), DATAIN(34) 
                           => DATAIN(34), DATAIN(33) => DATAIN(33), DATAIN(32) 
                           => DATAIN(32), DATAIN(31) => DATAIN(31), DATAIN(30) 
                           => DATAIN(30), DATAIN(29) => DATAIN(29), DATAIN(28) 
                           => DATAIN(28), DATAIN(27) => DATAIN(27), DATAIN(26) 
                           => DATAIN(26), DATAIN(25) => DATAIN(25), DATAIN(24) 
                           => DATAIN(24), DATAIN(23) => DATAIN(23), DATAIN(22) 
                           => DATAIN(22), DATAIN(21) => DATAIN(21), DATAIN(20) 
                           => DATAIN(20), DATAIN(19) => DATAIN(19), DATAIN(18) 
                           => DATAIN(18), DATAIN(17) => DATAIN(17), DATAIN(16) 
                           => DATAIN(16), DATAIN(15) => DATAIN(15), DATAIN(14) 
                           => DATAIN(14), DATAIN(13) => DATAIN(13), DATAIN(12) 
                           => DATAIN(12), DATAIN(11) => DATAIN(11), DATAIN(10) 
                           => DATAIN(10), DATAIN(9) => DATAIN(9), DATAIN(8) => 
                           DATAIN(8), DATAIN(7) => DATAIN(7), DATAIN(6) => 
                           DATAIN(6), DATAIN(5) => DATAIN(5), DATAIN(4) => 
                           DATAIN(4), DATAIN(3) => DATAIN(3), DATAIN(2) => 
                           DATAIN(2), DATAIN(1) => DATAIN(1), DATAIN(0) => 
                           DATAIN(0), OUT1(63) => loc_out1_3_63_port, OUT1(62) 
                           => loc_out1_3_62_port, OUT1(61) => 
                           loc_out1_3_61_port, OUT1(60) => loc_out1_3_60_port, 
                           OUT1(59) => loc_out1_3_59_port, OUT1(58) => 
                           loc_out1_3_58_port, OUT1(57) => loc_out1_3_57_port, 
                           OUT1(56) => loc_out1_3_56_port, OUT1(55) => 
                           loc_out1_3_55_port, OUT1(54) => loc_out1_3_54_port, 
                           OUT1(53) => loc_out1_3_53_port, OUT1(52) => 
                           loc_out1_3_52_port, OUT1(51) => loc_out1_3_51_port, 
                           OUT1(50) => loc_out1_3_50_port, OUT1(49) => 
                           loc_out1_3_49_port, OUT1(48) => loc_out1_3_48_port, 
                           OUT1(47) => loc_out1_3_47_port, OUT1(46) => 
                           loc_out1_3_46_port, OUT1(45) => loc_out1_3_45_port, 
                           OUT1(44) => loc_out1_3_44_port, OUT1(43) => 
                           loc_out1_3_43_port, OUT1(42) => loc_out1_3_42_port, 
                           OUT1(41) => loc_out1_3_41_port, OUT1(40) => 
                           loc_out1_3_40_port, OUT1(39) => loc_out1_3_39_port, 
                           OUT1(38) => loc_out1_3_38_port, OUT1(37) => 
                           loc_out1_3_37_port, OUT1(36) => loc_out1_3_36_port, 
                           OUT1(35) => loc_out1_3_35_port, OUT1(34) => 
                           loc_out1_3_34_port, OUT1(33) => loc_out1_3_33_port, 
                           OUT1(32) => loc_out1_3_32_port, OUT1(31) => 
                           loc_out1_3_31_port, OUT1(30) => loc_out1_3_30_port, 
                           OUT1(29) => loc_out1_3_29_port, OUT1(28) => 
                           loc_out1_3_28_port, OUT1(27) => loc_out1_3_27_port, 
                           OUT1(26) => loc_out1_3_26_port, OUT1(25) => 
                           loc_out1_3_25_port, OUT1(24) => loc_out1_3_24_port, 
                           OUT1(23) => loc_out1_3_23_port, OUT1(22) => 
                           loc_out1_3_22_port, OUT1(21) => loc_out1_3_21_port, 
                           OUT1(20) => loc_out1_3_20_port, OUT1(19) => 
                           loc_out1_3_19_port, OUT1(18) => loc_out1_3_18_port, 
                           OUT1(17) => loc_out1_3_17_port, OUT1(16) => 
                           loc_out1_3_16_port, OUT1(15) => loc_out1_3_15_port, 
                           OUT1(14) => loc_out1_3_14_port, OUT1(13) => 
                           loc_out1_3_13_port, OUT1(12) => loc_out1_3_12_port, 
                           OUT1(11) => loc_out1_3_11_port, OUT1(10) => 
                           loc_out1_3_10_port, OUT1(9) => loc_out1_3_9_port, 
                           OUT1(8) => loc_out1_3_8_port, OUT1(7) => 
                           loc_out1_3_7_port, OUT1(6) => loc_out1_3_6_port, 
                           OUT1(5) => loc_out1_3_5_port, OUT1(4) => 
                           loc_out1_3_4_port, OUT1(3) => loc_out1_3_3_port, 
                           OUT1(2) => loc_out1_3_2_port, OUT1(1) => 
                           loc_out1_3_1_port, OUT1(0) => loc_out1_3_0_port, 
                           OUT2(63) => loc_out2_3_63_port, OUT2(62) => 
                           loc_out2_3_62_port, OUT2(61) => loc_out2_3_61_port, 
                           OUT2(60) => loc_out2_3_60_port, OUT2(59) => 
                           loc_out2_3_59_port, OUT2(58) => loc_out2_3_58_port, 
                           OUT2(57) => loc_out2_3_57_port, OUT2(56) => 
                           loc_out2_3_56_port, OUT2(55) => loc_out2_3_55_port, 
                           OUT2(54) => loc_out2_3_54_port, OUT2(53) => 
                           loc_out2_3_53_port, OUT2(52) => loc_out2_3_52_port, 
                           OUT2(51) => loc_out2_3_51_port, OUT2(50) => 
                           loc_out2_3_50_port, OUT2(49) => loc_out2_3_49_port, 
                           OUT2(48) => loc_out2_3_48_port, OUT2(47) => 
                           loc_out2_3_47_port, OUT2(46) => loc_out2_3_46_port, 
                           OUT2(45) => loc_out2_3_45_port, OUT2(44) => 
                           loc_out2_3_44_port, OUT2(43) => loc_out2_3_43_port, 
                           OUT2(42) => loc_out2_3_42_port, OUT2(41) => 
                           loc_out2_3_41_port, OUT2(40) => loc_out2_3_40_port, 
                           OUT2(39) => loc_out2_3_39_port, OUT2(38) => 
                           loc_out2_3_38_port, OUT2(37) => loc_out2_3_37_port, 
                           OUT2(36) => loc_out2_3_36_port, OUT2(35) => 
                           loc_out2_3_35_port, OUT2(34) => loc_out2_3_34_port, 
                           OUT2(33) => loc_out2_3_33_port, OUT2(32) => 
                           loc_out2_3_32_port, OUT2(31) => loc_out2_3_31_port, 
                           OUT2(30) => loc_out2_3_30_port, OUT2(29) => 
                           loc_out2_3_29_port, OUT2(28) => loc_out2_3_28_port, 
                           OUT2(27) => loc_out2_3_27_port, OUT2(26) => 
                           loc_out2_3_26_port, OUT2(25) => loc_out2_3_25_port, 
                           OUT2(24) => loc_out2_3_24_port, OUT2(23) => 
                           loc_out2_3_23_port, OUT2(22) => loc_out2_3_22_port, 
                           OUT2(21) => loc_out2_3_21_port, OUT2(20) => 
                           loc_out2_3_20_port, OUT2(19) => loc_out2_3_19_port, 
                           OUT2(18) => loc_out2_3_18_port, OUT2(17) => 
                           loc_out2_3_17_port, OUT2(16) => loc_out2_3_16_port, 
                           OUT2(15) => loc_out2_3_15_port, OUT2(14) => 
                           loc_out2_3_14_port, OUT2(13) => loc_out2_3_13_port, 
                           OUT2(12) => loc_out2_3_12_port, OUT2(11) => 
                           loc_out2_3_11_port, OUT2(10) => loc_out2_3_10_port, 
                           OUT2(9) => loc_out2_3_9_port, OUT2(8) => 
                           loc_out2_3_8_port, OUT2(7) => loc_out2_3_7_port, 
                           OUT2(6) => loc_out2_3_6_port, OUT2(5) => 
                           loc_out2_3_5_port, OUT2(4) => loc_out2_3_4_port, 
                           OUT2(3) => loc_out2_3_3_port, OUT2(2) => 
                           loc_out2_3_2_port, OUT2(1) => loc_out2_3_1_port, 
                           OUT2(0) => loc_out2_3_0_port);
   OUT2_reg_63_inst : DLH_X1 port map( G => n3077, D => N1195, Q => OUT2(63));
   OUT2_reg_62_inst : DLH_X1 port map( G => n3075, D => N1194, Q => OUT2(62));
   OUT2_reg_61_inst : DLH_X1 port map( G => n3075, D => N1193, Q => OUT2(61));
   OUT2_reg_60_inst : DLH_X1 port map( G => n3075, D => N1192, Q => OUT2(60));
   OUT2_reg_59_inst : DLH_X1 port map( G => n3075, D => N1191, Q => OUT2(59));
   OUT2_reg_58_inst : DLH_X1 port map( G => n3075, D => N1190, Q => OUT2(58));
   OUT2_reg_57_inst : DLH_X1 port map( G => n3075, D => N1189, Q => OUT2(57));
   OUT2_reg_56_inst : DLH_X1 port map( G => n3075, D => N1188, Q => OUT2(56));
   OUT2_reg_55_inst : DLH_X1 port map( G => n3075, D => N1187, Q => OUT2(55));
   OUT2_reg_54_inst : DLH_X1 port map( G => n3075, D => N1186, Q => OUT2(54));
   OUT2_reg_53_inst : DLH_X1 port map( G => n3075, D => N1185, Q => OUT2(53));
   OUT2_reg_52_inst : DLH_X1 port map( G => n3076, D => N1184, Q => OUT2(52));
   OUT2_reg_51_inst : DLH_X1 port map( G => n3076, D => N1183, Q => OUT2(51));
   OUT2_reg_50_inst : DLH_X1 port map( G => n3076, D => N1182, Q => OUT2(50));
   OUT2_reg_49_inst : DLH_X1 port map( G => n3076, D => N1181, Q => OUT2(49));
   OUT2_reg_48_inst : DLH_X1 port map( G => n3076, D => N1180, Q => OUT2(48));
   OUT2_reg_47_inst : DLH_X1 port map( G => n3076, D => N1179, Q => OUT2(47));
   OUT2_reg_46_inst : DLH_X1 port map( G => n3076, D => N1178, Q => OUT2(46));
   OUT2_reg_45_inst : DLH_X1 port map( G => n3076, D => N1177, Q => OUT2(45));
   OUT2_reg_44_inst : DLH_X1 port map( G => n3076, D => N1176, Q => OUT2(44));
   OUT2_reg_43_inst : DLH_X1 port map( G => n3076, D => N1175, Q => OUT2(43));
   OUT2_reg_42_inst : DLH_X1 port map( G => n3076, D => N1174, Q => OUT2(42));
   OUT2_reg_41_inst : DLH_X1 port map( G => n3076, D => N1173, Q => OUT2(41));
   OUT2_reg_40_inst : DLH_X1 port map( G => n3077, D => N1172, Q => OUT2(40));
   OUT2_reg_39_inst : DLH_X1 port map( G => n3077, D => N1171, Q => OUT2(39));
   OUT2_reg_38_inst : DLH_X1 port map( G => n3077, D => N1170, Q => OUT2(38));
   OUT2_reg_37_inst : DLH_X1 port map( G => n3077, D => N1169, Q => OUT2(37));
   OUT2_reg_36_inst : DLH_X1 port map( G => n3077, D => N1168, Q => OUT2(36));
   OUT2_reg_35_inst : DLH_X1 port map( G => n3077, D => N1167, Q => OUT2(35));
   OUT2_reg_34_inst : DLH_X1 port map( G => n3077, D => N1166, Q => OUT2(34));
   OUT2_reg_33_inst : DLH_X1 port map( G => n3077, D => N1165, Q => OUT2(33));
   OUT2_reg_32_inst : DLH_X1 port map( G => n3077, D => N1164, Q => OUT2(32));
   OUT2_reg_31_inst : DLH_X1 port map( G => n3077, D => N1163, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => n3077, D => N1162, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => n3078, D => N1161, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => n3078, D => N1160, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => n3078, D => N1159, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => n3078, D => N1158, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => n3078, D => N1157, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => n3078, D => N1156, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => n3078, D => N1155, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => n3078, D => N1154, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => n3078, D => N1153, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => n3078, D => N1152, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => n3078, D => N1151, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => n3078, D => N1150, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => n3079, D => N1149, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => n3079, D => N1148, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => n3079, D => N1147, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => n3079, D => N1146, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => n3079, D => N1145, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => n3079, D => N1144, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => n3079, D => N1143, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => n3079, D => N1142, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => n3079, D => N1141, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => n3079, D => N1140, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => n3079, D => N1139, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => n3079, D => N1138, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => n3080, D => N1137, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => n3080, D => N1136, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => n3080, D => N1135, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => n3080, D => N1134, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => n3080, D => N1133, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => n3075, D => N1132, Q => OUT2(0));
   U2159 : NAND3_X1 port map( A1 => n1038, A2 => n2123, A3 => ADD_RD2(2), ZN =>
                           n2122);
   U2160 : NAND3_X1 port map( A1 => n2128, A2 => n2129, A3 => n3075, ZN => 
                           n2661);
   U2161 : NAND3_X1 port map( A1 => n2108, A2 => n2103, A3 => n2935, ZN => 
                           n2934);
   U2162 : NAND3_X1 port map( A1 => n1038, A2 => n2108, A3 => n2935, ZN => 
                           n2936);
   CWP_reg_0_inst : DFF_X1 port map( D => n1036, CK => CLK, Q => n1038, QN => 
                           n2103);
   CWP_reg_1_inst : DFF_X1 port map( D => n1035, CK => CLK, Q => n2937, QN => 
                           n2109);
   U2163 : NOR3_X1 port map( A1 => n2103, A2 => n2133, A3 => n2667, ZN => n2152
                           );
   U2164 : NOR3_X1 port map( A1 => n2133, A2 => n1038, A3 => n2667, ZN => n2155
                           );
   U2165 : BUF_X1 port map( A => n3064, Z => n3066);
   U2166 : BUF_X1 port map( A => n3065, Z => n3069);
   U2167 : BUF_X1 port map( A => n3064, Z => n3068);
   U2168 : BUF_X1 port map( A => n3064, Z => n3067);
   U2169 : BUF_X1 port map( A => n3065, Z => n3070);
   U2170 : BUF_X1 port map( A => n2139, Z => n3064);
   U2171 : BUF_X1 port map( A => n2139, Z => n3065);
   U2172 : BUF_X1 port map( A => n2157, Z => n3007);
   U2173 : BUF_X1 port map( A => n2157, Z => n3008);
   U2174 : BUF_X1 port map( A => n2157, Z => n3004);
   U2175 : BUF_X1 port map( A => n2157, Z => n3005);
   U2176 : BUF_X1 port map( A => n2157, Z => n3006);
   U2177 : INV_X1 port map( A => n2657, ZN => n2139);
   U2178 : INV_X1 port map( A => n2108, ZN => n2133);
   U2179 : INV_X1 port map( A => n3074, ZN => n3073);
   U2180 : INV_X1 port map( A => n3074, ZN => n3072);
   U2181 : INV_X1 port map( A => n3074, ZN => n3071);
   U2182 : NOR2_X1 port map( A1 => n2134, A2 => n2667, ZN => n2157);
   U2183 : BUF_X1 port map( A => n2159, Z => n2995);
   U2184 : BUF_X1 port map( A => n2159, Z => n2996);
   U2185 : BUF_X1 port map( A => n2147, Z => n3044);
   U2186 : BUF_X1 port map( A => n2147, Z => n3043);
   U2187 : BUF_X1 port map( A => n2160, Z => n2989);
   U2188 : BUF_X1 port map( A => n2160, Z => n2990);
   U2189 : BUF_X1 port map( A => n2156, Z => n3013);
   U2190 : BUF_X1 port map( A => n2156, Z => n3014);
   U2191 : BUF_X1 port map( A => n2158, Z => n3001);
   U2192 : BUF_X1 port map( A => n2158, Z => n3002);
   U2193 : BUF_X1 port map( A => n2143, Z => n3062);
   U2194 : BUF_X1 port map( A => n2143, Z => n3061);
   U2195 : BUF_X1 port map( A => n2153, Z => n3031);
   U2196 : BUF_X1 port map( A => n2153, Z => n3032);
   U2197 : BUF_X1 port map( A => n2144, Z => n3054);
   U2198 : BUF_X1 port map( A => n2144, Z => n3055);
   U2199 : BUF_X1 port map( A => n2144, Z => n3056);
   U2200 : BUF_X1 port map( A => n2154, Z => n3023);
   U2201 : BUF_X1 port map( A => n2154, Z => n3024);
   U2202 : BUF_X1 port map( A => n2154, Z => n3025);
   U2203 : BUF_X1 port map( A => n2154, Z => n3026);
   U2204 : BUF_X1 port map( A => n2152, Z => n3038);
   U2205 : BUF_X1 port map( A => n2145, Z => n3050);
   U2206 : BUF_X1 port map( A => n2159, Z => n2992);
   U2207 : BUF_X1 port map( A => n2159, Z => n2993);
   U2208 : BUF_X1 port map( A => n2159, Z => n2994);
   U2209 : BUF_X1 port map( A => n2147, Z => n3042);
   U2210 : BUF_X1 port map( A => n2147, Z => n3041);
   U2211 : BUF_X1 port map( A => n2147, Z => n3040);
   U2212 : BUF_X1 port map( A => n2156, Z => n3010);
   U2213 : BUF_X1 port map( A => n2160, Z => n2986);
   U2214 : BUF_X1 port map( A => n2158, Z => n2998);
   U2215 : BUF_X1 port map( A => n2156, Z => n3011);
   U2216 : BUF_X1 port map( A => n2160, Z => n2987);
   U2217 : BUF_X1 port map( A => n2158, Z => n2999);
   U2218 : BUF_X1 port map( A => n2156, Z => n3012);
   U2219 : BUF_X1 port map( A => n2160, Z => n2988);
   U2220 : BUF_X1 port map( A => n2158, Z => n3000);
   U2221 : BUF_X1 port map( A => n2143, Z => n3060);
   U2222 : BUF_X1 port map( A => n2143, Z => n3059);
   U2223 : BUF_X1 port map( A => n2143, Z => n3058);
   U2224 : BUF_X1 port map( A => n2153, Z => n3028);
   U2225 : BUF_X1 port map( A => n2153, Z => n3029);
   U2226 : BUF_X1 port map( A => n2153, Z => n3030);
   U2227 : BUF_X1 port map( A => n2144, Z => n3052);
   U2228 : BUF_X1 port map( A => n2144, Z => n3053);
   U2229 : BUF_X1 port map( A => n2154, Z => n3022);
   U2230 : BUF_X1 port map( A => n2152, Z => n3034);
   U2231 : BUF_X1 port map( A => n2152, Z => n3035);
   U2232 : BUF_X1 port map( A => n2152, Z => n3036);
   U2233 : BUF_X1 port map( A => n2152, Z => n3037);
   U2234 : BUF_X1 port map( A => n2145, Z => n3046);
   U2235 : BUF_X1 port map( A => n2145, Z => n3047);
   U2236 : BUF_X1 port map( A => n2145, Z => n3048);
   U2237 : BUF_X1 port map( A => n2145, Z => n3049);
   U2238 : NOR2_X1 port map( A1 => n2661, A2 => n2136, ZN => n2657);
   U2239 : BUF_X1 port map( A => n2672, Z => n2983);
   U2240 : BUF_X1 port map( A => n2674, Z => n2971);
   U2241 : BUF_X1 port map( A => n2672, Z => n2984);
   U2242 : BUF_X1 port map( A => n2674, Z => n2972);
   U2243 : BUF_X1 port map( A => n2676, Z => n2959);
   U2244 : BUF_X1 port map( A => n2676, Z => n2960);
   U2245 : BUF_X1 port map( A => n2675, Z => n2965);
   U2246 : BUF_X1 port map( A => n2675, Z => n2966);
   U2247 : BUF_X1 port map( A => n2672, Z => n2980);
   U2248 : BUF_X1 port map( A => n2674, Z => n2968);
   U2249 : BUF_X1 port map( A => n2674, Z => n2969);
   U2250 : BUF_X1 port map( A => n2676, Z => n2956);
   U2251 : BUF_X1 port map( A => n2672, Z => n2981);
   U2252 : BUF_X1 port map( A => n2676, Z => n2957);
   U2253 : BUF_X1 port map( A => n2672, Z => n2982);
   U2254 : BUF_X1 port map( A => n2674, Z => n2970);
   U2255 : BUF_X1 port map( A => n2676, Z => n2958);
   U2256 : BUF_X1 port map( A => n2673, Z => n2974);
   U2257 : BUF_X1 port map( A => n2677, Z => n2950);
   U2258 : BUF_X1 port map( A => n2673, Z => n2975);
   U2259 : BUF_X1 port map( A => n2677, Z => n2951);
   U2260 : BUF_X1 port map( A => n2673, Z => n2976);
   U2261 : BUF_X1 port map( A => n2677, Z => n2952);
   U2262 : BUF_X1 port map( A => n2673, Z => n2977);
   U2263 : BUF_X1 port map( A => n2677, Z => n2953);
   U2264 : BUF_X1 port map( A => n2673, Z => n2978);
   U2265 : BUF_X1 port map( A => n2677, Z => n2954);
   U2266 : BUF_X1 port map( A => n2679, Z => n2938);
   U2267 : BUF_X1 port map( A => n2679, Z => n2939);
   U2268 : BUF_X1 port map( A => n2679, Z => n2940);
   U2269 : BUF_X1 port map( A => n2679, Z => n2941);
   U2270 : BUF_X1 port map( A => n2679, Z => n2942);
   U2271 : BUF_X1 port map( A => n2675, Z => n2962);
   U2272 : BUF_X1 port map( A => n2675, Z => n2963);
   U2273 : BUF_X1 port map( A => n2675, Z => n2964);
   U2274 : INV_X1 port map( A => n2933, ZN => n2935);
   U2275 : NOR2_X1 port map( A1 => n2130, A2 => n2133, ZN => enable_io_2_port);
   U2276 : NAND2_X1 port map( A1 => n2131, A2 => n2112, ZN => n2108);
   U2277 : NAND2_X1 port map( A1 => n2133, A2 => n2137, ZN => n2134);
   U2278 : INV_X1 port map( A => n2132, ZN => enable_io_3_port);
   U2279 : AOI21_X1 port map( B1 => n2103, B2 => enable_io_2_port, A => 
                           enable_loc_3_port, ZN => n2132);
   U2280 : OAI21_X1 port map( B1 => n2130, B2 => n2134, A => n2135, ZN => 
                           enable_io_1_port);
   U2281 : INV_X1 port map( A => enable_loc_1_port, ZN => n2135);
   U2282 : AOI21_X1 port map( B1 => n2128, B2 => n2129, A => n3072, ZN => n2145
                           );
   U2283 : NOR2_X1 port map( A1 => n2661, A2 => n2137, ZN => n2143);
   U2284 : NOR2_X1 port map( A1 => n2661, A2 => n2112, ZN => n2147);
   U2285 : NOR2_X1 port map( A1 => n2137, A2 => n2667, ZN => n2159);
   U2286 : NOR2_X1 port map( A1 => n2137, A2 => n2118, ZN => n2160);
   U2287 : NOR2_X1 port map( A1 => n2112, A2 => n2118, ZN => n2153);
   U2288 : NOR2_X1 port map( A1 => n2131, A2 => n2118, ZN => n2156);
   U2289 : NOR2_X1 port map( A1 => n2136, A2 => n2118, ZN => n2158);
   U2290 : NOR2_X1 port map( A1 => n2661, A2 => n2131, ZN => n2144);
   U2291 : BUF_X1 port map( A => n2155, Z => n3016);
   U2292 : BUF_X1 port map( A => n2155, Z => n3017);
   U2293 : BUF_X1 port map( A => n2155, Z => n3018);
   U2294 : BUF_X1 port map( A => n2155, Z => n3019);
   U2295 : BUF_X1 port map( A => n2155, Z => n3020);
   U2296 : NOR2_X1 port map( A1 => n2118, A2 => n2119, ZN => loc_read1_3_port);
   U2297 : NOR2_X1 port map( A1 => n2116, A2 => n2117, ZN => loc_read2_3_port);
   U2298 : NOR2_X1 port map( A1 => n2130, A2 => n2137, ZN => enable_loc_3_port)
                           ;
   U2299 : INV_X1 port map( A => n2113, ZN => n2136);
   U2300 : NOR2_X1 port map( A1 => n2112, A2 => n2130, ZN => enable_loc_1_port)
                           ;
   U2301 : INV_X1 port map( A => n2126, ZN => n2667);
   U2302 : BUF_X1 port map( A => N1235, Z => n3074);
   U2303 : AND2_X1 port map( A1 => n2118, A2 => n2667, ZN => n2154);
   U2304 : BUF_X1 port map( A => N1235, Z => n3075);
   U2305 : NOR2_X1 port map( A1 => n2136, A2 => n2130, ZN => enable_loc_0_port)
                           ;
   U2306 : NOR3_X1 port map( A1 => n2128, A2 => n2129, A3 => n2119, ZN => 
                           global_read1);
   U2307 : NOR2_X1 port map( A1 => n2130, A2 => n2131, ZN => enable_loc_2_port)
                           ;
   U2308 : OR2_X1 port map( A1 => enable_loc_3_port, A2 => enable_loc_0_port, 
                           ZN => enable_io_0_port);
   U2309 : OAI22_X1 port map( A1 => n2137, A2 => n2933, B1 => n2932, B2 => 
                           n2136, ZN => n2677);
   U2310 : OAI22_X1 port map( A1 => n2932, A2 => n2112, B1 => n2134, B2 => 
                           n2933, ZN => n2673);
   U2311 : OAI21_X1 port map( B1 => n2932, B2 => n2137, A => n2934, ZN => n2679
                           );
   U2312 : NOR2_X1 port map( A1 => n2137, A2 => n2116, ZN => n2675);
   U2313 : NOR2_X1 port map( A1 => n2112, A2 => n2116, ZN => n2674);
   U2314 : NOR2_X1 port map( A1 => n2131, A2 => n2116, ZN => n2672);
   U2315 : NOR2_X1 port map( A1 => n2136, A2 => n2116, ZN => n2676);
   U2316 : BUF_X1 port map( A => n2678, Z => n2944);
   U2317 : BUF_X1 port map( A => n2678, Z => n2945);
   U2318 : BUF_X1 port map( A => n2678, Z => n2946);
   U2319 : BUF_X1 port map( A => n2678, Z => n2947);
   U2320 : BUF_X1 port map( A => n2678, Z => n2948);
   U2321 : INV_X1 port map( A => n2124, ZN => n2932);
   U2322 : NAND2_X1 port map( A1 => n2932, A2 => n2116, ZN => n2933);
   U2323 : BUF_X1 port map( A => N1235, Z => n3079);
   U2324 : BUF_X1 port map( A => N1235, Z => n3078);
   U2325 : BUF_X1 port map( A => N1235, Z => n3076);
   U2326 : BUF_X1 port map( A => N1235, Z => n3077);
   U2327 : BUF_X1 port map( A => N1235, Z => n3080);
   U2328 : NAND2_X1 port map( A1 => n1038, A2 => n2109, ZN => n2112);
   U2329 : NAND2_X1 port map( A1 => n2937, A2 => n2103, ZN => n2131);
   U2330 : AOI222_X1 port map( A1 => io_out1_2_4_port, A2 => n3037, B1 => 
                           loc_out1_1_4_port, B2 => n3031, C1 => 
                           global_out1_4_port, C2 => n3025, ZN => n2312);
   U2331 : AOI222_X1 port map( A1 => io_out1_2_5_port, A2 => n3038, B1 => 
                           loc_out1_1_5_port, B2 => n3032, C1 => 
                           global_out1_5_port, C2 => n3026, ZN => n2224);
   U2332 : AOI222_X1 port map( A1 => io_out1_2_6_port, A2 => n3039, B1 => 
                           loc_out1_1_6_port, B2 => n3033, C1 => 
                           global_out1_6_port, C2 => n3027, ZN => n2184);
   U2333 : AOI222_X1 port map( A1 => io_out1_2_7_port, A2 => n3039, B1 => 
                           loc_out1_1_7_port, B2 => n3033, C1 => 
                           global_out1_7_port, C2 => n3027, ZN => n2176);
   U2334 : AOI222_X1 port map( A1 => io_out1_2_8_port, A2 => n3039, B1 => 
                           loc_out1_1_8_port, B2 => n3033, C1 => 
                           global_out1_8_port, C2 => n3027, ZN => n2168);
   U2335 : AOI222_X1 port map( A1 => io_out1_2_9_port, A2 => n3039, B1 => 
                           loc_out1_1_9_port, B2 => n3033, C1 => 
                           global_out1_9_port, C2 => n3027, ZN => n2151);
   U2336 : AOI222_X1 port map( A1 => io_out1_2_42_port, A2 => n3037, B1 => 
                           loc_out1_1_42_port, B2 => n3031, C1 => 
                           global_out1_42_port, C2 => n3025, ZN => n2376);
   U2337 : AOI222_X1 port map( A1 => io_out1_2_43_port, A2 => n3037, B1 => 
                           loc_out1_1_43_port, B2 => n3031, C1 => 
                           global_out1_43_port, C2 => n3025, ZN => n2368);
   U2338 : AOI222_X1 port map( A1 => io_out1_2_44_port, A2 => n3037, B1 => 
                           loc_out1_1_44_port, B2 => n3031, C1 => 
                           global_out1_44_port, C2 => n3025, ZN => n2360);
   U2339 : AOI222_X1 port map( A1 => io_out1_2_45_port, A2 => n3037, B1 => 
                           loc_out1_1_45_port, B2 => n3031, C1 => 
                           global_out1_45_port, C2 => n3025, ZN => n2352);
   U2340 : AOI222_X1 port map( A1 => io_out1_2_46_port, A2 => n3037, B1 => 
                           loc_out1_1_46_port, B2 => n3031, C1 => 
                           global_out1_46_port, C2 => n3025, ZN => n2344);
   U2341 : AOI222_X1 port map( A1 => io_out1_2_47_port, A2 => n3037, B1 => 
                           loc_out1_1_47_port, B2 => n3031, C1 => 
                           global_out1_47_port, C2 => n3025, ZN => n2336);
   U2342 : AOI222_X1 port map( A1 => io_out1_2_48_port, A2 => n3037, B1 => 
                           loc_out1_1_48_port, B2 => n3031, C1 => 
                           global_out1_48_port, C2 => n3025, ZN => n2328);
   U2343 : AOI222_X1 port map( A1 => io_out1_2_49_port, A2 => n3037, B1 => 
                           loc_out1_1_49_port, B2 => n3031, C1 => 
                           global_out1_49_port, C2 => n3025, ZN => n2320);
   U2344 : AOI222_X1 port map( A1 => io_out1_2_50_port, A2 => n3037, B1 => 
                           loc_out1_1_50_port, B2 => n3031, C1 => 
                           global_out1_50_port, C2 => n3025, ZN => n2304);
   U2345 : AOI222_X1 port map( A1 => io_out1_2_51_port, A2 => n3037, B1 => 
                           loc_out1_1_51_port, B2 => n3031, C1 => 
                           global_out1_51_port, C2 => n3025, ZN => n2296);
   U2346 : AOI222_X1 port map( A1 => io_out1_2_52_port, A2 => n3037, B1 => 
                           loc_out1_1_52_port, B2 => n3031, C1 => 
                           global_out1_52_port, C2 => n3025, ZN => n2288);
   U2347 : AOI222_X1 port map( A1 => io_out1_2_53_port, A2 => n3038, B1 => 
                           loc_out1_1_53_port, B2 => n3032, C1 => 
                           global_out1_53_port, C2 => n3026, ZN => n2280);
   U2348 : AOI222_X1 port map( A1 => io_out1_2_54_port, A2 => n3038, B1 => 
                           loc_out1_1_54_port, B2 => n3032, C1 => 
                           global_out1_54_port, C2 => n3026, ZN => n2272);
   U2349 : AOI222_X1 port map( A1 => io_out1_2_55_port, A2 => n3038, B1 => 
                           loc_out1_1_55_port, B2 => n3032, C1 => 
                           global_out1_55_port, C2 => n3026, ZN => n2264);
   U2350 : AOI222_X1 port map( A1 => io_out1_2_56_port, A2 => n3038, B1 => 
                           loc_out1_1_56_port, B2 => n3032, C1 => 
                           global_out1_56_port, C2 => n3026, ZN => n2256);
   U2351 : AOI222_X1 port map( A1 => io_out1_2_57_port, A2 => n3038, B1 => 
                           loc_out1_1_57_port, B2 => n3032, C1 => 
                           global_out1_57_port, C2 => n3026, ZN => n2248);
   U2352 : AOI222_X1 port map( A1 => io_out1_2_58_port, A2 => n3038, B1 => 
                           loc_out1_1_58_port, B2 => n3032, C1 => 
                           global_out1_58_port, C2 => n3026, ZN => n2240);
   U2353 : AOI222_X1 port map( A1 => io_out1_2_59_port, A2 => n3038, B1 => 
                           loc_out1_1_59_port, B2 => n3032, C1 => 
                           global_out1_59_port, C2 => n3026, ZN => n2232);
   U2354 : AOI222_X1 port map( A1 => io_out1_2_60_port, A2 => n3038, B1 => 
                           loc_out1_1_60_port, B2 => n3032, C1 => 
                           global_out1_60_port, C2 => n3026, ZN => n2216);
   U2355 : AOI222_X1 port map( A1 => io_out1_2_61_port, A2 => n3038, B1 => 
                           loc_out1_1_61_port, B2 => n3032, C1 => 
                           global_out1_61_port, C2 => n3026, ZN => n2208);
   U2356 : AOI222_X1 port map( A1 => io_out1_2_62_port, A2 => n3038, B1 => 
                           loc_out1_1_62_port, B2 => n3032, C1 => 
                           global_out1_62_port, C2 => n3026, ZN => n2200);
   U2357 : AOI222_X1 port map( A1 => io_out1_2_63_port, A2 => n3038, B1 => 
                           loc_out1_1_63_port, B2 => n3032, C1 => 
                           global_out1_63_port, C2 => n3026, ZN => n2192);
   U2358 : AOI222_X1 port map( A1 => io_out1_2_2_port, A2 => n3035, B1 => 
                           loc_out1_1_2_port, B2 => n3029, C1 => 
                           global_out1_2_port, C2 => n3023, ZN => n2488);
   U2359 : AOI222_X1 port map( A1 => io_out1_2_3_port, A2 => n3036, B1 => 
                           loc_out1_1_3_port, B2 => n3030, C1 => 
                           global_out1_3_port, C2 => n3024, ZN => n2400);
   U2360 : AOI222_X1 port map( A1 => io_out1_2_20_port, A2 => n3035, B1 => 
                           loc_out1_1_20_port, B2 => n3029, C1 => 
                           global_out1_20_port, C2 => n3023, ZN => n2568);
   U2361 : AOI222_X1 port map( A1 => io_out1_2_21_port, A2 => n3035, B1 => 
                           loc_out1_1_21_port, B2 => n3029, C1 => 
                           global_out1_21_port, C2 => n3023, ZN => n2560);
   U2362 : AOI222_X1 port map( A1 => io_out1_2_22_port, A2 => n3035, B1 => 
                           loc_out1_1_22_port, B2 => n3029, C1 => 
                           global_out1_22_port, C2 => n3023, ZN => n2552);
   U2363 : AOI222_X1 port map( A1 => io_out1_2_23_port, A2 => n3035, B1 => 
                           loc_out1_1_23_port, B2 => n3029, C1 => 
                           global_out1_23_port, C2 => n3023, ZN => n2544);
   U2364 : AOI222_X1 port map( A1 => io_out1_2_24_port, A2 => n3035, B1 => 
                           loc_out1_1_24_port, B2 => n3029, C1 => 
                           global_out1_24_port, C2 => n3023, ZN => n2536);
   U2365 : AOI222_X1 port map( A1 => io_out1_2_25_port, A2 => n3035, B1 => 
                           loc_out1_1_25_port, B2 => n3029, C1 => 
                           global_out1_25_port, C2 => n3023, ZN => n2528);
   U2366 : AOI222_X1 port map( A1 => io_out1_2_26_port, A2 => n3035, B1 => 
                           loc_out1_1_26_port, B2 => n3029, C1 => 
                           global_out1_26_port, C2 => n3023, ZN => n2520);
   U2367 : AOI222_X1 port map( A1 => io_out1_2_27_port, A2 => n3035, B1 => 
                           loc_out1_1_27_port, B2 => n3029, C1 => 
                           global_out1_27_port, C2 => n3023, ZN => n2512);
   U2368 : AOI222_X1 port map( A1 => io_out1_2_28_port, A2 => n3035, B1 => 
                           loc_out1_1_28_port, B2 => n3029, C1 => 
                           global_out1_28_port, C2 => n3023, ZN => n2504);
   U2369 : AOI222_X1 port map( A1 => io_out1_2_29_port, A2 => n3035, B1 => 
                           loc_out1_1_29_port, B2 => n3029, C1 => 
                           global_out1_29_port, C2 => n3023, ZN => n2496);
   U2370 : AOI222_X1 port map( A1 => io_out1_2_30_port, A2 => n3035, B1 => 
                           loc_out1_1_30_port, B2 => n3029, C1 => 
                           global_out1_30_port, C2 => n3023, ZN => n2480);
   U2371 : AOI222_X1 port map( A1 => io_out1_2_31_port, A2 => n3036, B1 => 
                           loc_out1_1_31_port, B2 => n3030, C1 => 
                           global_out1_31_port, C2 => n3024, ZN => n2472);
   U2372 : AOI222_X1 port map( A1 => io_out1_2_32_port, A2 => n3036, B1 => 
                           loc_out1_1_32_port, B2 => n3030, C1 => 
                           global_out1_32_port, C2 => n3024, ZN => n2464);
   U2373 : AOI222_X1 port map( A1 => io_out1_2_33_port, A2 => n3036, B1 => 
                           loc_out1_1_33_port, B2 => n3030, C1 => 
                           global_out1_33_port, C2 => n3024, ZN => n2456);
   U2374 : AOI222_X1 port map( A1 => io_out1_2_34_port, A2 => n3036, B1 => 
                           loc_out1_1_34_port, B2 => n3030, C1 => 
                           global_out1_34_port, C2 => n3024, ZN => n2448);
   U2375 : AOI222_X1 port map( A1 => io_out1_2_35_port, A2 => n3036, B1 => 
                           loc_out1_1_35_port, B2 => n3030, C1 => 
                           global_out1_35_port, C2 => n3024, ZN => n2440);
   U2376 : AOI222_X1 port map( A1 => io_out1_2_36_port, A2 => n3036, B1 => 
                           loc_out1_1_36_port, B2 => n3030, C1 => 
                           global_out1_36_port, C2 => n3024, ZN => n2432);
   U2377 : AOI222_X1 port map( A1 => io_out1_2_37_port, A2 => n3036, B1 => 
                           loc_out1_1_37_port, B2 => n3030, C1 => 
                           global_out1_37_port, C2 => n3024, ZN => n2424);
   U2378 : AOI222_X1 port map( A1 => io_out1_2_38_port, A2 => n3036, B1 => 
                           loc_out1_1_38_port, B2 => n3030, C1 => 
                           global_out1_38_port, C2 => n3024, ZN => n2416);
   U2379 : AOI222_X1 port map( A1 => io_out1_2_39_port, A2 => n3036, B1 => 
                           loc_out1_1_39_port, B2 => n3030, C1 => 
                           global_out1_39_port, C2 => n3024, ZN => n2408);
   U2380 : AOI222_X1 port map( A1 => io_out1_2_40_port, A2 => n3036, B1 => 
                           loc_out1_1_40_port, B2 => n3030, C1 => 
                           global_out1_40_port, C2 => n3024, ZN => n2392);
   U2381 : AOI222_X1 port map( A1 => io_out1_2_41_port, A2 => n3036, B1 => 
                           loc_out1_1_41_port, B2 => n3030, C1 => 
                           global_out1_41_port, C2 => n3024, ZN => n2384);
   U2382 : AOI222_X1 port map( A1 => io_out1_2_0_port, A2 => n3034, B1 => 
                           loc_out1_1_0_port, B2 => n3028, C1 => 
                           global_out1_0_port, C2 => n3022, ZN => n2666);
   U2383 : AOI222_X1 port map( A1 => io_out1_2_1_port, A2 => n3034, B1 => 
                           loc_out1_1_1_port, B2 => n3028, C1 => 
                           global_out1_1_port, C2 => n3022, ZN => n2576);
   U2384 : AOI222_X1 port map( A1 => io_out1_2_10_port, A2 => n3034, B1 => 
                           loc_out1_1_10_port, B2 => n3028, C1 => 
                           global_out1_10_port, C2 => n3022, ZN => n2656);
   U2385 : AOI222_X1 port map( A1 => io_out1_2_11_port, A2 => n3034, B1 => 
                           loc_out1_1_11_port, B2 => n3028, C1 => 
                           global_out1_11_port, C2 => n3022, ZN => n2648);
   U2386 : AOI222_X1 port map( A1 => io_out1_2_12_port, A2 => n3034, B1 => 
                           loc_out1_1_12_port, B2 => n3028, C1 => 
                           global_out1_12_port, C2 => n3022, ZN => n2640);
   U2387 : AOI222_X1 port map( A1 => io_out1_2_13_port, A2 => n3034, B1 => 
                           loc_out1_1_13_port, B2 => n3028, C1 => 
                           global_out1_13_port, C2 => n3022, ZN => n2632);
   U2388 : AOI222_X1 port map( A1 => io_out1_2_14_port, A2 => n3034, B1 => 
                           loc_out1_1_14_port, B2 => n3028, C1 => 
                           global_out1_14_port, C2 => n3022, ZN => n2624);
   U2389 : AOI222_X1 port map( A1 => io_out1_2_15_port, A2 => n3034, B1 => 
                           loc_out1_1_15_port, B2 => n3028, C1 => 
                           global_out1_15_port, C2 => n3022, ZN => n2616);
   U2390 : AOI222_X1 port map( A1 => io_out1_2_16_port, A2 => n3034, B1 => 
                           loc_out1_1_16_port, B2 => n3028, C1 => 
                           global_out1_16_port, C2 => n3022, ZN => n2608);
   U2391 : AOI222_X1 port map( A1 => io_out1_2_17_port, A2 => n3034, B1 => 
                           loc_out1_1_17_port, B2 => n3028, C1 => 
                           global_out1_17_port, C2 => n3022, ZN => n2600);
   U2392 : AOI222_X1 port map( A1 => io_out1_2_18_port, A2 => n3034, B1 => 
                           loc_out1_1_18_port, B2 => n3028, C1 => 
                           global_out1_18_port, C2 => n3022, ZN => n2592);
   U2393 : AOI222_X1 port map( A1 => io_out1_2_19_port, A2 => n3034, B1 => 
                           loc_out1_1_19_port, B2 => n3028, C1 => 
                           global_out1_19_port, C2 => n3022, ZN => n2584);
   U2394 : OAI211_X1 port map( C1 => n3069, C2 => n2465, A => n2466, B => n2467
                           , ZN => OUT1(31));
   U2395 : INV_X1 port map( A => io_out1_0_31_port, ZN => n2465);
   U2396 : AOI22_X1 port map( A1 => n3048, A2 => n2468, B1 => io_out1_1_31_port
                           , B2 => n3043, ZN => n2466);
   U2397 : AOI222_X1 port map( A1 => global_out1_31_port, A2 => n3073, B1 => 
                           io_out1_3_31_port, B2 => n3061, C1 => 
                           io_out1_2_31_port, C2 => n3054, ZN => n2467);
   U2398 : OAI211_X1 port map( C1 => n3068, C2 => n2457, A => n2458, B => n2459
                           , ZN => OUT1(32));
   U2399 : INV_X1 port map( A => io_out1_0_32_port, ZN => n2457);
   U2400 : AOI22_X1 port map( A1 => n3048, A2 => n2460, B1 => io_out1_1_32_port
                           , B2 => n3043, ZN => n2458);
   U2401 : AOI222_X1 port map( A1 => global_out1_32_port, A2 => n3073, B1 => 
                           io_out1_3_32_port, B2 => n3061, C1 => 
                           io_out1_2_32_port, C2 => n3054, ZN => n2459);
   U2402 : OAI211_X1 port map( C1 => n3068, C2 => n2449, A => n2450, B => n2451
                           , ZN => OUT1(33));
   U2403 : INV_X1 port map( A => io_out1_0_33_port, ZN => n2449);
   U2404 : AOI22_X1 port map( A1 => n3048, A2 => n2452, B1 => io_out1_1_33_port
                           , B2 => n3043, ZN => n2450);
   U2405 : AOI222_X1 port map( A1 => global_out1_33_port, A2 => n3073, B1 => 
                           io_out1_3_33_port, B2 => n3061, C1 => 
                           io_out1_2_33_port, C2 => n3054, ZN => n2451);
   U2406 : OAI211_X1 port map( C1 => n3070, C2 => n2649, A => n2650, B => n2651
                           , ZN => OUT1(10));
   U2407 : INV_X1 port map( A => io_out1_0_10_port, ZN => n2649);
   U2408 : AOI22_X1 port map( A1 => n3046, A2 => n2652, B1 => io_out1_1_10_port
                           , B2 => n3045, ZN => n2650);
   U2409 : AOI222_X1 port map( A1 => global_out1_10_port, A2 => n3073, B1 => 
                           io_out1_3_10_port, B2 => n3063, C1 => 
                           io_out1_2_10_port, C2 => n3052, ZN => n2651);
   U2410 : OAI211_X1 port map( C1 => n3070, C2 => n2633, A => n2634, B => n2635
                           , ZN => OUT1(12));
   U2411 : INV_X1 port map( A => io_out1_0_12_port, ZN => n2633);
   U2412 : AOI22_X1 port map( A1 => n3046, A2 => n2636, B1 => io_out1_1_12_port
                           , B2 => n3045, ZN => n2634);
   U2413 : AOI222_X1 port map( A1 => global_out1_12_port, A2 => n3071, B1 => 
                           io_out1_3_12_port, B2 => n3063, C1 => 
                           io_out1_2_12_port, C2 => n3052, ZN => n2635);
   U2414 : NOR3_X1 port map( A1 => n2114, A2 => ADD_WR(2), A3 => n2115, ZN => 
                           loc_write_3_port);
   U2415 : INV_X1 port map( A => ADD_WR(3), ZN => n2115);
   U2416 : NOR3_X1 port map( A1 => n2120, A2 => ADD_WR(3), A3 => n2114, ZN => 
                           io_write_3_port);
   U2417 : XNOR2_X1 port map( A => n2103, B => ADD_WR(2), ZN => n2120);
   U2418 : NAND2_X1 port map( A1 => n2937, A2 => n1038, ZN => n2137);
   U2419 : OR2_X1 port map( A1 => n2123, A2 => ADD_RD2(2), ZN => n2116);
   U2420 : AOI21_X1 port map( B1 => n2121, B2 => n2122, A => n2117, ZN => 
                           io_read2_3_port);
   U2421 : NAND2_X1 port map( A1 => n2124, A2 => n2103, ZN => n2121);
   U2422 : NAND2_X1 port map( A1 => ADD_RD1(3), A2 => n2128, ZN => n2118);
   U2423 : INV_X1 port map( A => ENABLE, ZN => n2130);
   U2424 : NOR2_X1 port map( A1 => n2125, A2 => n2119, ZN => io_read1_3_port);
   U2425 : AOI21_X1 port map( B1 => n2126, B2 => n1038, A => n2127, ZN => n2125
                           );
   U2426 : NOR3_X1 port map( A1 => ADD_RD1(2), A2 => n1038, A3 => ADD_RD1(3), 
                           ZN => n2127);
   U2427 : NOR2_X1 port map( A1 => n2937, A2 => n1038, ZN => n2113);
   U2428 : NOR2_X1 port map( A1 => n2128, A2 => ADD_RD1(3), ZN => n2126);
   U2429 : NOR2_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(2), ZN => n2124);
   U2430 : AOI21_X1 port map( B1 => n1038, B2 => n2112, A => n2113, ZN => n2110
                           );
   U2431 : INV_X1 port map( A => ADD_RD1(2), ZN => n2128);
   U2432 : NAND2_X1 port map( A1 => ADD_RD2(3), A2 => n2116, ZN => N1235);
   U2433 : NAND4_X1 port map( A1 => n2309, A2 => n2310, A3 => n2311, A4 => 
                           n2312, ZN => n2308);
   U2434 : AOI22_X1 port map( A1 => io_out1_0_4_port, A2 => n2995, B1 => 
                           loc_out1_3_4_port, B2 => n2989, ZN => n2309);
   U2435 : AOI22_X1 port map( A1 => io_out1_1_4_port, A2 => n3007, B1 => 
                           loc_out1_0_4_port, B2 => n3001, ZN => n2310);
   U2436 : AOI22_X1 port map( A1 => io_out1_3_4_port, A2 => n3019, B1 => 
                           loc_out1_2_4_port, B2 => n3013, ZN => n2311);
   U2437 : NAND4_X1 port map( A1 => n2221, A2 => n2222, A3 => n2223, A4 => 
                           n2224, ZN => n2220);
   U2438 : AOI22_X1 port map( A1 => io_out1_0_5_port, A2 => n2996, B1 => 
                           loc_out1_3_5_port, B2 => n2990, ZN => n2221);
   U2439 : AOI22_X1 port map( A1 => io_out1_1_5_port, A2 => n3008, B1 => 
                           loc_out1_0_5_port, B2 => n3002, ZN => n2222);
   U2440 : AOI22_X1 port map( A1 => io_out1_3_5_port, A2 => n3020, B1 => 
                           loc_out1_2_5_port, B2 => n3014, ZN => n2223);
   U2441 : NAND4_X1 port map( A1 => n2181, A2 => n2182, A3 => n2183, A4 => 
                           n2184, ZN => n2180);
   U2442 : AOI22_X1 port map( A1 => io_out1_0_6_port, A2 => n2997, B1 => 
                           loc_out1_3_6_port, B2 => n2991, ZN => n2181);
   U2443 : AOI22_X1 port map( A1 => io_out1_1_6_port, A2 => n3009, B1 => 
                           loc_out1_0_6_port, B2 => n3003, ZN => n2182);
   U2444 : AOI22_X1 port map( A1 => io_out1_3_6_port, A2 => n3021, B1 => 
                           loc_out1_2_6_port, B2 => n3015, ZN => n2183);
   U2445 : NAND4_X1 port map( A1 => n2173, A2 => n2174, A3 => n2175, A4 => 
                           n2176, ZN => n2172);
   U2446 : AOI22_X1 port map( A1 => io_out1_0_7_port, A2 => n2997, B1 => 
                           loc_out1_3_7_port, B2 => n2991, ZN => n2173);
   U2447 : AOI22_X1 port map( A1 => io_out1_1_7_port, A2 => n3009, B1 => 
                           loc_out1_0_7_port, B2 => n3003, ZN => n2174);
   U2448 : AOI22_X1 port map( A1 => io_out1_3_7_port, A2 => n3021, B1 => 
                           loc_out1_2_7_port, B2 => n3015, ZN => n2175);
   U2449 : NAND4_X1 port map( A1 => n2165, A2 => n2166, A3 => n2167, A4 => 
                           n2168, ZN => n2164);
   U2450 : AOI22_X1 port map( A1 => io_out1_0_8_port, A2 => n2997, B1 => 
                           loc_out1_3_8_port, B2 => n2991, ZN => n2165);
   U2451 : AOI22_X1 port map( A1 => io_out1_1_8_port, A2 => n3009, B1 => 
                           loc_out1_0_8_port, B2 => n3003, ZN => n2166);
   U2452 : AOI22_X1 port map( A1 => io_out1_3_8_port, A2 => n3021, B1 => 
                           loc_out1_2_8_port, B2 => n3015, ZN => n2167);
   U2453 : NAND4_X1 port map( A1 => n2148, A2 => n2149, A3 => n2150, A4 => 
                           n2151, ZN => n2146);
   U2454 : AOI22_X1 port map( A1 => io_out1_0_9_port, A2 => n2997, B1 => 
                           loc_out1_3_9_port, B2 => n2991, ZN => n2148);
   U2455 : AOI22_X1 port map( A1 => io_out1_1_9_port, A2 => n3009, B1 => 
                           loc_out1_0_9_port, B2 => n3003, ZN => n2149);
   U2456 : AOI22_X1 port map( A1 => io_out1_3_9_port, A2 => n3021, B1 => 
                           loc_out1_2_9_port, B2 => n3015, ZN => n2150);
   U2457 : NAND4_X1 port map( A1 => n2373, A2 => n2374, A3 => n2375, A4 => 
                           n2376, ZN => n2372);
   U2458 : AOI22_X1 port map( A1 => io_out1_0_42_port, A2 => n2995, B1 => 
                           loc_out1_3_42_port, B2 => n2989, ZN => n2373);
   U2459 : AOI22_X1 port map( A1 => io_out1_1_42_port, A2 => n3007, B1 => 
                           loc_out1_0_42_port, B2 => n3001, ZN => n2374);
   U2460 : AOI22_X1 port map( A1 => io_out1_3_42_port, A2 => n3019, B1 => 
                           loc_out1_2_42_port, B2 => n3013, ZN => n2375);
   U2461 : NAND4_X1 port map( A1 => n2365, A2 => n2366, A3 => n2367, A4 => 
                           n2368, ZN => n2364);
   U2462 : AOI22_X1 port map( A1 => io_out1_0_43_port, A2 => n2995, B1 => 
                           loc_out1_3_43_port, B2 => n2989, ZN => n2365);
   U2463 : AOI22_X1 port map( A1 => io_out1_1_43_port, A2 => n3007, B1 => 
                           loc_out1_0_43_port, B2 => n3001, ZN => n2366);
   U2464 : AOI22_X1 port map( A1 => io_out1_3_43_port, A2 => n3019, B1 => 
                           loc_out1_2_43_port, B2 => n3013, ZN => n2367);
   U2465 : NAND4_X1 port map( A1 => n2357, A2 => n2358, A3 => n2359, A4 => 
                           n2360, ZN => n2356);
   U2466 : AOI22_X1 port map( A1 => io_out1_0_44_port, A2 => n2995, B1 => 
                           loc_out1_3_44_port, B2 => n2989, ZN => n2357);
   U2467 : AOI22_X1 port map( A1 => io_out1_1_44_port, A2 => n3007, B1 => 
                           loc_out1_0_44_port, B2 => n3001, ZN => n2358);
   U2468 : AOI22_X1 port map( A1 => io_out1_3_44_port, A2 => n3019, B1 => 
                           loc_out1_2_44_port, B2 => n3013, ZN => n2359);
   U2469 : NAND4_X1 port map( A1 => n2349, A2 => n2350, A3 => n2351, A4 => 
                           n2352, ZN => n2348);
   U2470 : AOI22_X1 port map( A1 => io_out1_0_45_port, A2 => n2995, B1 => 
                           loc_out1_3_45_port, B2 => n2989, ZN => n2349);
   U2471 : AOI22_X1 port map( A1 => io_out1_1_45_port, A2 => n3007, B1 => 
                           loc_out1_0_45_port, B2 => n3001, ZN => n2350);
   U2472 : AOI22_X1 port map( A1 => io_out1_3_45_port, A2 => n3019, B1 => 
                           loc_out1_2_45_port, B2 => n3013, ZN => n2351);
   U2473 : NAND4_X1 port map( A1 => n2341, A2 => n2342, A3 => n2343, A4 => 
                           n2344, ZN => n2340);
   U2474 : AOI22_X1 port map( A1 => io_out1_0_46_port, A2 => n2995, B1 => 
                           loc_out1_3_46_port, B2 => n2989, ZN => n2341);
   U2475 : AOI22_X1 port map( A1 => io_out1_1_46_port, A2 => n3007, B1 => 
                           loc_out1_0_46_port, B2 => n3001, ZN => n2342);
   U2476 : AOI22_X1 port map( A1 => io_out1_3_46_port, A2 => n3019, B1 => 
                           loc_out1_2_46_port, B2 => n3013, ZN => n2343);
   U2477 : NAND4_X1 port map( A1 => n2333, A2 => n2334, A3 => n2335, A4 => 
                           n2336, ZN => n2332);
   U2478 : AOI22_X1 port map( A1 => io_out1_0_47_port, A2 => n2995, B1 => 
                           loc_out1_3_47_port, B2 => n2989, ZN => n2333);
   U2479 : AOI22_X1 port map( A1 => io_out1_1_47_port, A2 => n3007, B1 => 
                           loc_out1_0_47_port, B2 => n3001, ZN => n2334);
   U2480 : AOI22_X1 port map( A1 => io_out1_3_47_port, A2 => n3019, B1 => 
                           loc_out1_2_47_port, B2 => n3013, ZN => n2335);
   U2481 : NAND4_X1 port map( A1 => n2325, A2 => n2326, A3 => n2327, A4 => 
                           n2328, ZN => n2324);
   U2482 : AOI22_X1 port map( A1 => io_out1_0_48_port, A2 => n2995, B1 => 
                           loc_out1_3_48_port, B2 => n2989, ZN => n2325);
   U2483 : AOI22_X1 port map( A1 => io_out1_1_48_port, A2 => n3007, B1 => 
                           loc_out1_0_48_port, B2 => n3001, ZN => n2326);
   U2484 : AOI22_X1 port map( A1 => io_out1_3_48_port, A2 => n3019, B1 => 
                           loc_out1_2_48_port, B2 => n3013, ZN => n2327);
   U2485 : NAND4_X1 port map( A1 => n2317, A2 => n2318, A3 => n2319, A4 => 
                           n2320, ZN => n2316);
   U2486 : AOI22_X1 port map( A1 => io_out1_0_49_port, A2 => n2995, B1 => 
                           loc_out1_3_49_port, B2 => n2989, ZN => n2317);
   U2487 : AOI22_X1 port map( A1 => io_out1_1_49_port, A2 => n3007, B1 => 
                           loc_out1_0_49_port, B2 => n3001, ZN => n2318);
   U2488 : AOI22_X1 port map( A1 => io_out1_3_49_port, A2 => n3019, B1 => 
                           loc_out1_2_49_port, B2 => n3013, ZN => n2319);
   U2489 : NAND4_X1 port map( A1 => n2301, A2 => n2302, A3 => n2303, A4 => 
                           n2304, ZN => n2300);
   U2490 : AOI22_X1 port map( A1 => io_out1_0_50_port, A2 => n2995, B1 => 
                           loc_out1_3_50_port, B2 => n2989, ZN => n2301);
   U2491 : AOI22_X1 port map( A1 => io_out1_1_50_port, A2 => n3007, B1 => 
                           loc_out1_0_50_port, B2 => n3001, ZN => n2302);
   U2492 : AOI22_X1 port map( A1 => io_out1_3_50_port, A2 => n3019, B1 => 
                           loc_out1_2_50_port, B2 => n3013, ZN => n2303);
   U2493 : NAND4_X1 port map( A1 => n2293, A2 => n2294, A3 => n2295, A4 => 
                           n2296, ZN => n2292);
   U2494 : AOI22_X1 port map( A1 => io_out1_0_51_port, A2 => n2995, B1 => 
                           loc_out1_3_51_port, B2 => n2989, ZN => n2293);
   U2495 : AOI22_X1 port map( A1 => io_out1_1_51_port, A2 => n3007, B1 => 
                           loc_out1_0_51_port, B2 => n3001, ZN => n2294);
   U2496 : AOI22_X1 port map( A1 => io_out1_3_51_port, A2 => n3019, B1 => 
                           loc_out1_2_51_port, B2 => n3013, ZN => n2295);
   U2497 : NAND4_X1 port map( A1 => n2285, A2 => n2286, A3 => n2287, A4 => 
                           n2288, ZN => n2284);
   U2498 : AOI22_X1 port map( A1 => io_out1_0_52_port, A2 => n2995, B1 => 
                           loc_out1_3_52_port, B2 => n2989, ZN => n2285);
   U2499 : AOI22_X1 port map( A1 => io_out1_1_52_port, A2 => n3007, B1 => 
                           loc_out1_0_52_port, B2 => n3001, ZN => n2286);
   U2500 : AOI22_X1 port map( A1 => io_out1_3_52_port, A2 => n3019, B1 => 
                           loc_out1_2_52_port, B2 => n3013, ZN => n2287);
   U2501 : NAND4_X1 port map( A1 => n2277, A2 => n2278, A3 => n2279, A4 => 
                           n2280, ZN => n2276);
   U2502 : AOI22_X1 port map( A1 => io_out1_0_53_port, A2 => n2996, B1 => 
                           loc_out1_3_53_port, B2 => n2990, ZN => n2277);
   U2503 : AOI22_X1 port map( A1 => io_out1_1_53_port, A2 => n3008, B1 => 
                           loc_out1_0_53_port, B2 => n3002, ZN => n2278);
   U2504 : AOI22_X1 port map( A1 => io_out1_3_53_port, A2 => n3020, B1 => 
                           loc_out1_2_53_port, B2 => n3014, ZN => n2279);
   U2505 : NAND4_X1 port map( A1 => n2269, A2 => n2270, A3 => n2271, A4 => 
                           n2272, ZN => n2268);
   U2506 : AOI22_X1 port map( A1 => io_out1_0_54_port, A2 => n2996, B1 => 
                           loc_out1_3_54_port, B2 => n2990, ZN => n2269);
   U2507 : AOI22_X1 port map( A1 => io_out1_1_54_port, A2 => n3008, B1 => 
                           loc_out1_0_54_port, B2 => n3002, ZN => n2270);
   U2508 : AOI22_X1 port map( A1 => io_out1_3_54_port, A2 => n3020, B1 => 
                           loc_out1_2_54_port, B2 => n3014, ZN => n2271);
   U2509 : NAND4_X1 port map( A1 => n2261, A2 => n2262, A3 => n2263, A4 => 
                           n2264, ZN => n2260);
   U2510 : AOI22_X1 port map( A1 => io_out1_0_55_port, A2 => n2996, B1 => 
                           loc_out1_3_55_port, B2 => n2990, ZN => n2261);
   U2511 : AOI22_X1 port map( A1 => io_out1_1_55_port, A2 => n3008, B1 => 
                           loc_out1_0_55_port, B2 => n3002, ZN => n2262);
   U2512 : AOI22_X1 port map( A1 => io_out1_3_55_port, A2 => n3020, B1 => 
                           loc_out1_2_55_port, B2 => n3014, ZN => n2263);
   U2513 : NAND4_X1 port map( A1 => n2253, A2 => n2254, A3 => n2255, A4 => 
                           n2256, ZN => n2252);
   U2514 : AOI22_X1 port map( A1 => io_out1_0_56_port, A2 => n2996, B1 => 
                           loc_out1_3_56_port, B2 => n2990, ZN => n2253);
   U2515 : AOI22_X1 port map( A1 => io_out1_1_56_port, A2 => n3008, B1 => 
                           loc_out1_0_56_port, B2 => n3002, ZN => n2254);
   U2516 : AOI22_X1 port map( A1 => io_out1_3_56_port, A2 => n3020, B1 => 
                           loc_out1_2_56_port, B2 => n3014, ZN => n2255);
   U2517 : NAND4_X1 port map( A1 => n2245, A2 => n2246, A3 => n2247, A4 => 
                           n2248, ZN => n2244);
   U2518 : AOI22_X1 port map( A1 => io_out1_0_57_port, A2 => n2996, B1 => 
                           loc_out1_3_57_port, B2 => n2990, ZN => n2245);
   U2519 : AOI22_X1 port map( A1 => io_out1_1_57_port, A2 => n3008, B1 => 
                           loc_out1_0_57_port, B2 => n3002, ZN => n2246);
   U2520 : AOI22_X1 port map( A1 => io_out1_3_57_port, A2 => n3020, B1 => 
                           loc_out1_2_57_port, B2 => n3014, ZN => n2247);
   U2521 : NAND4_X1 port map( A1 => n2237, A2 => n2238, A3 => n2239, A4 => 
                           n2240, ZN => n2236);
   U2522 : AOI22_X1 port map( A1 => io_out1_0_58_port, A2 => n2996, B1 => 
                           loc_out1_3_58_port, B2 => n2990, ZN => n2237);
   U2523 : AOI22_X1 port map( A1 => io_out1_1_58_port, A2 => n3008, B1 => 
                           loc_out1_0_58_port, B2 => n3002, ZN => n2238);
   U2524 : AOI22_X1 port map( A1 => io_out1_3_58_port, A2 => n3020, B1 => 
                           loc_out1_2_58_port, B2 => n3014, ZN => n2239);
   U2525 : NAND4_X1 port map( A1 => n2229, A2 => n2230, A3 => n2231, A4 => 
                           n2232, ZN => n2228);
   U2526 : AOI22_X1 port map( A1 => io_out1_0_59_port, A2 => n2996, B1 => 
                           loc_out1_3_59_port, B2 => n2990, ZN => n2229);
   U2527 : AOI22_X1 port map( A1 => io_out1_1_59_port, A2 => n3008, B1 => 
                           loc_out1_0_59_port, B2 => n3002, ZN => n2230);
   U2528 : AOI22_X1 port map( A1 => io_out1_3_59_port, A2 => n3020, B1 => 
                           loc_out1_2_59_port, B2 => n3014, ZN => n2231);
   U2529 : NAND4_X1 port map( A1 => n2213, A2 => n2214, A3 => n2215, A4 => 
                           n2216, ZN => n2212);
   U2530 : AOI22_X1 port map( A1 => io_out1_0_60_port, A2 => n2996, B1 => 
                           loc_out1_3_60_port, B2 => n2990, ZN => n2213);
   U2531 : AOI22_X1 port map( A1 => io_out1_1_60_port, A2 => n3008, B1 => 
                           loc_out1_0_60_port, B2 => n3002, ZN => n2214);
   U2532 : AOI22_X1 port map( A1 => io_out1_3_60_port, A2 => n3020, B1 => 
                           loc_out1_2_60_port, B2 => n3014, ZN => n2215);
   U2533 : NAND4_X1 port map( A1 => n2205, A2 => n2206, A3 => n2207, A4 => 
                           n2208, ZN => n2204);
   U2534 : AOI22_X1 port map( A1 => io_out1_0_61_port, A2 => n2996, B1 => 
                           loc_out1_3_61_port, B2 => n2990, ZN => n2205);
   U2535 : AOI22_X1 port map( A1 => io_out1_1_61_port, A2 => n3008, B1 => 
                           loc_out1_0_61_port, B2 => n3002, ZN => n2206);
   U2536 : AOI22_X1 port map( A1 => io_out1_3_61_port, A2 => n3020, B1 => 
                           loc_out1_2_61_port, B2 => n3014, ZN => n2207);
   U2537 : NAND4_X1 port map( A1 => n2197, A2 => n2198, A3 => n2199, A4 => 
                           n2200, ZN => n2196);
   U2538 : AOI22_X1 port map( A1 => io_out1_0_62_port, A2 => n2996, B1 => 
                           loc_out1_3_62_port, B2 => n2990, ZN => n2197);
   U2539 : AOI22_X1 port map( A1 => io_out1_1_62_port, A2 => n3008, B1 => 
                           loc_out1_0_62_port, B2 => n3002, ZN => n2198);
   U2540 : AOI22_X1 port map( A1 => io_out1_3_62_port, A2 => n3020, B1 => 
                           loc_out1_2_62_port, B2 => n3014, ZN => n2199);
   U2541 : NAND4_X1 port map( A1 => n2189, A2 => n2190, A3 => n2191, A4 => 
                           n2192, ZN => n2188);
   U2542 : AOI22_X1 port map( A1 => io_out1_0_63_port, A2 => n2996, B1 => 
                           loc_out1_3_63_port, B2 => n2990, ZN => n2189);
   U2543 : AOI22_X1 port map( A1 => io_out1_1_63_port, A2 => n3008, B1 => 
                           loc_out1_0_63_port, B2 => n3002, ZN => n2190);
   U2544 : AOI22_X1 port map( A1 => io_out1_3_63_port, A2 => n3020, B1 => 
                           loc_out1_2_63_port, B2 => n3014, ZN => n2191);
   U2545 : NAND4_X1 port map( A1 => n2485, A2 => n2486, A3 => n2487, A4 => 
                           n2488, ZN => n2484);
   U2546 : AOI22_X1 port map( A1 => io_out1_0_2_port, A2 => n2993, B1 => 
                           loc_out1_3_2_port, B2 => n2987, ZN => n2485);
   U2547 : AOI22_X1 port map( A1 => io_out1_1_2_port, A2 => n3005, B1 => 
                           loc_out1_0_2_port, B2 => n2999, ZN => n2486);
   U2548 : AOI22_X1 port map( A1 => io_out1_3_2_port, A2 => n3017, B1 => 
                           loc_out1_2_2_port, B2 => n3011, ZN => n2487);
   U2549 : NAND4_X1 port map( A1 => n2397, A2 => n2398, A3 => n2399, A4 => 
                           n2400, ZN => n2396);
   U2550 : AOI22_X1 port map( A1 => io_out1_0_3_port, A2 => n2994, B1 => 
                           loc_out1_3_3_port, B2 => n2988, ZN => n2397);
   U2551 : AOI22_X1 port map( A1 => io_out1_1_3_port, A2 => n3006, B1 => 
                           loc_out1_0_3_port, B2 => n3000, ZN => n2398);
   U2552 : AOI22_X1 port map( A1 => io_out1_3_3_port, A2 => n3018, B1 => 
                           loc_out1_2_3_port, B2 => n3012, ZN => n2399);
   U2553 : NAND4_X1 port map( A1 => n2565, A2 => n2566, A3 => n2567, A4 => 
                           n2568, ZN => n2564);
   U2554 : AOI22_X1 port map( A1 => io_out1_0_20_port, A2 => n2993, B1 => 
                           loc_out1_3_20_port, B2 => n2987, ZN => n2565);
   U2555 : AOI22_X1 port map( A1 => io_out1_1_20_port, A2 => n3005, B1 => 
                           loc_out1_0_20_port, B2 => n2999, ZN => n2566);
   U2556 : AOI22_X1 port map( A1 => io_out1_3_20_port, A2 => n3017, B1 => 
                           loc_out1_2_20_port, B2 => n3011, ZN => n2567);
   U2557 : NAND4_X1 port map( A1 => n2557, A2 => n2558, A3 => n2559, A4 => 
                           n2560, ZN => n2556);
   U2558 : AOI22_X1 port map( A1 => io_out1_0_21_port, A2 => n2993, B1 => 
                           loc_out1_3_21_port, B2 => n2987, ZN => n2557);
   U2559 : AOI22_X1 port map( A1 => io_out1_1_21_port, A2 => n3005, B1 => 
                           loc_out1_0_21_port, B2 => n2999, ZN => n2558);
   U2560 : AOI22_X1 port map( A1 => io_out1_3_21_port, A2 => n3017, B1 => 
                           loc_out1_2_21_port, B2 => n3011, ZN => n2559);
   U2561 : NAND4_X1 port map( A1 => n2549, A2 => n2550, A3 => n2551, A4 => 
                           n2552, ZN => n2548);
   U2562 : AOI22_X1 port map( A1 => io_out1_0_22_port, A2 => n2993, B1 => 
                           loc_out1_3_22_port, B2 => n2987, ZN => n2549);
   U2563 : AOI22_X1 port map( A1 => io_out1_1_22_port, A2 => n3005, B1 => 
                           loc_out1_0_22_port, B2 => n2999, ZN => n2550);
   U2564 : AOI22_X1 port map( A1 => io_out1_3_22_port, A2 => n3017, B1 => 
                           loc_out1_2_22_port, B2 => n3011, ZN => n2551);
   U2565 : NAND4_X1 port map( A1 => n2541, A2 => n2542, A3 => n2543, A4 => 
                           n2544, ZN => n2540);
   U2566 : AOI22_X1 port map( A1 => io_out1_0_23_port, A2 => n2993, B1 => 
                           loc_out1_3_23_port, B2 => n2987, ZN => n2541);
   U2567 : AOI22_X1 port map( A1 => io_out1_1_23_port, A2 => n3005, B1 => 
                           loc_out1_0_23_port, B2 => n2999, ZN => n2542);
   U2568 : AOI22_X1 port map( A1 => io_out1_3_23_port, A2 => n3017, B1 => 
                           loc_out1_2_23_port, B2 => n3011, ZN => n2543);
   U2569 : NAND4_X1 port map( A1 => n2533, A2 => n2534, A3 => n2535, A4 => 
                           n2536, ZN => n2532);
   U2570 : AOI22_X1 port map( A1 => io_out1_0_24_port, A2 => n2993, B1 => 
                           loc_out1_3_24_port, B2 => n2987, ZN => n2533);
   U2571 : AOI22_X1 port map( A1 => io_out1_1_24_port, A2 => n3005, B1 => 
                           loc_out1_0_24_port, B2 => n2999, ZN => n2534);
   U2572 : AOI22_X1 port map( A1 => io_out1_3_24_port, A2 => n3017, B1 => 
                           loc_out1_2_24_port, B2 => n3011, ZN => n2535);
   U2573 : NAND4_X1 port map( A1 => n2525, A2 => n2526, A3 => n2527, A4 => 
                           n2528, ZN => n2524);
   U2574 : AOI22_X1 port map( A1 => io_out1_0_25_port, A2 => n2993, B1 => 
                           loc_out1_3_25_port, B2 => n2987, ZN => n2525);
   U2575 : AOI22_X1 port map( A1 => io_out1_1_25_port, A2 => n3005, B1 => 
                           loc_out1_0_25_port, B2 => n2999, ZN => n2526);
   U2576 : AOI22_X1 port map( A1 => io_out1_3_25_port, A2 => n3017, B1 => 
                           loc_out1_2_25_port, B2 => n3011, ZN => n2527);
   U2577 : NAND4_X1 port map( A1 => n2517, A2 => n2518, A3 => n2519, A4 => 
                           n2520, ZN => n2516);
   U2578 : AOI22_X1 port map( A1 => io_out1_0_26_port, A2 => n2993, B1 => 
                           loc_out1_3_26_port, B2 => n2987, ZN => n2517);
   U2579 : AOI22_X1 port map( A1 => io_out1_1_26_port, A2 => n3005, B1 => 
                           loc_out1_0_26_port, B2 => n2999, ZN => n2518);
   U2580 : AOI22_X1 port map( A1 => io_out1_3_26_port, A2 => n3017, B1 => 
                           loc_out1_2_26_port, B2 => n3011, ZN => n2519);
   U2581 : NAND4_X1 port map( A1 => n2509, A2 => n2510, A3 => n2511, A4 => 
                           n2512, ZN => n2508);
   U2582 : AOI22_X1 port map( A1 => io_out1_0_27_port, A2 => n2993, B1 => 
                           loc_out1_3_27_port, B2 => n2987, ZN => n2509);
   U2583 : AOI22_X1 port map( A1 => io_out1_1_27_port, A2 => n3005, B1 => 
                           loc_out1_0_27_port, B2 => n2999, ZN => n2510);
   U2584 : AOI22_X1 port map( A1 => io_out1_3_27_port, A2 => n3017, B1 => 
                           loc_out1_2_27_port, B2 => n3011, ZN => n2511);
   U2585 : NAND4_X1 port map( A1 => n2501, A2 => n2502, A3 => n2503, A4 => 
                           n2504, ZN => n2500);
   U2586 : AOI22_X1 port map( A1 => io_out1_0_28_port, A2 => n2993, B1 => 
                           loc_out1_3_28_port, B2 => n2987, ZN => n2501);
   U2587 : AOI22_X1 port map( A1 => io_out1_1_28_port, A2 => n3005, B1 => 
                           loc_out1_0_28_port, B2 => n2999, ZN => n2502);
   U2588 : AOI22_X1 port map( A1 => io_out1_3_28_port, A2 => n3017, B1 => 
                           loc_out1_2_28_port, B2 => n3011, ZN => n2503);
   U2589 : NAND4_X1 port map( A1 => n2493, A2 => n2494, A3 => n2495, A4 => 
                           n2496, ZN => n2492);
   U2590 : AOI22_X1 port map( A1 => io_out1_0_29_port, A2 => n2993, B1 => 
                           loc_out1_3_29_port, B2 => n2987, ZN => n2493);
   U2591 : AOI22_X1 port map( A1 => io_out1_1_29_port, A2 => n3005, B1 => 
                           loc_out1_0_29_port, B2 => n2999, ZN => n2494);
   U2592 : AOI22_X1 port map( A1 => io_out1_3_29_port, A2 => n3017, B1 => 
                           loc_out1_2_29_port, B2 => n3011, ZN => n2495);
   U2593 : NAND4_X1 port map( A1 => n2477, A2 => n2478, A3 => n2479, A4 => 
                           n2480, ZN => n2476);
   U2594 : AOI22_X1 port map( A1 => io_out1_0_30_port, A2 => n2993, B1 => 
                           loc_out1_3_30_port, B2 => n2987, ZN => n2477);
   U2595 : AOI22_X1 port map( A1 => io_out1_1_30_port, A2 => n3005, B1 => 
                           loc_out1_0_30_port, B2 => n2999, ZN => n2478);
   U2596 : AOI22_X1 port map( A1 => io_out1_3_30_port, A2 => n3017, B1 => 
                           loc_out1_2_30_port, B2 => n3011, ZN => n2479);
   U2597 : NAND4_X1 port map( A1 => n2469, A2 => n2470, A3 => n2471, A4 => 
                           n2472, ZN => n2468);
   U2598 : AOI22_X1 port map( A1 => io_out1_0_31_port, A2 => n2994, B1 => 
                           loc_out1_3_31_port, B2 => n2988, ZN => n2469);
   U2599 : AOI22_X1 port map( A1 => io_out1_1_31_port, A2 => n3006, B1 => 
                           loc_out1_0_31_port, B2 => n3000, ZN => n2470);
   U2600 : AOI22_X1 port map( A1 => io_out1_3_31_port, A2 => n3018, B1 => 
                           loc_out1_2_31_port, B2 => n3012, ZN => n2471);
   U2601 : NAND4_X1 port map( A1 => n2461, A2 => n2462, A3 => n2463, A4 => 
                           n2464, ZN => n2460);
   U2602 : AOI22_X1 port map( A1 => io_out1_0_32_port, A2 => n2994, B1 => 
                           loc_out1_3_32_port, B2 => n2988, ZN => n2461);
   U2603 : AOI22_X1 port map( A1 => io_out1_1_32_port, A2 => n3006, B1 => 
                           loc_out1_0_32_port, B2 => n3000, ZN => n2462);
   U2604 : AOI22_X1 port map( A1 => io_out1_3_32_port, A2 => n3018, B1 => 
                           loc_out1_2_32_port, B2 => n3012, ZN => n2463);
   U2605 : NAND4_X1 port map( A1 => n2453, A2 => n2454, A3 => n2455, A4 => 
                           n2456, ZN => n2452);
   U2606 : AOI22_X1 port map( A1 => io_out1_0_33_port, A2 => n2994, B1 => 
                           loc_out1_3_33_port, B2 => n2988, ZN => n2453);
   U2607 : AOI22_X1 port map( A1 => io_out1_1_33_port, A2 => n3006, B1 => 
                           loc_out1_0_33_port, B2 => n3000, ZN => n2454);
   U2608 : AOI22_X1 port map( A1 => io_out1_3_33_port, A2 => n3018, B1 => 
                           loc_out1_2_33_port, B2 => n3012, ZN => n2455);
   U2609 : NAND4_X1 port map( A1 => n2445, A2 => n2446, A3 => n2447, A4 => 
                           n2448, ZN => n2444);
   U2610 : AOI22_X1 port map( A1 => io_out1_0_34_port, A2 => n2994, B1 => 
                           loc_out1_3_34_port, B2 => n2988, ZN => n2445);
   U2611 : AOI22_X1 port map( A1 => io_out1_1_34_port, A2 => n3006, B1 => 
                           loc_out1_0_34_port, B2 => n3000, ZN => n2446);
   U2612 : AOI22_X1 port map( A1 => io_out1_3_34_port, A2 => n3018, B1 => 
                           loc_out1_2_34_port, B2 => n3012, ZN => n2447);
   U2613 : NAND4_X1 port map( A1 => n2437, A2 => n2438, A3 => n2439, A4 => 
                           n2440, ZN => n2436);
   U2614 : AOI22_X1 port map( A1 => io_out1_0_35_port, A2 => n2994, B1 => 
                           loc_out1_3_35_port, B2 => n2988, ZN => n2437);
   U2615 : AOI22_X1 port map( A1 => io_out1_1_35_port, A2 => n3006, B1 => 
                           loc_out1_0_35_port, B2 => n3000, ZN => n2438);
   U2616 : AOI22_X1 port map( A1 => io_out1_3_35_port, A2 => n3018, B1 => 
                           loc_out1_2_35_port, B2 => n3012, ZN => n2439);
   U2617 : NAND4_X1 port map( A1 => n2429, A2 => n2430, A3 => n2431, A4 => 
                           n2432, ZN => n2428);
   U2618 : AOI22_X1 port map( A1 => io_out1_0_36_port, A2 => n2994, B1 => 
                           loc_out1_3_36_port, B2 => n2988, ZN => n2429);
   U2619 : AOI22_X1 port map( A1 => io_out1_1_36_port, A2 => n3006, B1 => 
                           loc_out1_0_36_port, B2 => n3000, ZN => n2430);
   U2620 : AOI22_X1 port map( A1 => io_out1_3_36_port, A2 => n3018, B1 => 
                           loc_out1_2_36_port, B2 => n3012, ZN => n2431);
   U2621 : NAND4_X1 port map( A1 => n2421, A2 => n2422, A3 => n2423, A4 => 
                           n2424, ZN => n2420);
   U2622 : AOI22_X1 port map( A1 => io_out1_0_37_port, A2 => n2994, B1 => 
                           loc_out1_3_37_port, B2 => n2988, ZN => n2421);
   U2623 : AOI22_X1 port map( A1 => io_out1_1_37_port, A2 => n3006, B1 => 
                           loc_out1_0_37_port, B2 => n3000, ZN => n2422);
   U2624 : AOI22_X1 port map( A1 => io_out1_3_37_port, A2 => n3018, B1 => 
                           loc_out1_2_37_port, B2 => n3012, ZN => n2423);
   U2625 : NAND4_X1 port map( A1 => n2413, A2 => n2414, A3 => n2415, A4 => 
                           n2416, ZN => n2412);
   U2626 : AOI22_X1 port map( A1 => io_out1_0_38_port, A2 => n2994, B1 => 
                           loc_out1_3_38_port, B2 => n2988, ZN => n2413);
   U2627 : AOI22_X1 port map( A1 => io_out1_1_38_port, A2 => n3006, B1 => 
                           loc_out1_0_38_port, B2 => n3000, ZN => n2414);
   U2628 : AOI22_X1 port map( A1 => io_out1_3_38_port, A2 => n3018, B1 => 
                           loc_out1_2_38_port, B2 => n3012, ZN => n2415);
   U2629 : NAND4_X1 port map( A1 => n2405, A2 => n2406, A3 => n2407, A4 => 
                           n2408, ZN => n2404);
   U2630 : AOI22_X1 port map( A1 => io_out1_0_39_port, A2 => n2994, B1 => 
                           loc_out1_3_39_port, B2 => n2988, ZN => n2405);
   U2631 : AOI22_X1 port map( A1 => io_out1_1_39_port, A2 => n3006, B1 => 
                           loc_out1_0_39_port, B2 => n3000, ZN => n2406);
   U2632 : AOI22_X1 port map( A1 => io_out1_3_39_port, A2 => n3018, B1 => 
                           loc_out1_2_39_port, B2 => n3012, ZN => n2407);
   U2633 : NAND4_X1 port map( A1 => n2389, A2 => n2390, A3 => n2391, A4 => 
                           n2392, ZN => n2388);
   U2634 : AOI22_X1 port map( A1 => io_out1_0_40_port, A2 => n2994, B1 => 
                           loc_out1_3_40_port, B2 => n2988, ZN => n2389);
   U2635 : AOI22_X1 port map( A1 => io_out1_1_40_port, A2 => n3006, B1 => 
                           loc_out1_0_40_port, B2 => n3000, ZN => n2390);
   U2636 : AOI22_X1 port map( A1 => io_out1_3_40_port, A2 => n3018, B1 => 
                           loc_out1_2_40_port, B2 => n3012, ZN => n2391);
   U2637 : NAND4_X1 port map( A1 => n2381, A2 => n2382, A3 => n2383, A4 => 
                           n2384, ZN => n2380);
   U2638 : AOI22_X1 port map( A1 => io_out1_0_41_port, A2 => n2994, B1 => 
                           loc_out1_3_41_port, B2 => n2988, ZN => n2381);
   U2639 : AOI22_X1 port map( A1 => io_out1_1_41_port, A2 => n3006, B1 => 
                           loc_out1_0_41_port, B2 => n3000, ZN => n2382);
   U2640 : AOI22_X1 port map( A1 => io_out1_3_41_port, A2 => n3018, B1 => 
                           loc_out1_2_41_port, B2 => n3012, ZN => n2383);
   U2641 : NAND4_X1 port map( A1 => n2663, A2 => n2664, A3 => n2665, A4 => 
                           n2666, ZN => n2662);
   U2642 : AOI22_X1 port map( A1 => io_out1_0_0_port, A2 => n2992, B1 => 
                           loc_out1_3_0_port, B2 => n2986, ZN => n2663);
   U2643 : AOI22_X1 port map( A1 => io_out1_1_0_port, A2 => n3004, B1 => 
                           loc_out1_0_0_port, B2 => n2998, ZN => n2664);
   U2644 : AOI22_X1 port map( A1 => io_out1_3_0_port, A2 => n3016, B1 => 
                           loc_out1_2_0_port, B2 => n3010, ZN => n2665);
   U2645 : NAND4_X1 port map( A1 => n2573, A2 => n2574, A3 => n2575, A4 => 
                           n2576, ZN => n2572);
   U2646 : AOI22_X1 port map( A1 => io_out1_0_1_port, A2 => n2992, B1 => 
                           loc_out1_3_1_port, B2 => n2986, ZN => n2573);
   U2647 : AOI22_X1 port map( A1 => io_out1_1_1_port, A2 => n3004, B1 => 
                           loc_out1_0_1_port, B2 => n2998, ZN => n2574);
   U2648 : AOI22_X1 port map( A1 => io_out1_3_1_port, A2 => n3016, B1 => 
                           loc_out1_2_1_port, B2 => n3010, ZN => n2575);
   U2649 : NAND4_X1 port map( A1 => n2653, A2 => n2654, A3 => n2655, A4 => 
                           n2656, ZN => n2652);
   U2650 : AOI22_X1 port map( A1 => io_out1_0_10_port, A2 => n2992, B1 => 
                           loc_out1_3_10_port, B2 => n2986, ZN => n2653);
   U2651 : AOI22_X1 port map( A1 => io_out1_1_10_port, A2 => n3004, B1 => 
                           loc_out1_0_10_port, B2 => n2998, ZN => n2654);
   U2652 : AOI22_X1 port map( A1 => io_out1_3_10_port, A2 => n3016, B1 => 
                           loc_out1_2_10_port, B2 => n3010, ZN => n2655);
   U2653 : NAND4_X1 port map( A1 => n2645, A2 => n2646, A3 => n2647, A4 => 
                           n2648, ZN => n2644);
   U2654 : AOI22_X1 port map( A1 => io_out1_0_11_port, A2 => n2992, B1 => 
                           loc_out1_3_11_port, B2 => n2986, ZN => n2645);
   U2655 : AOI22_X1 port map( A1 => io_out1_1_11_port, A2 => n3004, B1 => 
                           loc_out1_0_11_port, B2 => n2998, ZN => n2646);
   U2656 : AOI22_X1 port map( A1 => io_out1_3_11_port, A2 => n3016, B1 => 
                           loc_out1_2_11_port, B2 => n3010, ZN => n2647);
   U2657 : NAND4_X1 port map( A1 => n2637, A2 => n2638, A3 => n2639, A4 => 
                           n2640, ZN => n2636);
   U2658 : AOI22_X1 port map( A1 => io_out1_0_12_port, A2 => n2992, B1 => 
                           loc_out1_3_12_port, B2 => n2986, ZN => n2637);
   U2659 : AOI22_X1 port map( A1 => io_out1_1_12_port, A2 => n3004, B1 => 
                           loc_out1_0_12_port, B2 => n2998, ZN => n2638);
   U2660 : AOI22_X1 port map( A1 => io_out1_3_12_port, A2 => n3016, B1 => 
                           loc_out1_2_12_port, B2 => n3010, ZN => n2639);
   U2661 : NAND4_X1 port map( A1 => n2629, A2 => n2630, A3 => n2631, A4 => 
                           n2632, ZN => n2628);
   U2662 : AOI22_X1 port map( A1 => io_out1_0_13_port, A2 => n2992, B1 => 
                           loc_out1_3_13_port, B2 => n2986, ZN => n2629);
   U2663 : AOI22_X1 port map( A1 => io_out1_1_13_port, A2 => n3004, B1 => 
                           loc_out1_0_13_port, B2 => n2998, ZN => n2630);
   U2664 : AOI22_X1 port map( A1 => io_out1_3_13_port, A2 => n3016, B1 => 
                           loc_out1_2_13_port, B2 => n3010, ZN => n2631);
   U2665 : NAND4_X1 port map( A1 => n2621, A2 => n2622, A3 => n2623, A4 => 
                           n2624, ZN => n2620);
   U2666 : AOI22_X1 port map( A1 => io_out1_0_14_port, A2 => n2992, B1 => 
                           loc_out1_3_14_port, B2 => n2986, ZN => n2621);
   U2667 : AOI22_X1 port map( A1 => io_out1_1_14_port, A2 => n3004, B1 => 
                           loc_out1_0_14_port, B2 => n2998, ZN => n2622);
   U2668 : AOI22_X1 port map( A1 => io_out1_3_14_port, A2 => n3016, B1 => 
                           loc_out1_2_14_port, B2 => n3010, ZN => n2623);
   U2669 : NAND4_X1 port map( A1 => n2613, A2 => n2614, A3 => n2615, A4 => 
                           n2616, ZN => n2612);
   U2670 : AOI22_X1 port map( A1 => io_out1_0_15_port, A2 => n2992, B1 => 
                           loc_out1_3_15_port, B2 => n2986, ZN => n2613);
   U2671 : AOI22_X1 port map( A1 => io_out1_1_15_port, A2 => n3004, B1 => 
                           loc_out1_0_15_port, B2 => n2998, ZN => n2614);
   U2672 : AOI22_X1 port map( A1 => io_out1_3_15_port, A2 => n3016, B1 => 
                           loc_out1_2_15_port, B2 => n3010, ZN => n2615);
   U2673 : NAND4_X1 port map( A1 => n2605, A2 => n2606, A3 => n2607, A4 => 
                           n2608, ZN => n2604);
   U2674 : AOI22_X1 port map( A1 => io_out1_0_16_port, A2 => n2992, B1 => 
                           loc_out1_3_16_port, B2 => n2986, ZN => n2605);
   U2675 : AOI22_X1 port map( A1 => io_out1_1_16_port, A2 => n3004, B1 => 
                           loc_out1_0_16_port, B2 => n2998, ZN => n2606);
   U2676 : AOI22_X1 port map( A1 => io_out1_3_16_port, A2 => n3016, B1 => 
                           loc_out1_2_16_port, B2 => n3010, ZN => n2607);
   U2677 : NAND4_X1 port map( A1 => n2597, A2 => n2598, A3 => n2599, A4 => 
                           n2600, ZN => n2596);
   U2678 : AOI22_X1 port map( A1 => io_out1_0_17_port, A2 => n2992, B1 => 
                           loc_out1_3_17_port, B2 => n2986, ZN => n2597);
   U2679 : AOI22_X1 port map( A1 => io_out1_1_17_port, A2 => n3004, B1 => 
                           loc_out1_0_17_port, B2 => n2998, ZN => n2598);
   U2680 : AOI22_X1 port map( A1 => io_out1_3_17_port, A2 => n3016, B1 => 
                           loc_out1_2_17_port, B2 => n3010, ZN => n2599);
   U2681 : NAND4_X1 port map( A1 => n2589, A2 => n2590, A3 => n2591, A4 => 
                           n2592, ZN => n2588);
   U2682 : AOI22_X1 port map( A1 => io_out1_0_18_port, A2 => n2992, B1 => 
                           loc_out1_3_18_port, B2 => n2986, ZN => n2589);
   U2683 : AOI22_X1 port map( A1 => io_out1_1_18_port, A2 => n3004, B1 => 
                           loc_out1_0_18_port, B2 => n2998, ZN => n2590);
   U2684 : AOI22_X1 port map( A1 => io_out1_3_18_port, A2 => n3016, B1 => 
                           loc_out1_2_18_port, B2 => n3010, ZN => n2591);
   U2685 : NAND4_X1 port map( A1 => n2581, A2 => n2582, A3 => n2583, A4 => 
                           n2584, ZN => n2580);
   U2686 : AOI22_X1 port map( A1 => io_out1_0_19_port, A2 => n2992, B1 => 
                           loc_out1_3_19_port, B2 => n2986, ZN => n2581);
   U2687 : AOI22_X1 port map( A1 => io_out1_1_19_port, A2 => n3004, B1 => 
                           loc_out1_0_19_port, B2 => n2998, ZN => n2582);
   U2688 : AOI22_X1 port map( A1 => io_out1_3_19_port, A2 => n3016, B1 => 
                           loc_out1_2_19_port, B2 => n3010, ZN => n2583);
   U2689 : AND3_X1 port map( A1 => ADD_RD2(2), A2 => ADD_RD2(3), A3 => RD2, ZN 
                           => global_read2);
   U2690 : INV_X1 port map( A => RD1, ZN => n2119);
   U2691 : OAI211_X1 port map( C1 => n3074, C2 => n2658, A => n2659, B => n2660
                           , ZN => OUT1(0));
   U2692 : INV_X1 port map( A => global_out1_0_port, ZN => n2658);
   U2693 : AOI22_X1 port map( A1 => n3046, A2 => n2662, B1 => io_out1_2_0_port,
                           B2 => n3052, ZN => n2659);
   U2694 : AOI222_X1 port map( A1 => io_out1_3_0_port, A2 => n3063, B1 => 
                           io_out1_1_0_port, B2 => n3045, C1 => 
                           io_out1_0_0_port, C2 => n2657, ZN => n2660);
   U2695 : OAI211_X1 port map( C1 => n3066, C2 => n2217, A => n2218, B => n2219
                           , ZN => OUT1(5));
   U2696 : INV_X1 port map( A => io_out1_0_5_port, ZN => n2217);
   U2697 : AOI22_X1 port map( A1 => n3050, A2 => n2220, B1 => io_out1_1_5_port,
                           B2 => n3040, ZN => n2218);
   U2698 : AOI222_X1 port map( A1 => global_out1_5_port, A2 => n3072, B1 => 
                           io_out1_3_5_port, B2 => n3058, C1 => 
                           io_out1_2_5_port, C2 => n3056, ZN => n2219);
   U2699 : OAI211_X1 port map( C1 => n3066, C2 => n2177, A => n2178, B => n2179
                           , ZN => OUT1(6));
   U2700 : INV_X1 port map( A => io_out1_0_6_port, ZN => n2177);
   U2701 : AOI22_X1 port map( A1 => n3051, A2 => n2180, B1 => io_out1_1_6_port,
                           B2 => n3040, ZN => n2178);
   U2702 : AOI222_X1 port map( A1 => global_out1_6_port, A2 => n3073, B1 => 
                           io_out1_3_6_port, B2 => n3058, C1 => 
                           io_out1_2_6_port, C2 => n3057, ZN => n2179);
   U2703 : OAI211_X1 port map( C1 => n3066, C2 => n2169, A => n2170, B => n2171
                           , ZN => OUT1(7));
   U2704 : INV_X1 port map( A => io_out1_0_7_port, ZN => n2169);
   U2705 : AOI22_X1 port map( A1 => n3051, A2 => n2172, B1 => io_out1_1_7_port,
                           B2 => n3040, ZN => n2170);
   U2706 : AOI222_X1 port map( A1 => global_out1_7_port, A2 => n3071, B1 => 
                           io_out1_3_7_port, B2 => n3058, C1 => 
                           io_out1_2_7_port, C2 => n3057, ZN => n2171);
   U2707 : OAI211_X1 port map( C1 => n3066, C2 => n2161, A => n2162, B => n2163
                           , ZN => OUT1(8));
   U2708 : INV_X1 port map( A => io_out1_0_8_port, ZN => n2161);
   U2709 : AOI22_X1 port map( A1 => n3051, A2 => n2164, B1 => io_out1_1_8_port,
                           B2 => n3040, ZN => n2162);
   U2710 : AOI222_X1 port map( A1 => global_out1_8_port, A2 => n3072, B1 => 
                           io_out1_3_8_port, B2 => n3058, C1 => 
                           io_out1_2_8_port, C2 => n3057, ZN => n2163);
   U2711 : OAI211_X1 port map( C1 => n3066, C2 => n2249, A => n2250, B => n2251
                           , ZN => OUT1(56));
   U2712 : INV_X1 port map( A => io_out1_0_56_port, ZN => n2249);
   U2713 : AOI22_X1 port map( A1 => n3050, A2 => n2252, B1 => io_out1_1_56_port
                           , B2 => n3040, ZN => n2250);
   U2714 : AOI222_X1 port map( A1 => global_out1_56_port, A2 => n3071, B1 => 
                           io_out1_3_56_port, B2 => n3058, C1 => 
                           io_out1_2_56_port, C2 => n3056, ZN => n2251);
   U2715 : OAI211_X1 port map( C1 => n3066, C2 => n2241, A => n2242, B => n2243
                           , ZN => OUT1(57));
   U2716 : INV_X1 port map( A => io_out1_0_57_port, ZN => n2241);
   U2717 : AOI22_X1 port map( A1 => n3050, A2 => n2244, B1 => io_out1_1_57_port
                           , B2 => n3040, ZN => n2242);
   U2718 : AOI222_X1 port map( A1 => global_out1_57_port, A2 => n3073, B1 => 
                           io_out1_3_57_port, B2 => n3058, C1 => 
                           io_out1_2_57_port, C2 => n3056, ZN => n2243);
   U2719 : OAI211_X1 port map( C1 => n3066, C2 => n2233, A => n2234, B => n2235
                           , ZN => OUT1(58));
   U2720 : INV_X1 port map( A => io_out1_0_58_port, ZN => n2233);
   U2721 : AOI22_X1 port map( A1 => n3050, A2 => n2236, B1 => io_out1_1_58_port
                           , B2 => n3040, ZN => n2234);
   U2722 : AOI222_X1 port map( A1 => global_out1_58_port, A2 => n3071, B1 => 
                           io_out1_3_58_port, B2 => n3058, C1 => 
                           io_out1_2_58_port, C2 => n3056, ZN => n2235);
   U2723 : OAI211_X1 port map( C1 => n3066, C2 => n2225, A => n2226, B => n2227
                           , ZN => OUT1(59));
   U2724 : INV_X1 port map( A => io_out1_0_59_port, ZN => n2225);
   U2725 : AOI22_X1 port map( A1 => n3050, A2 => n2228, B1 => io_out1_1_59_port
                           , B2 => n3040, ZN => n2226);
   U2726 : AOI222_X1 port map( A1 => global_out1_59_port, A2 => n3072, B1 => 
                           io_out1_3_59_port, B2 => n3058, C1 => 
                           io_out1_2_59_port, C2 => n3056, ZN => n2227);
   U2727 : OAI211_X1 port map( C1 => n3066, C2 => n2209, A => n2210, B => n2211
                           , ZN => OUT1(60));
   U2728 : INV_X1 port map( A => io_out1_0_60_port, ZN => n2209);
   U2729 : AOI22_X1 port map( A1 => n3050, A2 => n2212, B1 => io_out1_1_60_port
                           , B2 => n3040, ZN => n2210);
   U2730 : AOI222_X1 port map( A1 => global_out1_60_port, A2 => n3073, B1 => 
                           io_out1_3_60_port, B2 => n3058, C1 => 
                           io_out1_2_60_port, C2 => n3056, ZN => n2211);
   U2731 : OAI211_X1 port map( C1 => n3066, C2 => n2201, A => n2202, B => n2203
                           , ZN => OUT1(61));
   U2732 : INV_X1 port map( A => io_out1_0_61_port, ZN => n2201);
   U2733 : AOI22_X1 port map( A1 => n3050, A2 => n2204, B1 => io_out1_1_61_port
                           , B2 => n3040, ZN => n2202);
   U2734 : AOI222_X1 port map( A1 => global_out1_61_port, A2 => n3071, B1 => 
                           io_out1_3_61_port, B2 => n3058, C1 => 
                           io_out1_2_61_port, C2 => n3056, ZN => n2203);
   U2735 : OAI211_X1 port map( C1 => n3066, C2 => n2193, A => n2194, B => n2195
                           , ZN => OUT1(62));
   U2736 : INV_X1 port map( A => io_out1_0_62_port, ZN => n2193);
   U2737 : AOI22_X1 port map( A1 => n3050, A2 => n2196, B1 => io_out1_1_62_port
                           , B2 => n3040, ZN => n2194);
   U2738 : AOI222_X1 port map( A1 => global_out1_62_port, A2 => n3072, B1 => 
                           io_out1_3_62_port, B2 => n3058, C1 => 
                           io_out1_2_62_port, C2 => n3056, ZN => n2195);
   U2739 : OAI211_X1 port map( C1 => n3066, C2 => n2185, A => n2186, B => n2187
                           , ZN => OUT1(63));
   U2740 : INV_X1 port map( A => io_out1_0_63_port, ZN => n2185);
   U2741 : AOI22_X1 port map( A1 => n3050, A2 => n2188, B1 => io_out1_1_63_port
                           , B2 => n3040, ZN => n2186);
   U2742 : AOI222_X1 port map( A1 => global_out1_63_port, A2 => n3073, B1 => 
                           io_out1_3_63_port, B2 => n3058, C1 => 
                           io_out1_2_63_port, C2 => n3056, ZN => n2187);
   U2743 : OAI211_X1 port map( C1 => n3069, C2 => n2481, A => n2482, B => n2483
                           , ZN => OUT1(2));
   U2744 : INV_X1 port map( A => io_out1_0_2_port, ZN => n2481);
   U2745 : AOI22_X1 port map( A1 => n3047, A2 => n2484, B1 => io_out1_1_2_port,
                           B2 => n3043, ZN => n2482);
   U2746 : AOI222_X1 port map( A1 => global_out1_2_port, A2 => n3073, B1 => 
                           io_out1_3_2_port, B2 => n3061, C1 => 
                           io_out1_2_2_port, C2 => n3053, ZN => n2483);
   U2747 : OAI211_X1 port map( C1 => n3068, C2 => n2393, A => n2394, B => n2395
                           , ZN => OUT1(3));
   U2748 : INV_X1 port map( A => io_out1_0_3_port, ZN => n2393);
   U2749 : AOI22_X1 port map( A1 => n3048, A2 => n2396, B1 => io_out1_1_3_port,
                           B2 => n3042, ZN => n2394);
   U2750 : AOI222_X1 port map( A1 => global_out1_3_port, A2 => n3072, B1 => 
                           io_out1_3_3_port, B2 => n3060, C1 => 
                           io_out1_2_3_port, C2 => n3054, ZN => n2395);
   U2751 : OAI211_X1 port map( C1 => n3067, C2 => n2305, A => n2306, B => n2307
                           , ZN => OUT1(4));
   U2752 : INV_X1 port map( A => io_out1_0_4_port, ZN => n2305);
   U2753 : AOI22_X1 port map( A1 => n3049, A2 => n2308, B1 => io_out1_1_4_port,
                           B2 => n3041, ZN => n2306);
   U2754 : AOI222_X1 port map( A1 => global_out1_4_port, A2 => n3071, B1 => 
                           io_out1_3_4_port, B2 => n3059, C1 => 
                           io_out1_2_4_port, C2 => n3055, ZN => n2307);
   U2755 : OAI211_X1 port map( C1 => n3069, C2 => n2561, A => n2562, B => n2563
                           , ZN => OUT1(20));
   U2756 : INV_X1 port map( A => io_out1_0_20_port, ZN => n2561);
   U2757 : AOI22_X1 port map( A1 => n3047, A2 => n2564, B1 => io_out1_1_20_port
                           , B2 => n3044, ZN => n2562);
   U2758 : AOI222_X1 port map( A1 => global_out1_20_port, A2 => n3071, B1 => 
                           io_out1_3_20_port, B2 => n3062, C1 => 
                           io_out1_2_20_port, C2 => n3053, ZN => n2563);
   U2759 : OAI211_X1 port map( C1 => n3069, C2 => n2553, A => n2554, B => n2555
                           , ZN => OUT1(21));
   U2760 : INV_X1 port map( A => io_out1_0_21_port, ZN => n2553);
   U2761 : AOI22_X1 port map( A1 => n3047, A2 => n2556, B1 => io_out1_1_21_port
                           , B2 => n3044, ZN => n2554);
   U2762 : AOI222_X1 port map( A1 => global_out1_21_port, A2 => n3073, B1 => 
                           io_out1_3_21_port, B2 => n3062, C1 => 
                           io_out1_2_21_port, C2 => n3053, ZN => n2555);
   U2763 : OAI211_X1 port map( C1 => n3069, C2 => n2545, A => n2546, B => n2547
                           , ZN => OUT1(22));
   U2764 : INV_X1 port map( A => io_out1_0_22_port, ZN => n2545);
   U2765 : AOI22_X1 port map( A1 => n3047, A2 => n2548, B1 => io_out1_1_22_port
                           , B2 => n3043, ZN => n2546);
   U2766 : AOI222_X1 port map( A1 => global_out1_22_port, A2 => n3071, B1 => 
                           io_out1_3_22_port, B2 => n3061, C1 => 
                           io_out1_2_22_port, C2 => n3053, ZN => n2547);
   U2767 : OAI211_X1 port map( C1 => n3069, C2 => n2537, A => n2538, B => n2539
                           , ZN => OUT1(23));
   U2768 : INV_X1 port map( A => io_out1_0_23_port, ZN => n2537);
   U2769 : AOI22_X1 port map( A1 => n3047, A2 => n2540, B1 => io_out1_1_23_port
                           , B2 => n3044, ZN => n2538);
   U2770 : AOI222_X1 port map( A1 => global_out1_23_port, A2 => n3073, B1 => 
                           io_out1_3_23_port, B2 => n3062, C1 => 
                           io_out1_2_23_port, C2 => n3053, ZN => n2539);
   U2771 : OAI211_X1 port map( C1 => n3069, C2 => n2529, A => n2530, B => n2531
                           , ZN => OUT1(24));
   U2772 : INV_X1 port map( A => io_out1_0_24_port, ZN => n2529);
   U2773 : AOI22_X1 port map( A1 => n3047, A2 => n2532, B1 => io_out1_1_24_port
                           , B2 => n3043, ZN => n2530);
   U2774 : AOI222_X1 port map( A1 => global_out1_24_port, A2 => n3073, B1 => 
                           io_out1_3_24_port, B2 => n3061, C1 => 
                           io_out1_2_24_port, C2 => n3053, ZN => n2531);
   U2775 : OAI211_X1 port map( C1 => n3069, C2 => n2521, A => n2522, B => n2523
                           , ZN => OUT1(25));
   U2776 : INV_X1 port map( A => io_out1_0_25_port, ZN => n2521);
   U2777 : AOI22_X1 port map( A1 => n3047, A2 => n2524, B1 => io_out1_1_25_port
                           , B2 => n3043, ZN => n2522);
   U2778 : AOI222_X1 port map( A1 => global_out1_25_port, A2 => n3073, B1 => 
                           io_out1_3_25_port, B2 => n3061, C1 => 
                           io_out1_2_25_port, C2 => n3053, ZN => n2523);
   U2779 : OAI211_X1 port map( C1 => n3069, C2 => n2513, A => n2514, B => n2515
                           , ZN => OUT1(26));
   U2780 : INV_X1 port map( A => io_out1_0_26_port, ZN => n2513);
   U2781 : AOI22_X1 port map( A1 => n3047, A2 => n2516, B1 => io_out1_1_26_port
                           , B2 => n3043, ZN => n2514);
   U2782 : AOI222_X1 port map( A1 => global_out1_26_port, A2 => n3073, B1 => 
                           io_out1_3_26_port, B2 => n3061, C1 => 
                           io_out1_2_26_port, C2 => n3053, ZN => n2515);
   U2783 : OAI211_X1 port map( C1 => n3069, C2 => n2505, A => n2506, B => n2507
                           , ZN => OUT1(27));
   U2784 : INV_X1 port map( A => io_out1_0_27_port, ZN => n2505);
   U2785 : AOI22_X1 port map( A1 => n3047, A2 => n2508, B1 => io_out1_1_27_port
                           , B2 => n3043, ZN => n2506);
   U2786 : AOI222_X1 port map( A1 => global_out1_27_port, A2 => n3073, B1 => 
                           io_out1_3_27_port, B2 => n3061, C1 => 
                           io_out1_2_27_port, C2 => n3053, ZN => n2507);
   U2787 : OAI211_X1 port map( C1 => n3069, C2 => n2497, A => n2498, B => n2499
                           , ZN => OUT1(28));
   U2788 : INV_X1 port map( A => io_out1_0_28_port, ZN => n2497);
   U2789 : AOI22_X1 port map( A1 => n3047, A2 => n2500, B1 => io_out1_1_28_port
                           , B2 => n3043, ZN => n2498);
   U2790 : AOI222_X1 port map( A1 => global_out1_28_port, A2 => n3073, B1 => 
                           io_out1_3_28_port, B2 => n3061, C1 => 
                           io_out1_2_28_port, C2 => n3053, ZN => n2499);
   U2791 : OAI211_X1 port map( C1 => n3069, C2 => n2489, A => n2490, B => n2491
                           , ZN => OUT1(29));
   U2792 : INV_X1 port map( A => io_out1_0_29_port, ZN => n2489);
   U2793 : AOI22_X1 port map( A1 => n3047, A2 => n2492, B1 => io_out1_1_29_port
                           , B2 => n3043, ZN => n2490);
   U2794 : AOI222_X1 port map( A1 => global_out1_29_port, A2 => n3073, B1 => 
                           io_out1_3_29_port, B2 => n3061, C1 => 
                           io_out1_2_29_port, C2 => n3053, ZN => n2491);
   U2795 : OAI211_X1 port map( C1 => n3069, C2 => n2473, A => n2474, B => n2475
                           , ZN => OUT1(30));
   U2796 : INV_X1 port map( A => io_out1_0_30_port, ZN => n2473);
   U2797 : AOI22_X1 port map( A1 => n3047, A2 => n2476, B1 => io_out1_1_30_port
                           , B2 => n3043, ZN => n2474);
   U2798 : AOI222_X1 port map( A1 => global_out1_30_port, A2 => n3073, B1 => 
                           io_out1_3_30_port, B2 => n3061, C1 => 
                           io_out1_2_30_port, C2 => n3053, ZN => n2475);
   U2799 : OAI211_X1 port map( C1 => n3068, C2 => n2441, A => n2442, B => n2443
                           , ZN => OUT1(34));
   U2800 : INV_X1 port map( A => io_out1_0_34_port, ZN => n2441);
   U2801 : AOI22_X1 port map( A1 => n3048, A2 => n2444, B1 => io_out1_1_34_port
                           , B2 => n3042, ZN => n2442);
   U2802 : AOI222_X1 port map( A1 => global_out1_34_port, A2 => n3073, B1 => 
                           io_out1_3_34_port, B2 => n3060, C1 => 
                           io_out1_2_34_port, C2 => n3054, ZN => n2443);
   U2803 : OAI211_X1 port map( C1 => n3068, C2 => n2433, A => n2434, B => n2435
                           , ZN => OUT1(35));
   U2804 : INV_X1 port map( A => io_out1_0_35_port, ZN => n2433);
   U2805 : AOI22_X1 port map( A1 => n3048, A2 => n2436, B1 => io_out1_1_35_port
                           , B2 => n3042, ZN => n2434);
   U2806 : AOI222_X1 port map( A1 => global_out1_35_port, A2 => n3072, B1 => 
                           io_out1_3_35_port, B2 => n3060, C1 => 
                           io_out1_2_35_port, C2 => n3054, ZN => n2435);
   U2807 : OAI211_X1 port map( C1 => n3068, C2 => n2425, A => n2426, B => n2427
                           , ZN => OUT1(36));
   U2808 : INV_X1 port map( A => io_out1_0_36_port, ZN => n2425);
   U2809 : AOI22_X1 port map( A1 => n3048, A2 => n2428, B1 => io_out1_1_36_port
                           , B2 => n3042, ZN => n2426);
   U2810 : AOI222_X1 port map( A1 => global_out1_36_port, A2 => n3072, B1 => 
                           io_out1_3_36_port, B2 => n3060, C1 => 
                           io_out1_2_36_port, C2 => n3054, ZN => n2427);
   U2811 : OAI211_X1 port map( C1 => n3068, C2 => n2417, A => n2418, B => n2419
                           , ZN => OUT1(37));
   U2812 : INV_X1 port map( A => io_out1_0_37_port, ZN => n2417);
   U2813 : AOI22_X1 port map( A1 => n3048, A2 => n2420, B1 => io_out1_1_37_port
                           , B2 => n3042, ZN => n2418);
   U2814 : AOI222_X1 port map( A1 => global_out1_37_port, A2 => n3072, B1 => 
                           io_out1_3_37_port, B2 => n3060, C1 => 
                           io_out1_2_37_port, C2 => n3054, ZN => n2419);
   U2815 : OAI211_X1 port map( C1 => n3068, C2 => n2409, A => n2410, B => n2411
                           , ZN => OUT1(38));
   U2816 : INV_X1 port map( A => io_out1_0_38_port, ZN => n2409);
   U2817 : AOI22_X1 port map( A1 => n3048, A2 => n2412, B1 => io_out1_1_38_port
                           , B2 => n3042, ZN => n2410);
   U2818 : AOI222_X1 port map( A1 => global_out1_38_port, A2 => n3072, B1 => 
                           io_out1_3_38_port, B2 => n3060, C1 => 
                           io_out1_2_38_port, C2 => n3054, ZN => n2411);
   U2819 : OAI211_X1 port map( C1 => n3068, C2 => n2401, A => n2402, B => n2403
                           , ZN => OUT1(39));
   U2820 : INV_X1 port map( A => io_out1_0_39_port, ZN => n2401);
   U2821 : AOI22_X1 port map( A1 => n3048, A2 => n2404, B1 => io_out1_1_39_port
                           , B2 => n3042, ZN => n2402);
   U2822 : AOI222_X1 port map( A1 => global_out1_39_port, A2 => n3072, B1 => 
                           io_out1_3_39_port, B2 => n3060, C1 => 
                           io_out1_2_39_port, C2 => n3054, ZN => n2403);
   U2823 : OAI211_X1 port map( C1 => n3068, C2 => n2385, A => n2386, B => n2387
                           , ZN => OUT1(40));
   U2824 : INV_X1 port map( A => io_out1_0_40_port, ZN => n2385);
   U2825 : AOI22_X1 port map( A1 => n3048, A2 => n2388, B1 => io_out1_1_40_port
                           , B2 => n3042, ZN => n2386);
   U2826 : AOI222_X1 port map( A1 => global_out1_40_port, A2 => n3072, B1 => 
                           io_out1_3_40_port, B2 => n3060, C1 => 
                           io_out1_2_40_port, C2 => n3054, ZN => n2387);
   U2827 : OAI211_X1 port map( C1 => n3068, C2 => n2377, A => n2378, B => n2379
                           , ZN => OUT1(41));
   U2828 : INV_X1 port map( A => io_out1_0_41_port, ZN => n2377);
   U2829 : AOI22_X1 port map( A1 => n3048, A2 => n2380, B1 => io_out1_1_41_port
                           , B2 => n3042, ZN => n2378);
   U2830 : AOI222_X1 port map( A1 => global_out1_41_port, A2 => n3072, B1 => 
                           io_out1_3_41_port, B2 => n3060, C1 => 
                           io_out1_2_41_port, C2 => n3054, ZN => n2379);
   U2831 : OAI211_X1 port map( C1 => n3068, C2 => n2369, A => n2370, B => n2371
                           , ZN => OUT1(42));
   U2832 : INV_X1 port map( A => io_out1_0_42_port, ZN => n2369);
   U2833 : AOI22_X1 port map( A1 => n3049, A2 => n2372, B1 => io_out1_1_42_port
                           , B2 => n3042, ZN => n2370);
   U2834 : AOI222_X1 port map( A1 => global_out1_42_port, A2 => n3072, B1 => 
                           io_out1_3_42_port, B2 => n3060, C1 => 
                           io_out1_2_42_port, C2 => n3055, ZN => n2371);
   U2835 : OAI211_X1 port map( C1 => n3068, C2 => n2361, A => n2362, B => n2363
                           , ZN => OUT1(43));
   U2836 : INV_X1 port map( A => io_out1_0_43_port, ZN => n2361);
   U2837 : AOI22_X1 port map( A1 => n3049, A2 => n2364, B1 => io_out1_1_43_port
                           , B2 => n3042, ZN => n2362);
   U2838 : AOI222_X1 port map( A1 => global_out1_43_port, A2 => n3072, B1 => 
                           io_out1_3_43_port, B2 => n3060, C1 => 
                           io_out1_2_43_port, C2 => n3055, ZN => n2363);
   U2839 : OAI211_X1 port map( C1 => n3067, C2 => n2353, A => n2354, B => n2355
                           , ZN => OUT1(44));
   U2840 : INV_X1 port map( A => io_out1_0_44_port, ZN => n2353);
   U2841 : AOI22_X1 port map( A1 => n3049, A2 => n2356, B1 => io_out1_1_44_port
                           , B2 => n3041, ZN => n2354);
   U2842 : AOI222_X1 port map( A1 => global_out1_44_port, A2 => n3072, B1 => 
                           io_out1_3_44_port, B2 => n3059, C1 => 
                           io_out1_2_44_port, C2 => n3055, ZN => n2355);
   U2843 : OAI211_X1 port map( C1 => n3067, C2 => n2345, A => n2346, B => n2347
                           , ZN => OUT1(45));
   U2844 : INV_X1 port map( A => io_out1_0_45_port, ZN => n2345);
   U2845 : AOI22_X1 port map( A1 => n3049, A2 => n2348, B1 => io_out1_1_45_port
                           , B2 => n3041, ZN => n2346);
   U2846 : AOI222_X1 port map( A1 => global_out1_45_port, A2 => n3072, B1 => 
                           io_out1_3_45_port, B2 => n3059, C1 => 
                           io_out1_2_45_port, C2 => n3055, ZN => n2347);
   U2847 : OAI211_X1 port map( C1 => n3067, C2 => n2337, A => n2338, B => n2339
                           , ZN => OUT1(46));
   U2848 : INV_X1 port map( A => io_out1_0_46_port, ZN => n2337);
   U2849 : AOI22_X1 port map( A1 => n3049, A2 => n2340, B1 => io_out1_1_46_port
                           , B2 => n3041, ZN => n2338);
   U2850 : AOI222_X1 port map( A1 => global_out1_46_port, A2 => n3071, B1 => 
                           io_out1_3_46_port, B2 => n3059, C1 => 
                           io_out1_2_46_port, C2 => n3055, ZN => n2339);
   U2851 : OAI211_X1 port map( C1 => n3067, C2 => n2329, A => n2330, B => n2331
                           , ZN => OUT1(47));
   U2852 : INV_X1 port map( A => io_out1_0_47_port, ZN => n2329);
   U2853 : AOI22_X1 port map( A1 => n3049, A2 => n2332, B1 => io_out1_1_47_port
                           , B2 => n3041, ZN => n2330);
   U2854 : AOI222_X1 port map( A1 => global_out1_47_port, A2 => n3071, B1 => 
                           io_out1_3_47_port, B2 => n3059, C1 => 
                           io_out1_2_47_port, C2 => n3055, ZN => n2331);
   U2855 : OAI211_X1 port map( C1 => n3067, C2 => n2321, A => n2322, B => n2323
                           , ZN => OUT1(48));
   U2856 : INV_X1 port map( A => io_out1_0_48_port, ZN => n2321);
   U2857 : AOI22_X1 port map( A1 => n3049, A2 => n2324, B1 => io_out1_1_48_port
                           , B2 => n3041, ZN => n2322);
   U2858 : AOI222_X1 port map( A1 => global_out1_48_port, A2 => n3071, B1 => 
                           io_out1_3_48_port, B2 => n3059, C1 => 
                           io_out1_2_48_port, C2 => n3055, ZN => n2323);
   U2859 : OAI211_X1 port map( C1 => n3067, C2 => n2313, A => n2314, B => n2315
                           , ZN => OUT1(49));
   U2860 : INV_X1 port map( A => io_out1_0_49_port, ZN => n2313);
   U2861 : AOI22_X1 port map( A1 => n3049, A2 => n2316, B1 => io_out1_1_49_port
                           , B2 => n3041, ZN => n2314);
   U2862 : AOI222_X1 port map( A1 => global_out1_49_port, A2 => n3071, B1 => 
                           io_out1_3_49_port, B2 => n3059, C1 => 
                           io_out1_2_49_port, C2 => n3055, ZN => n2315);
   U2863 : OAI211_X1 port map( C1 => n3067, C2 => n2297, A => n2298, B => n2299
                           , ZN => OUT1(50));
   U2864 : INV_X1 port map( A => io_out1_0_50_port, ZN => n2297);
   U2865 : AOI22_X1 port map( A1 => n3049, A2 => n2300, B1 => io_out1_1_50_port
                           , B2 => n3041, ZN => n2298);
   U2866 : AOI222_X1 port map( A1 => global_out1_50_port, A2 => n3071, B1 => 
                           io_out1_3_50_port, B2 => n3059, C1 => 
                           io_out1_2_50_port, C2 => n3055, ZN => n2299);
   U2867 : OAI211_X1 port map( C1 => n3067, C2 => n2289, A => n2290, B => n2291
                           , ZN => OUT1(51));
   U2868 : INV_X1 port map( A => io_out1_0_51_port, ZN => n2289);
   U2869 : AOI22_X1 port map( A1 => n3049, A2 => n2292, B1 => io_out1_1_51_port
                           , B2 => n3041, ZN => n2290);
   U2870 : AOI222_X1 port map( A1 => global_out1_51_port, A2 => n3071, B1 => 
                           io_out1_3_51_port, B2 => n3059, C1 => 
                           io_out1_2_51_port, C2 => n3055, ZN => n2291);
   U2871 : OAI211_X1 port map( C1 => n3067, C2 => n2281, A => n2282, B => n2283
                           , ZN => OUT1(52));
   U2872 : INV_X1 port map( A => io_out1_0_52_port, ZN => n2281);
   U2873 : AOI22_X1 port map( A1 => n3049, A2 => n2284, B1 => io_out1_1_52_port
                           , B2 => n3042, ZN => n2282);
   U2874 : AOI222_X1 port map( A1 => global_out1_52_port, A2 => n3071, B1 => 
                           io_out1_3_52_port, B2 => n3060, C1 => 
                           io_out1_2_52_port, C2 => n3055, ZN => n2283);
   U2875 : OAI211_X1 port map( C1 => n3067, C2 => n2273, A => n2274, B => n2275
                           , ZN => OUT1(53));
   U2876 : INV_X1 port map( A => io_out1_0_53_port, ZN => n2273);
   U2877 : AOI22_X1 port map( A1 => n3050, A2 => n2276, B1 => io_out1_1_53_port
                           , B2 => n3041, ZN => n2274);
   U2878 : AOI222_X1 port map( A1 => global_out1_53_port, A2 => n3071, B1 => 
                           io_out1_3_53_port, B2 => n3059, C1 => 
                           io_out1_2_53_port, C2 => n3056, ZN => n2275);
   U2879 : OAI211_X1 port map( C1 => n3067, C2 => n2265, A => n2266, B => n2267
                           , ZN => OUT1(54));
   U2880 : INV_X1 port map( A => io_out1_0_54_port, ZN => n2265);
   U2881 : AOI22_X1 port map( A1 => n3050, A2 => n2268, B1 => io_out1_1_54_port
                           , B2 => n3041, ZN => n2266);
   U2882 : AOI222_X1 port map( A1 => global_out1_54_port, A2 => n3071, B1 => 
                           io_out1_3_54_port, B2 => n3059, C1 => 
                           io_out1_2_54_port, C2 => n3056, ZN => n2267);
   U2883 : OAI211_X1 port map( C1 => n3067, C2 => n2257, A => n2258, B => n2259
                           , ZN => OUT1(55));
   U2884 : INV_X1 port map( A => io_out1_0_55_port, ZN => n2257);
   U2885 : AOI22_X1 port map( A1 => n3050, A2 => n2260, B1 => io_out1_1_55_port
                           , B2 => n3041, ZN => n2258);
   U2886 : AOI222_X1 port map( A1 => global_out1_55_port, A2 => n3071, B1 => 
                           io_out1_3_55_port, B2 => n3059, C1 => 
                           io_out1_2_55_port, C2 => n3056, ZN => n2259);
   U2887 : OAI211_X1 port map( C1 => n3070, C2 => n2569, A => n2570, B => n2571
                           , ZN => OUT1(1));
   U2888 : INV_X1 port map( A => io_out1_0_1_port, ZN => n2569);
   U2889 : AOI22_X1 port map( A1 => n3046, A2 => n2572, B1 => io_out1_1_1_port,
                           B2 => n3044, ZN => n2570);
   U2890 : AOI222_X1 port map( A1 => global_out1_1_port, A2 => n3071, B1 => 
                           io_out1_3_1_port, B2 => n3062, C1 => 
                           io_out1_2_1_port, C2 => n3052, ZN => n2571);
   U2891 : OAI211_X1 port map( C1 => n3070, C2 => n2641, A => n2642, B => n2643
                           , ZN => OUT1(11));
   U2892 : INV_X1 port map( A => io_out1_0_11_port, ZN => n2641);
   U2893 : AOI22_X1 port map( A1 => n3046, A2 => n2644, B1 => io_out1_1_11_port
                           , B2 => n3044, ZN => n2642);
   U2894 : AOI222_X1 port map( A1 => global_out1_11_port, A2 => n3072, B1 => 
                           io_out1_3_11_port, B2 => n3062, C1 => 
                           io_out1_2_11_port, C2 => n3052, ZN => n2643);
   U2895 : OAI211_X1 port map( C1 => n3070, C2 => n2625, A => n2626, B => n2627
                           , ZN => OUT1(13));
   U2896 : INV_X1 port map( A => io_out1_0_13_port, ZN => n2625);
   U2897 : AOI22_X1 port map( A1 => n3046, A2 => n2628, B1 => io_out1_1_13_port
                           , B2 => n3044, ZN => n2626);
   U2898 : AOI222_X1 port map( A1 => global_out1_13_port, A2 => n3073, B1 => 
                           io_out1_3_13_port, B2 => n3062, C1 => 
                           io_out1_2_13_port, C2 => n3052, ZN => n2627);
   U2899 : OAI211_X1 port map( C1 => n3070, C2 => n2617, A => n2618, B => n2619
                           , ZN => OUT1(14));
   U2900 : INV_X1 port map( A => io_out1_0_14_port, ZN => n2617);
   U2901 : AOI22_X1 port map( A1 => n3046, A2 => n2620, B1 => io_out1_1_14_port
                           , B2 => n3044, ZN => n2618);
   U2902 : AOI222_X1 port map( A1 => global_out1_14_port, A2 => n3071, B1 => 
                           io_out1_3_14_port, B2 => n3062, C1 => 
                           io_out1_2_14_port, C2 => n3052, ZN => n2619);
   U2903 : OAI211_X1 port map( C1 => n3070, C2 => n2609, A => n2610, B => n2611
                           , ZN => OUT1(15));
   U2904 : INV_X1 port map( A => io_out1_0_15_port, ZN => n2609);
   U2905 : AOI22_X1 port map( A1 => n3046, A2 => n2612, B1 => io_out1_1_15_port
                           , B2 => n3044, ZN => n2610);
   U2906 : AOI222_X1 port map( A1 => global_out1_15_port, A2 => n3073, B1 => 
                           io_out1_3_15_port, B2 => n3062, C1 => 
                           io_out1_2_15_port, C2 => n3052, ZN => n2611);
   U2907 : OAI211_X1 port map( C1 => n3070, C2 => n2601, A => n2602, B => n2603
                           , ZN => OUT1(16));
   U2908 : INV_X1 port map( A => io_out1_0_16_port, ZN => n2601);
   U2909 : AOI22_X1 port map( A1 => n3046, A2 => n2604, B1 => io_out1_1_16_port
                           , B2 => n3044, ZN => n2602);
   U2910 : AOI222_X1 port map( A1 => global_out1_16_port, A2 => n3071, B1 => 
                           io_out1_3_16_port, B2 => n3062, C1 => 
                           io_out1_2_16_port, C2 => n3052, ZN => n2603);
   U2911 : OAI211_X1 port map( C1 => n3070, C2 => n2593, A => n2594, B => n2595
                           , ZN => OUT1(17));
   U2912 : INV_X1 port map( A => io_out1_0_17_port, ZN => n2593);
   U2913 : AOI22_X1 port map( A1 => n3046, A2 => n2596, B1 => io_out1_1_17_port
                           , B2 => n3044, ZN => n2594);
   U2914 : AOI222_X1 port map( A1 => global_out1_17_port, A2 => n3073, B1 => 
                           io_out1_3_17_port, B2 => n3062, C1 => 
                           io_out1_2_17_port, C2 => n3052, ZN => n2595);
   U2915 : OAI211_X1 port map( C1 => n3070, C2 => n2585, A => n2586, B => n2587
                           , ZN => OUT1(18));
   U2916 : INV_X1 port map( A => io_out1_0_18_port, ZN => n2585);
   U2917 : AOI22_X1 port map( A1 => n3046, A2 => n2588, B1 => io_out1_1_18_port
                           , B2 => n3044, ZN => n2586);
   U2918 : AOI222_X1 port map( A1 => global_out1_18_port, A2 => n3073, B1 => 
                           io_out1_3_18_port, B2 => n3062, C1 => 
                           io_out1_2_18_port, C2 => n3052, ZN => n2587);
   U2919 : OAI211_X1 port map( C1 => n3070, C2 => n2577, A => n2578, B => n2579
                           , ZN => OUT1(19));
   U2920 : INV_X1 port map( A => io_out1_0_19_port, ZN => n2577);
   U2921 : AOI22_X1 port map( A1 => n3046, A2 => n2580, B1 => io_out1_1_19_port
                           , B2 => n3044, ZN => n2578);
   U2922 : AOI222_X1 port map( A1 => global_out1_19_port, A2 => n3071, B1 => 
                           io_out1_3_19_port, B2 => n3062, C1 => 
                           io_out1_2_19_port, C2 => n3052, ZN => n2579);
   U2923 : OAI211_X1 port map( C1 => n2138, C2 => n3066, A => n2140, B => n2141
                           , ZN => OUT1(9));
   U2924 : INV_X1 port map( A => io_out1_0_9_port, ZN => n2138);
   U2925 : AOI22_X1 port map( A1 => n3051, A2 => n2146, B1 => n3045, B2 => 
                           io_out1_1_9_port, ZN => n2140);
   U2926 : AOI222_X1 port map( A1 => global_out1_9_port, A2 => n3071, B1 => 
                           n3063, B2 => io_out1_3_9_port, C1 => n3057, C2 => 
                           io_out1_2_9_port, ZN => n2141);
   U2927 : INV_X1 port map( A => ADD_RD1(3), ZN => n2129);
   U2928 : AND3_X1 port map( A1 => ADD_WR(2), A2 => ADD_WR(3), A3 => WR, ZN => 
                           global_write);
   U2929 : INV_X1 port map( A => WR, ZN => n2114);
   U2930 : NOR2_X1 port map( A1 => RESET, A2 => n2105, ZN => n1035);
   U2931 : AOI22_X1 port map( A1 => n2106, A2 => n2107, B1 => CALL, B2 => n2108
                           , ZN => n2105);
   U2932 : INV_X1 port map( A => CALL, ZN => n2107);
   U2933 : OAI22_X1 port map( A1 => RETN, A2 => n2109, B1 => n2110, B2 => n2111
                           , ZN => n2106);
   U2934 : NOR2_X1 port map( A1 => RESET, A2 => n2102, ZN => n1036);
   U2935 : XNOR2_X1 port map( A => n2103, B => n2104, ZN => n2102);
   U2936 : NOR2_X1 port map( A1 => CALL, A2 => RETN, ZN => n2104);
   U2937 : INV_X1 port map( A => RD2, ZN => n2117);
   U2938 : INV_X1 port map( A => ADD_RD2(3), ZN => n2123);
   U2939 : INV_X1 port map( A => RETN, ZN => n2111);
   U2940 : OAI21_X1 port map( B1 => n2932, B2 => n2131, A => n2936, ZN => n2678
                           );
   U2941 : AOI22_X1 port map( A1 => loc_out2_2_36_port, A2 => n2983, B1 => 
                           io_out2_1_36_port, B2 => n2977, ZN => n2787);
   U2942 : AOI22_X1 port map( A1 => loc_out2_2_37_port, A2 => n2983, B1 => 
                           io_out2_1_37_port, B2 => n2977, ZN => n2783);
   U2943 : AOI22_X1 port map( A1 => loc_out2_2_38_port, A2 => n2983, B1 => 
                           io_out2_1_38_port, B2 => n2977, ZN => n2779);
   U2944 : AOI22_X1 port map( A1 => loc_out2_2_39_port, A2 => n2983, B1 => 
                           io_out2_1_39_port, B2 => n2977, ZN => n2775);
   U2945 : AOI22_X1 port map( A1 => loc_out2_2_40_port, A2 => n2983, B1 => 
                           io_out2_1_40_port, B2 => n2977, ZN => n2771);
   U2946 : AOI22_X1 port map( A1 => loc_out2_2_41_port, A2 => n2983, B1 => 
                           io_out2_1_41_port, B2 => n2977, ZN => n2767);
   U2947 : AOI22_X1 port map( A1 => loc_out2_2_42_port, A2 => n2983, B1 => 
                           io_out2_1_42_port, B2 => n2977, ZN => n2763);
   U2948 : AOI22_X1 port map( A1 => loc_out2_2_43_port, A2 => n2983, B1 => 
                           io_out2_1_43_port, B2 => n2977, ZN => n2759);
   U2949 : AOI22_X1 port map( A1 => loc_out2_2_44_port, A2 => n2983, B1 => 
                           io_out2_1_44_port, B2 => n2977, ZN => n2755);
   U2950 : AOI22_X1 port map( A1 => loc_out2_2_45_port, A2 => n2983, B1 => 
                           io_out2_1_45_port, B2 => n2977, ZN => n2751);
   U2951 : AOI22_X1 port map( A1 => loc_out2_2_46_port, A2 => n2983, B1 => 
                           io_out2_1_46_port, B2 => n2977, ZN => n2747);
   U2952 : AOI22_X1 port map( A1 => loc_out2_2_47_port, A2 => n2983, B1 => 
                           io_out2_1_47_port, B2 => n2977, ZN => n2743);
   U2953 : AOI22_X1 port map( A1 => loc_out2_2_48_port, A2 => n2984, B1 => 
                           io_out2_1_48_port, B2 => n2978, ZN => n2739);
   U2954 : AOI22_X1 port map( A1 => loc_out2_2_49_port, A2 => n2984, B1 => 
                           io_out2_1_49_port, B2 => n2978, ZN => n2735);
   U2955 : AOI22_X1 port map( A1 => loc_out2_2_50_port, A2 => n2984, B1 => 
                           io_out2_1_50_port, B2 => n2978, ZN => n2731);
   U2956 : AOI22_X1 port map( A1 => loc_out2_2_51_port, A2 => n2984, B1 => 
                           io_out2_1_51_port, B2 => n2978, ZN => n2727);
   U2957 : AOI22_X1 port map( A1 => loc_out2_2_52_port, A2 => n2984, B1 => 
                           io_out2_1_52_port, B2 => n2978, ZN => n2723);
   U2958 : AOI22_X1 port map( A1 => loc_out2_2_53_port, A2 => n2984, B1 => 
                           io_out2_1_53_port, B2 => n2978, ZN => n2719);
   U2959 : AOI22_X1 port map( A1 => loc_out2_2_54_port, A2 => n2984, B1 => 
                           io_out2_1_54_port, B2 => n2978, ZN => n2715);
   U2960 : AOI22_X1 port map( A1 => loc_out2_2_55_port, A2 => n2984, B1 => 
                           io_out2_1_55_port, B2 => n2978, ZN => n2711);
   U2961 : AOI22_X1 port map( A1 => loc_out2_2_56_port, A2 => n2984, B1 => 
                           io_out2_1_56_port, B2 => n2978, ZN => n2707);
   U2962 : AOI22_X1 port map( A1 => loc_out2_2_57_port, A2 => n2984, B1 => 
                           io_out2_1_57_port, B2 => n2978, ZN => n2703);
   U2963 : AOI22_X1 port map( A1 => loc_out2_2_58_port, A2 => n2984, B1 => 
                           io_out2_1_58_port, B2 => n2978, ZN => n2699);
   U2964 : AOI22_X1 port map( A1 => loc_out2_2_59_port, A2 => n2984, B1 => 
                           io_out2_1_59_port, B2 => n2978, ZN => n2695);
   U2965 : AOI22_X1 port map( A1 => loc_out2_2_60_port, A2 => n2985, B1 => 
                           io_out2_1_60_port, B2 => n2979, ZN => n2691);
   U2966 : AOI22_X1 port map( A1 => loc_out2_2_61_port, A2 => n2985, B1 => 
                           io_out2_1_61_port, B2 => n2979, ZN => n2687);
   U2967 : AOI22_X1 port map( A1 => loc_out2_2_62_port, A2 => n2985, B1 => 
                           io_out2_1_62_port, B2 => n2979, ZN => n2683);
   U2968 : AOI22_X1 port map( A1 => loc_out2_2_63_port, A2 => n2985, B1 => 
                           io_out2_1_63_port, B2 => n2979, ZN => n2671);
   U2969 : AOI22_X1 port map( A1 => loc_out2_2_0_port, A2 => n2980, B1 => 
                           io_out2_1_0_port, B2 => n2974, ZN => n2931);
   U2970 : AOI22_X1 port map( A1 => loc_out2_2_1_port, A2 => n2980, B1 => 
                           io_out2_1_1_port, B2 => n2974, ZN => n2927);
   U2971 : AOI22_X1 port map( A1 => loc_out2_2_2_port, A2 => n2980, B1 => 
                           io_out2_1_2_port, B2 => n2974, ZN => n2923);
   U2972 : AOI22_X1 port map( A1 => loc_out2_2_3_port, A2 => n2980, B1 => 
                           io_out2_1_3_port, B2 => n2974, ZN => n2919);
   U2973 : AOI22_X1 port map( A1 => loc_out2_2_4_port, A2 => n2980, B1 => 
                           io_out2_1_4_port, B2 => n2974, ZN => n2915);
   U2974 : AOI22_X1 port map( A1 => loc_out2_2_5_port, A2 => n2980, B1 => 
                           io_out2_1_5_port, B2 => n2974, ZN => n2911);
   U2975 : AOI22_X1 port map( A1 => loc_out2_2_6_port, A2 => n2980, B1 => 
                           io_out2_1_6_port, B2 => n2974, ZN => n2907);
   U2976 : AOI22_X1 port map( A1 => loc_out2_2_7_port, A2 => n2980, B1 => 
                           io_out2_1_7_port, B2 => n2974, ZN => n2903);
   U2977 : AOI22_X1 port map( A1 => loc_out2_2_8_port, A2 => n2980, B1 => 
                           io_out2_1_8_port, B2 => n2974, ZN => n2899);
   U2978 : AOI22_X1 port map( A1 => loc_out2_2_9_port, A2 => n2980, B1 => 
                           io_out2_1_9_port, B2 => n2974, ZN => n2895);
   U2979 : AOI22_X1 port map( A1 => loc_out2_2_10_port, A2 => n2980, B1 => 
                           io_out2_1_10_port, B2 => n2974, ZN => n2891);
   U2980 : AOI22_X1 port map( A1 => loc_out2_2_11_port, A2 => n2980, B1 => 
                           io_out2_1_11_port, B2 => n2974, ZN => n2887);
   U2981 : AOI22_X1 port map( A1 => loc_out2_2_12_port, A2 => n2981, B1 => 
                           io_out2_1_12_port, B2 => n2975, ZN => n2883);
   U2982 : AOI22_X1 port map( A1 => loc_out2_2_13_port, A2 => n2981, B1 => 
                           io_out2_1_13_port, B2 => n2975, ZN => n2879);
   U2983 : AOI22_X1 port map( A1 => loc_out2_2_14_port, A2 => n2981, B1 => 
                           io_out2_1_14_port, B2 => n2975, ZN => n2875);
   U2984 : AOI22_X1 port map( A1 => loc_out2_2_15_port, A2 => n2981, B1 => 
                           io_out2_1_15_port, B2 => n2975, ZN => n2871);
   U2985 : AOI22_X1 port map( A1 => loc_out2_2_16_port, A2 => n2981, B1 => 
                           io_out2_1_16_port, B2 => n2975, ZN => n2867);
   U2986 : AOI22_X1 port map( A1 => loc_out2_2_17_port, A2 => n2981, B1 => 
                           io_out2_1_17_port, B2 => n2975, ZN => n2863);
   U2987 : AOI22_X1 port map( A1 => loc_out2_2_18_port, A2 => n2981, B1 => 
                           io_out2_1_18_port, B2 => n2975, ZN => n2859);
   U2988 : AOI22_X1 port map( A1 => loc_out2_2_19_port, A2 => n2981, B1 => 
                           io_out2_1_19_port, B2 => n2975, ZN => n2855);
   U2989 : AOI22_X1 port map( A1 => loc_out2_2_20_port, A2 => n2981, B1 => 
                           io_out2_1_20_port, B2 => n2975, ZN => n2851);
   U2990 : AOI22_X1 port map( A1 => loc_out2_2_21_port, A2 => n2981, B1 => 
                           io_out2_1_21_port, B2 => n2975, ZN => n2847);
   U2991 : AOI22_X1 port map( A1 => loc_out2_2_22_port, A2 => n2981, B1 => 
                           io_out2_1_22_port, B2 => n2975, ZN => n2843);
   U2992 : AOI22_X1 port map( A1 => loc_out2_2_23_port, A2 => n2981, B1 => 
                           io_out2_1_23_port, B2 => n2975, ZN => n2839);
   U2993 : AOI22_X1 port map( A1 => loc_out2_2_24_port, A2 => n2982, B1 => 
                           io_out2_1_24_port, B2 => n2976, ZN => n2835);
   U2994 : AOI22_X1 port map( A1 => loc_out2_2_25_port, A2 => n2982, B1 => 
                           io_out2_1_25_port, B2 => n2976, ZN => n2831);
   U2995 : AOI22_X1 port map( A1 => loc_out2_2_26_port, A2 => n2982, B1 => 
                           io_out2_1_26_port, B2 => n2976, ZN => n2827);
   U2996 : AOI22_X1 port map( A1 => loc_out2_2_27_port, A2 => n2982, B1 => 
                           io_out2_1_27_port, B2 => n2976, ZN => n2823);
   U2997 : AOI22_X1 port map( A1 => loc_out2_2_28_port, A2 => n2982, B1 => 
                           io_out2_1_28_port, B2 => n2976, ZN => n2819);
   U2998 : AOI22_X1 port map( A1 => loc_out2_2_29_port, A2 => n2982, B1 => 
                           io_out2_1_29_port, B2 => n2976, ZN => n2815);
   U2999 : AOI22_X1 port map( A1 => loc_out2_2_30_port, A2 => n2982, B1 => 
                           io_out2_1_30_port, B2 => n2976, ZN => n2811);
   U3000 : AOI22_X1 port map( A1 => loc_out2_2_31_port, A2 => n2982, B1 => 
                           io_out2_1_31_port, B2 => n2976, ZN => n2807);
   U3001 : AOI22_X1 port map( A1 => loc_out2_2_32_port, A2 => n2982, B1 => 
                           io_out2_1_32_port, B2 => n2976, ZN => n2803);
   U3002 : AOI22_X1 port map( A1 => loc_out2_2_33_port, A2 => n2982, B1 => 
                           io_out2_1_33_port, B2 => n2976, ZN => n2799);
   U3003 : AOI22_X1 port map( A1 => loc_out2_2_34_port, A2 => n2982, B1 => 
                           io_out2_1_34_port, B2 => n2976, ZN => n2795);
   U3004 : AOI22_X1 port map( A1 => loc_out2_2_35_port, A2 => n2982, B1 => 
                           io_out2_1_35_port, B2 => n2976, ZN => n2791);
   U3005 : NAND4_X1 port map( A1 => n2688, A2 => n2689, A3 => n2690, A4 => 
                           n2691, ZN => N1192);
   U3006 : AOI22_X1 port map( A1 => io_out2_2_60_port, A2 => n2949, B1 => 
                           io_out2_3_60_port, B2 => n2943, ZN => n2688);
   U3007 : AOI22_X1 port map( A1 => loc_out2_0_60_port, A2 => n2961, B1 => 
                           io_out2_0_60_port, B2 => n2955, ZN => n2689);
   U3008 : AOI22_X1 port map( A1 => loc_out2_1_60_port, A2 => n2973, B1 => 
                           loc_out2_3_60_port, B2 => n2967, ZN => n2690);
   U3009 : NAND4_X1 port map( A1 => n2684, A2 => n2685, A3 => n2686, A4 => 
                           n2687, ZN => N1193);
   U3010 : AOI22_X1 port map( A1 => io_out2_2_61_port, A2 => n2949, B1 => 
                           io_out2_3_61_port, B2 => n2943, ZN => n2684);
   U3011 : AOI22_X1 port map( A1 => loc_out2_0_61_port, A2 => n2961, B1 => 
                           io_out2_0_61_port, B2 => n2955, ZN => n2685);
   U3012 : AOI22_X1 port map( A1 => loc_out2_1_61_port, A2 => n2973, B1 => 
                           loc_out2_3_61_port, B2 => n2967, ZN => n2686);
   U3013 : NAND4_X1 port map( A1 => n2680, A2 => n2681, A3 => n2682, A4 => 
                           n2683, ZN => N1194);
   U3014 : AOI22_X1 port map( A1 => io_out2_2_62_port, A2 => n2949, B1 => 
                           io_out2_3_62_port, B2 => n2943, ZN => n2680);
   U3015 : AOI22_X1 port map( A1 => loc_out2_0_62_port, A2 => n2961, B1 => 
                           io_out2_0_62_port, B2 => n2955, ZN => n2681);
   U3016 : AOI22_X1 port map( A1 => loc_out2_1_62_port, A2 => n2973, B1 => 
                           loc_out2_3_62_port, B2 => n2967, ZN => n2682);
   U3017 : NAND4_X1 port map( A1 => n2668, A2 => n2669, A3 => n2670, A4 => 
                           n2671, ZN => N1195);
   U3018 : AOI22_X1 port map( A1 => io_out2_2_63_port, A2 => n2949, B1 => 
                           io_out2_3_63_port, B2 => n2943, ZN => n2668);
   U3019 : AOI22_X1 port map( A1 => loc_out2_0_63_port, A2 => n2961, B1 => 
                           io_out2_0_63_port, B2 => n2955, ZN => n2669);
   U3020 : AOI22_X1 port map( A1 => loc_out2_1_63_port, A2 => n2973, B1 => 
                           loc_out2_3_63_port, B2 => n2967, ZN => n2670);
   U3021 : NAND4_X1 port map( A1 => n2928, A2 => n2929, A3 => n2930, A4 => 
                           n2931, ZN => N1132);
   U3022 : AOI22_X1 port map( A1 => io_out2_2_0_port, A2 => n2944, B1 => 
                           io_out2_3_0_port, B2 => n2938, ZN => n2928);
   U3023 : AOI22_X1 port map( A1 => loc_out2_0_0_port, A2 => n2956, B1 => 
                           io_out2_0_0_port, B2 => n2950, ZN => n2929);
   U3024 : AOI22_X1 port map( A1 => loc_out2_1_0_port, A2 => n2968, B1 => 
                           loc_out2_3_0_port, B2 => n2962, ZN => n2930);
   U3025 : NAND4_X1 port map( A1 => n2924, A2 => n2925, A3 => n2926, A4 => 
                           n2927, ZN => N1133);
   U3026 : AOI22_X1 port map( A1 => io_out2_2_1_port, A2 => n2944, B1 => 
                           io_out2_3_1_port, B2 => n2938, ZN => n2924);
   U3027 : AOI22_X1 port map( A1 => loc_out2_0_1_port, A2 => n2956, B1 => 
                           io_out2_0_1_port, B2 => n2950, ZN => n2925);
   U3028 : AOI22_X1 port map( A1 => loc_out2_1_1_port, A2 => n2968, B1 => 
                           loc_out2_3_1_port, B2 => n2962, ZN => n2926);
   U3029 : NAND4_X1 port map( A1 => n2920, A2 => n2921, A3 => n2922, A4 => 
                           n2923, ZN => N1134);
   U3030 : AOI22_X1 port map( A1 => io_out2_2_2_port, A2 => n2944, B1 => 
                           io_out2_3_2_port, B2 => n2938, ZN => n2920);
   U3031 : AOI22_X1 port map( A1 => loc_out2_0_2_port, A2 => n2956, B1 => 
                           io_out2_0_2_port, B2 => n2950, ZN => n2921);
   U3032 : AOI22_X1 port map( A1 => loc_out2_1_2_port, A2 => n2968, B1 => 
                           loc_out2_3_2_port, B2 => n2962, ZN => n2922);
   U3033 : NAND4_X1 port map( A1 => n2916, A2 => n2917, A3 => n2918, A4 => 
                           n2919, ZN => N1135);
   U3034 : AOI22_X1 port map( A1 => io_out2_2_3_port, A2 => n2944, B1 => 
                           io_out2_3_3_port, B2 => n2938, ZN => n2916);
   U3035 : AOI22_X1 port map( A1 => loc_out2_0_3_port, A2 => n2956, B1 => 
                           io_out2_0_3_port, B2 => n2950, ZN => n2917);
   U3036 : AOI22_X1 port map( A1 => loc_out2_1_3_port, A2 => n2968, B1 => 
                           loc_out2_3_3_port, B2 => n2962, ZN => n2918);
   U3037 : NAND4_X1 port map( A1 => n2912, A2 => n2913, A3 => n2914, A4 => 
                           n2915, ZN => N1136);
   U3038 : AOI22_X1 port map( A1 => io_out2_2_4_port, A2 => n2944, B1 => 
                           io_out2_3_4_port, B2 => n2938, ZN => n2912);
   U3039 : AOI22_X1 port map( A1 => loc_out2_0_4_port, A2 => n2956, B1 => 
                           io_out2_0_4_port, B2 => n2950, ZN => n2913);
   U3040 : AOI22_X1 port map( A1 => loc_out2_1_4_port, A2 => n2968, B1 => 
                           loc_out2_3_4_port, B2 => n2962, ZN => n2914);
   U3041 : NAND4_X1 port map( A1 => n2908, A2 => n2909, A3 => n2910, A4 => 
                           n2911, ZN => N1137);
   U3042 : AOI22_X1 port map( A1 => io_out2_2_5_port, A2 => n2944, B1 => 
                           io_out2_3_5_port, B2 => n2938, ZN => n2908);
   U3043 : AOI22_X1 port map( A1 => loc_out2_0_5_port, A2 => n2956, B1 => 
                           io_out2_0_5_port, B2 => n2950, ZN => n2909);
   U3044 : AOI22_X1 port map( A1 => loc_out2_1_5_port, A2 => n2968, B1 => 
                           loc_out2_3_5_port, B2 => n2962, ZN => n2910);
   U3045 : NAND4_X1 port map( A1 => n2904, A2 => n2905, A3 => n2906, A4 => 
                           n2907, ZN => N1138);
   U3046 : AOI22_X1 port map( A1 => io_out2_2_6_port, A2 => n2944, B1 => 
                           io_out2_3_6_port, B2 => n2938, ZN => n2904);
   U3047 : AOI22_X1 port map( A1 => loc_out2_0_6_port, A2 => n2956, B1 => 
                           io_out2_0_6_port, B2 => n2950, ZN => n2905);
   U3048 : AOI22_X1 port map( A1 => loc_out2_1_6_port, A2 => n2968, B1 => 
                           loc_out2_3_6_port, B2 => n2962, ZN => n2906);
   U3049 : NAND4_X1 port map( A1 => n2900, A2 => n2901, A3 => n2902, A4 => 
                           n2903, ZN => N1139);
   U3050 : AOI22_X1 port map( A1 => io_out2_2_7_port, A2 => n2944, B1 => 
                           io_out2_3_7_port, B2 => n2938, ZN => n2900);
   U3051 : AOI22_X1 port map( A1 => loc_out2_0_7_port, A2 => n2956, B1 => 
                           io_out2_0_7_port, B2 => n2950, ZN => n2901);
   U3052 : AOI22_X1 port map( A1 => loc_out2_1_7_port, A2 => n2968, B1 => 
                           loc_out2_3_7_port, B2 => n2962, ZN => n2902);
   U3053 : NAND4_X1 port map( A1 => n2896, A2 => n2897, A3 => n2898, A4 => 
                           n2899, ZN => N1140);
   U3054 : AOI22_X1 port map( A1 => io_out2_2_8_port, A2 => n2944, B1 => 
                           io_out2_3_8_port, B2 => n2938, ZN => n2896);
   U3055 : AOI22_X1 port map( A1 => loc_out2_0_8_port, A2 => n2956, B1 => 
                           io_out2_0_8_port, B2 => n2950, ZN => n2897);
   U3056 : AOI22_X1 port map( A1 => loc_out2_1_8_port, A2 => n2968, B1 => 
                           loc_out2_3_8_port, B2 => n2962, ZN => n2898);
   U3057 : NAND4_X1 port map( A1 => n2892, A2 => n2893, A3 => n2894, A4 => 
                           n2895, ZN => N1141);
   U3058 : AOI22_X1 port map( A1 => io_out2_2_9_port, A2 => n2944, B1 => 
                           io_out2_3_9_port, B2 => n2938, ZN => n2892);
   U3059 : AOI22_X1 port map( A1 => loc_out2_0_9_port, A2 => n2956, B1 => 
                           io_out2_0_9_port, B2 => n2950, ZN => n2893);
   U3060 : AOI22_X1 port map( A1 => loc_out2_1_9_port, A2 => n2968, B1 => 
                           loc_out2_3_9_port, B2 => n2962, ZN => n2894);
   U3061 : NAND4_X1 port map( A1 => n2888, A2 => n2889, A3 => n2890, A4 => 
                           n2891, ZN => N1142);
   U3062 : AOI22_X1 port map( A1 => io_out2_2_10_port, A2 => n2944, B1 => 
                           io_out2_3_10_port, B2 => n2938, ZN => n2888);
   U3063 : AOI22_X1 port map( A1 => loc_out2_0_10_port, A2 => n2956, B1 => 
                           io_out2_0_10_port, B2 => n2950, ZN => n2889);
   U3064 : AOI22_X1 port map( A1 => loc_out2_1_10_port, A2 => n2968, B1 => 
                           loc_out2_3_10_port, B2 => n2962, ZN => n2890);
   U3065 : NAND4_X1 port map( A1 => n2884, A2 => n2885, A3 => n2886, A4 => 
                           n2887, ZN => N1143);
   U3066 : AOI22_X1 port map( A1 => io_out2_2_11_port, A2 => n2944, B1 => 
                           io_out2_3_11_port, B2 => n2938, ZN => n2884);
   U3067 : AOI22_X1 port map( A1 => loc_out2_0_11_port, A2 => n2956, B1 => 
                           io_out2_0_11_port, B2 => n2950, ZN => n2885);
   U3068 : AOI22_X1 port map( A1 => loc_out2_1_11_port, A2 => n2968, B1 => 
                           loc_out2_3_11_port, B2 => n2962, ZN => n2886);
   U3069 : NAND4_X1 port map( A1 => n2880, A2 => n2881, A3 => n2882, A4 => 
                           n2883, ZN => N1144);
   U3070 : AOI22_X1 port map( A1 => io_out2_2_12_port, A2 => n2945, B1 => 
                           io_out2_3_12_port, B2 => n2939, ZN => n2880);
   U3071 : AOI22_X1 port map( A1 => loc_out2_0_12_port, A2 => n2957, B1 => 
                           io_out2_0_12_port, B2 => n2951, ZN => n2881);
   U3072 : AOI22_X1 port map( A1 => loc_out2_1_12_port, A2 => n2969, B1 => 
                           loc_out2_3_12_port, B2 => n2963, ZN => n2882);
   U3073 : NAND4_X1 port map( A1 => n2876, A2 => n2877, A3 => n2878, A4 => 
                           n2879, ZN => N1145);
   U3074 : AOI22_X1 port map( A1 => io_out2_2_13_port, A2 => n2945, B1 => 
                           io_out2_3_13_port, B2 => n2939, ZN => n2876);
   U3075 : AOI22_X1 port map( A1 => loc_out2_0_13_port, A2 => n2957, B1 => 
                           io_out2_0_13_port, B2 => n2951, ZN => n2877);
   U3076 : AOI22_X1 port map( A1 => loc_out2_1_13_port, A2 => n2969, B1 => 
                           loc_out2_3_13_port, B2 => n2963, ZN => n2878);
   U3077 : NAND4_X1 port map( A1 => n2872, A2 => n2873, A3 => n2874, A4 => 
                           n2875, ZN => N1146);
   U3078 : AOI22_X1 port map( A1 => io_out2_2_14_port, A2 => n2945, B1 => 
                           io_out2_3_14_port, B2 => n2939, ZN => n2872);
   U3079 : AOI22_X1 port map( A1 => loc_out2_0_14_port, A2 => n2957, B1 => 
                           io_out2_0_14_port, B2 => n2951, ZN => n2873);
   U3080 : AOI22_X1 port map( A1 => loc_out2_1_14_port, A2 => n2969, B1 => 
                           loc_out2_3_14_port, B2 => n2963, ZN => n2874);
   U3081 : NAND4_X1 port map( A1 => n2868, A2 => n2869, A3 => n2870, A4 => 
                           n2871, ZN => N1147);
   U3082 : AOI22_X1 port map( A1 => io_out2_2_15_port, A2 => n2945, B1 => 
                           io_out2_3_15_port, B2 => n2939, ZN => n2868);
   U3083 : AOI22_X1 port map( A1 => loc_out2_0_15_port, A2 => n2957, B1 => 
                           io_out2_0_15_port, B2 => n2951, ZN => n2869);
   U3084 : AOI22_X1 port map( A1 => loc_out2_1_15_port, A2 => n2969, B1 => 
                           loc_out2_3_15_port, B2 => n2963, ZN => n2870);
   U3085 : NAND4_X1 port map( A1 => n2864, A2 => n2865, A3 => n2866, A4 => 
                           n2867, ZN => N1148);
   U3086 : AOI22_X1 port map( A1 => io_out2_2_16_port, A2 => n2945, B1 => 
                           io_out2_3_16_port, B2 => n2939, ZN => n2864);
   U3087 : AOI22_X1 port map( A1 => loc_out2_0_16_port, A2 => n2957, B1 => 
                           io_out2_0_16_port, B2 => n2951, ZN => n2865);
   U3088 : AOI22_X1 port map( A1 => loc_out2_1_16_port, A2 => n2969, B1 => 
                           loc_out2_3_16_port, B2 => n2963, ZN => n2866);
   U3089 : NAND4_X1 port map( A1 => n2860, A2 => n2861, A3 => n2862, A4 => 
                           n2863, ZN => N1149);
   U3090 : AOI22_X1 port map( A1 => io_out2_2_17_port, A2 => n2945, B1 => 
                           io_out2_3_17_port, B2 => n2939, ZN => n2860);
   U3091 : AOI22_X1 port map( A1 => loc_out2_0_17_port, A2 => n2957, B1 => 
                           io_out2_0_17_port, B2 => n2951, ZN => n2861);
   U3092 : AOI22_X1 port map( A1 => loc_out2_1_17_port, A2 => n2969, B1 => 
                           loc_out2_3_17_port, B2 => n2963, ZN => n2862);
   U3093 : NAND4_X1 port map( A1 => n2856, A2 => n2857, A3 => n2858, A4 => 
                           n2859, ZN => N1150);
   U3094 : AOI22_X1 port map( A1 => io_out2_2_18_port, A2 => n2945, B1 => 
                           io_out2_3_18_port, B2 => n2939, ZN => n2856);
   U3095 : AOI22_X1 port map( A1 => loc_out2_0_18_port, A2 => n2957, B1 => 
                           io_out2_0_18_port, B2 => n2951, ZN => n2857);
   U3096 : AOI22_X1 port map( A1 => loc_out2_1_18_port, A2 => n2969, B1 => 
                           loc_out2_3_18_port, B2 => n2963, ZN => n2858);
   U3097 : NAND4_X1 port map( A1 => n2852, A2 => n2853, A3 => n2854, A4 => 
                           n2855, ZN => N1151);
   U3098 : AOI22_X1 port map( A1 => io_out2_2_19_port, A2 => n2945, B1 => 
                           io_out2_3_19_port, B2 => n2939, ZN => n2852);
   U3099 : AOI22_X1 port map( A1 => loc_out2_0_19_port, A2 => n2957, B1 => 
                           io_out2_0_19_port, B2 => n2951, ZN => n2853);
   U3100 : AOI22_X1 port map( A1 => loc_out2_1_19_port, A2 => n2969, B1 => 
                           loc_out2_3_19_port, B2 => n2963, ZN => n2854);
   U3101 : NAND4_X1 port map( A1 => n2848, A2 => n2849, A3 => n2850, A4 => 
                           n2851, ZN => N1152);
   U3102 : AOI22_X1 port map( A1 => io_out2_2_20_port, A2 => n2945, B1 => 
                           io_out2_3_20_port, B2 => n2939, ZN => n2848);
   U3103 : AOI22_X1 port map( A1 => loc_out2_0_20_port, A2 => n2957, B1 => 
                           io_out2_0_20_port, B2 => n2951, ZN => n2849);
   U3104 : AOI22_X1 port map( A1 => loc_out2_1_20_port, A2 => n2969, B1 => 
                           loc_out2_3_20_port, B2 => n2963, ZN => n2850);
   U3105 : NAND4_X1 port map( A1 => n2844, A2 => n2845, A3 => n2846, A4 => 
                           n2847, ZN => N1153);
   U3106 : AOI22_X1 port map( A1 => io_out2_2_21_port, A2 => n2945, B1 => 
                           io_out2_3_21_port, B2 => n2939, ZN => n2844);
   U3107 : AOI22_X1 port map( A1 => loc_out2_0_21_port, A2 => n2957, B1 => 
                           io_out2_0_21_port, B2 => n2951, ZN => n2845);
   U3108 : AOI22_X1 port map( A1 => loc_out2_1_21_port, A2 => n2969, B1 => 
                           loc_out2_3_21_port, B2 => n2963, ZN => n2846);
   U3109 : NAND4_X1 port map( A1 => n2840, A2 => n2841, A3 => n2842, A4 => 
                           n2843, ZN => N1154);
   U3110 : AOI22_X1 port map( A1 => io_out2_2_22_port, A2 => n2945, B1 => 
                           io_out2_3_22_port, B2 => n2939, ZN => n2840);
   U3111 : AOI22_X1 port map( A1 => loc_out2_0_22_port, A2 => n2957, B1 => 
                           io_out2_0_22_port, B2 => n2951, ZN => n2841);
   U3112 : AOI22_X1 port map( A1 => loc_out2_1_22_port, A2 => n2969, B1 => 
                           loc_out2_3_22_port, B2 => n2963, ZN => n2842);
   U3113 : NAND4_X1 port map( A1 => n2836, A2 => n2837, A3 => n2838, A4 => 
                           n2839, ZN => N1155);
   U3114 : AOI22_X1 port map( A1 => io_out2_2_23_port, A2 => n2945, B1 => 
                           io_out2_3_23_port, B2 => n2939, ZN => n2836);
   U3115 : AOI22_X1 port map( A1 => loc_out2_0_23_port, A2 => n2957, B1 => 
                           io_out2_0_23_port, B2 => n2951, ZN => n2837);
   U3116 : AOI22_X1 port map( A1 => loc_out2_1_23_port, A2 => n2969, B1 => 
                           loc_out2_3_23_port, B2 => n2963, ZN => n2838);
   U3117 : NAND4_X1 port map( A1 => n2832, A2 => n2833, A3 => n2834, A4 => 
                           n2835, ZN => N1156);
   U3118 : AOI22_X1 port map( A1 => io_out2_2_24_port, A2 => n2946, B1 => 
                           io_out2_3_24_port, B2 => n2940, ZN => n2832);
   U3119 : AOI22_X1 port map( A1 => loc_out2_0_24_port, A2 => n2958, B1 => 
                           io_out2_0_24_port, B2 => n2952, ZN => n2833);
   U3120 : AOI22_X1 port map( A1 => loc_out2_1_24_port, A2 => n2970, B1 => 
                           loc_out2_3_24_port, B2 => n2964, ZN => n2834);
   U3121 : NAND4_X1 port map( A1 => n2828, A2 => n2829, A3 => n2830, A4 => 
                           n2831, ZN => N1157);
   U3122 : AOI22_X1 port map( A1 => io_out2_2_25_port, A2 => n2946, B1 => 
                           io_out2_3_25_port, B2 => n2940, ZN => n2828);
   U3123 : AOI22_X1 port map( A1 => loc_out2_0_25_port, A2 => n2958, B1 => 
                           io_out2_0_25_port, B2 => n2952, ZN => n2829);
   U3124 : AOI22_X1 port map( A1 => loc_out2_1_25_port, A2 => n2970, B1 => 
                           loc_out2_3_25_port, B2 => n2964, ZN => n2830);
   U3125 : NAND4_X1 port map( A1 => n2824, A2 => n2825, A3 => n2826, A4 => 
                           n2827, ZN => N1158);
   U3126 : AOI22_X1 port map( A1 => io_out2_2_26_port, A2 => n2946, B1 => 
                           io_out2_3_26_port, B2 => n2940, ZN => n2824);
   U3127 : AOI22_X1 port map( A1 => loc_out2_0_26_port, A2 => n2958, B1 => 
                           io_out2_0_26_port, B2 => n2952, ZN => n2825);
   U3128 : AOI22_X1 port map( A1 => loc_out2_1_26_port, A2 => n2970, B1 => 
                           loc_out2_3_26_port, B2 => n2964, ZN => n2826);
   U3129 : NAND4_X1 port map( A1 => n2820, A2 => n2821, A3 => n2822, A4 => 
                           n2823, ZN => N1159);
   U3130 : AOI22_X1 port map( A1 => io_out2_2_27_port, A2 => n2946, B1 => 
                           io_out2_3_27_port, B2 => n2940, ZN => n2820);
   U3131 : AOI22_X1 port map( A1 => loc_out2_0_27_port, A2 => n2958, B1 => 
                           io_out2_0_27_port, B2 => n2952, ZN => n2821);
   U3132 : AOI22_X1 port map( A1 => loc_out2_1_27_port, A2 => n2970, B1 => 
                           loc_out2_3_27_port, B2 => n2964, ZN => n2822);
   U3133 : NAND4_X1 port map( A1 => n2816, A2 => n2817, A3 => n2818, A4 => 
                           n2819, ZN => N1160);
   U3134 : AOI22_X1 port map( A1 => io_out2_2_28_port, A2 => n2946, B1 => 
                           io_out2_3_28_port, B2 => n2940, ZN => n2816);
   U3135 : AOI22_X1 port map( A1 => loc_out2_0_28_port, A2 => n2958, B1 => 
                           io_out2_0_28_port, B2 => n2952, ZN => n2817);
   U3136 : AOI22_X1 port map( A1 => loc_out2_1_28_port, A2 => n2970, B1 => 
                           loc_out2_3_28_port, B2 => n2964, ZN => n2818);
   U3137 : NAND4_X1 port map( A1 => n2812, A2 => n2813, A3 => n2814, A4 => 
                           n2815, ZN => N1161);
   U3138 : AOI22_X1 port map( A1 => io_out2_2_29_port, A2 => n2946, B1 => 
                           io_out2_3_29_port, B2 => n2940, ZN => n2812);
   U3139 : AOI22_X1 port map( A1 => loc_out2_0_29_port, A2 => n2958, B1 => 
                           io_out2_0_29_port, B2 => n2952, ZN => n2813);
   U3140 : AOI22_X1 port map( A1 => loc_out2_1_29_port, A2 => n2970, B1 => 
                           loc_out2_3_29_port, B2 => n2964, ZN => n2814);
   U3141 : NAND4_X1 port map( A1 => n2808, A2 => n2809, A3 => n2810, A4 => 
                           n2811, ZN => N1162);
   U3142 : AOI22_X1 port map( A1 => io_out2_2_30_port, A2 => n2946, B1 => 
                           io_out2_3_30_port, B2 => n2940, ZN => n2808);
   U3143 : AOI22_X1 port map( A1 => loc_out2_0_30_port, A2 => n2958, B1 => 
                           io_out2_0_30_port, B2 => n2952, ZN => n2809);
   U3144 : AOI22_X1 port map( A1 => loc_out2_1_30_port, A2 => n2970, B1 => 
                           loc_out2_3_30_port, B2 => n2964, ZN => n2810);
   U3145 : NAND4_X1 port map( A1 => n2804, A2 => n2805, A3 => n2806, A4 => 
                           n2807, ZN => N1163);
   U3146 : AOI22_X1 port map( A1 => io_out2_2_31_port, A2 => n2946, B1 => 
                           io_out2_3_31_port, B2 => n2940, ZN => n2804);
   U3147 : AOI22_X1 port map( A1 => loc_out2_0_31_port, A2 => n2958, B1 => 
                           io_out2_0_31_port, B2 => n2952, ZN => n2805);
   U3148 : AOI22_X1 port map( A1 => loc_out2_1_31_port, A2 => n2970, B1 => 
                           loc_out2_3_31_port, B2 => n2964, ZN => n2806);
   U3149 : NAND4_X1 port map( A1 => n2800, A2 => n2801, A3 => n2802, A4 => 
                           n2803, ZN => N1164);
   U3150 : AOI22_X1 port map( A1 => io_out2_2_32_port, A2 => n2946, B1 => 
                           io_out2_3_32_port, B2 => n2940, ZN => n2800);
   U3151 : AOI22_X1 port map( A1 => loc_out2_0_32_port, A2 => n2958, B1 => 
                           io_out2_0_32_port, B2 => n2952, ZN => n2801);
   U3152 : AOI22_X1 port map( A1 => loc_out2_1_32_port, A2 => n2970, B1 => 
                           loc_out2_3_32_port, B2 => n2964, ZN => n2802);
   U3153 : NAND4_X1 port map( A1 => n2796, A2 => n2797, A3 => n2798, A4 => 
                           n2799, ZN => N1165);
   U3154 : AOI22_X1 port map( A1 => io_out2_2_33_port, A2 => n2946, B1 => 
                           io_out2_3_33_port, B2 => n2940, ZN => n2796);
   U3155 : AOI22_X1 port map( A1 => loc_out2_0_33_port, A2 => n2958, B1 => 
                           io_out2_0_33_port, B2 => n2952, ZN => n2797);
   U3156 : AOI22_X1 port map( A1 => loc_out2_1_33_port, A2 => n2970, B1 => 
                           loc_out2_3_33_port, B2 => n2964, ZN => n2798);
   U3157 : NAND4_X1 port map( A1 => n2792, A2 => n2793, A3 => n2794, A4 => 
                           n2795, ZN => N1166);
   U3158 : AOI22_X1 port map( A1 => io_out2_2_34_port, A2 => n2946, B1 => 
                           io_out2_3_34_port, B2 => n2940, ZN => n2792);
   U3159 : AOI22_X1 port map( A1 => loc_out2_0_34_port, A2 => n2958, B1 => 
                           io_out2_0_34_port, B2 => n2952, ZN => n2793);
   U3160 : AOI22_X1 port map( A1 => loc_out2_1_34_port, A2 => n2970, B1 => 
                           loc_out2_3_34_port, B2 => n2964, ZN => n2794);
   U3161 : NAND4_X1 port map( A1 => n2788, A2 => n2789, A3 => n2790, A4 => 
                           n2791, ZN => N1167);
   U3162 : AOI22_X1 port map( A1 => io_out2_2_35_port, A2 => n2946, B1 => 
                           io_out2_3_35_port, B2 => n2940, ZN => n2788);
   U3163 : AOI22_X1 port map( A1 => loc_out2_0_35_port, A2 => n2958, B1 => 
                           io_out2_0_35_port, B2 => n2952, ZN => n2789);
   U3164 : AOI22_X1 port map( A1 => loc_out2_1_35_port, A2 => n2970, B1 => 
                           loc_out2_3_35_port, B2 => n2964, ZN => n2790);
   U3165 : NAND4_X1 port map( A1 => n2784, A2 => n2785, A3 => n2786, A4 => 
                           n2787, ZN => N1168);
   U3166 : AOI22_X1 port map( A1 => io_out2_2_36_port, A2 => n2947, B1 => 
                           io_out2_3_36_port, B2 => n2941, ZN => n2784);
   U3167 : AOI22_X1 port map( A1 => loc_out2_0_36_port, A2 => n2959, B1 => 
                           io_out2_0_36_port, B2 => n2953, ZN => n2785);
   U3168 : AOI22_X1 port map( A1 => loc_out2_1_36_port, A2 => n2971, B1 => 
                           loc_out2_3_36_port, B2 => n2965, ZN => n2786);
   U3169 : NAND4_X1 port map( A1 => n2780, A2 => n2781, A3 => n2782, A4 => 
                           n2783, ZN => N1169);
   U3170 : AOI22_X1 port map( A1 => io_out2_2_37_port, A2 => n2947, B1 => 
                           io_out2_3_37_port, B2 => n2941, ZN => n2780);
   U3171 : AOI22_X1 port map( A1 => loc_out2_0_37_port, A2 => n2959, B1 => 
                           io_out2_0_37_port, B2 => n2953, ZN => n2781);
   U3172 : AOI22_X1 port map( A1 => loc_out2_1_37_port, A2 => n2971, B1 => 
                           loc_out2_3_37_port, B2 => n2965, ZN => n2782);
   U3173 : NAND4_X1 port map( A1 => n2776, A2 => n2777, A3 => n2778, A4 => 
                           n2779, ZN => N1170);
   U3174 : AOI22_X1 port map( A1 => io_out2_2_38_port, A2 => n2947, B1 => 
                           io_out2_3_38_port, B2 => n2941, ZN => n2776);
   U3175 : AOI22_X1 port map( A1 => loc_out2_0_38_port, A2 => n2959, B1 => 
                           io_out2_0_38_port, B2 => n2953, ZN => n2777);
   U3176 : AOI22_X1 port map( A1 => loc_out2_1_38_port, A2 => n2971, B1 => 
                           loc_out2_3_38_port, B2 => n2965, ZN => n2778);
   U3177 : NAND4_X1 port map( A1 => n2772, A2 => n2773, A3 => n2774, A4 => 
                           n2775, ZN => N1171);
   U3178 : AOI22_X1 port map( A1 => io_out2_2_39_port, A2 => n2947, B1 => 
                           io_out2_3_39_port, B2 => n2941, ZN => n2772);
   U3179 : AOI22_X1 port map( A1 => loc_out2_0_39_port, A2 => n2959, B1 => 
                           io_out2_0_39_port, B2 => n2953, ZN => n2773);
   U3180 : AOI22_X1 port map( A1 => loc_out2_1_39_port, A2 => n2971, B1 => 
                           loc_out2_3_39_port, B2 => n2965, ZN => n2774);
   U3181 : NAND4_X1 port map( A1 => n2768, A2 => n2769, A3 => n2770, A4 => 
                           n2771, ZN => N1172);
   U3182 : AOI22_X1 port map( A1 => io_out2_2_40_port, A2 => n2947, B1 => 
                           io_out2_3_40_port, B2 => n2941, ZN => n2768);
   U3183 : AOI22_X1 port map( A1 => loc_out2_0_40_port, A2 => n2959, B1 => 
                           io_out2_0_40_port, B2 => n2953, ZN => n2769);
   U3184 : AOI22_X1 port map( A1 => loc_out2_1_40_port, A2 => n2971, B1 => 
                           loc_out2_3_40_port, B2 => n2965, ZN => n2770);
   U3185 : NAND4_X1 port map( A1 => n2764, A2 => n2765, A3 => n2766, A4 => 
                           n2767, ZN => N1173);
   U3186 : AOI22_X1 port map( A1 => io_out2_2_41_port, A2 => n2947, B1 => 
                           io_out2_3_41_port, B2 => n2941, ZN => n2764);
   U3187 : AOI22_X1 port map( A1 => loc_out2_0_41_port, A2 => n2959, B1 => 
                           io_out2_0_41_port, B2 => n2953, ZN => n2765);
   U3188 : AOI22_X1 port map( A1 => loc_out2_1_41_port, A2 => n2971, B1 => 
                           loc_out2_3_41_port, B2 => n2965, ZN => n2766);
   U3189 : NAND4_X1 port map( A1 => n2760, A2 => n2761, A3 => n2762, A4 => 
                           n2763, ZN => N1174);
   U3190 : AOI22_X1 port map( A1 => io_out2_2_42_port, A2 => n2947, B1 => 
                           io_out2_3_42_port, B2 => n2941, ZN => n2760);
   U3191 : AOI22_X1 port map( A1 => loc_out2_0_42_port, A2 => n2959, B1 => 
                           io_out2_0_42_port, B2 => n2953, ZN => n2761);
   U3192 : AOI22_X1 port map( A1 => loc_out2_1_42_port, A2 => n2971, B1 => 
                           loc_out2_3_42_port, B2 => n2965, ZN => n2762);
   U3193 : NAND4_X1 port map( A1 => n2756, A2 => n2757, A3 => n2758, A4 => 
                           n2759, ZN => N1175);
   U3194 : AOI22_X1 port map( A1 => io_out2_2_43_port, A2 => n2947, B1 => 
                           io_out2_3_43_port, B2 => n2941, ZN => n2756);
   U3195 : AOI22_X1 port map( A1 => loc_out2_0_43_port, A2 => n2959, B1 => 
                           io_out2_0_43_port, B2 => n2953, ZN => n2757);
   U3196 : AOI22_X1 port map( A1 => loc_out2_1_43_port, A2 => n2971, B1 => 
                           loc_out2_3_43_port, B2 => n2965, ZN => n2758);
   U3197 : NAND4_X1 port map( A1 => n2752, A2 => n2753, A3 => n2754, A4 => 
                           n2755, ZN => N1176);
   U3198 : AOI22_X1 port map( A1 => io_out2_2_44_port, A2 => n2947, B1 => 
                           io_out2_3_44_port, B2 => n2941, ZN => n2752);
   U3199 : AOI22_X1 port map( A1 => loc_out2_0_44_port, A2 => n2959, B1 => 
                           io_out2_0_44_port, B2 => n2953, ZN => n2753);
   U3200 : AOI22_X1 port map( A1 => loc_out2_1_44_port, A2 => n2971, B1 => 
                           loc_out2_3_44_port, B2 => n2965, ZN => n2754);
   U3201 : NAND4_X1 port map( A1 => n2748, A2 => n2749, A3 => n2750, A4 => 
                           n2751, ZN => N1177);
   U3202 : AOI22_X1 port map( A1 => io_out2_2_45_port, A2 => n2947, B1 => 
                           io_out2_3_45_port, B2 => n2941, ZN => n2748);
   U3203 : AOI22_X1 port map( A1 => loc_out2_0_45_port, A2 => n2959, B1 => 
                           io_out2_0_45_port, B2 => n2953, ZN => n2749);
   U3204 : AOI22_X1 port map( A1 => loc_out2_1_45_port, A2 => n2971, B1 => 
                           loc_out2_3_45_port, B2 => n2965, ZN => n2750);
   U3205 : NAND4_X1 port map( A1 => n2744, A2 => n2745, A3 => n2746, A4 => 
                           n2747, ZN => N1178);
   U3206 : AOI22_X1 port map( A1 => io_out2_2_46_port, A2 => n2947, B1 => 
                           io_out2_3_46_port, B2 => n2941, ZN => n2744);
   U3207 : AOI22_X1 port map( A1 => loc_out2_0_46_port, A2 => n2959, B1 => 
                           io_out2_0_46_port, B2 => n2953, ZN => n2745);
   U3208 : AOI22_X1 port map( A1 => loc_out2_1_46_port, A2 => n2971, B1 => 
                           loc_out2_3_46_port, B2 => n2965, ZN => n2746);
   U3209 : NAND4_X1 port map( A1 => n2740, A2 => n2741, A3 => n2742, A4 => 
                           n2743, ZN => N1179);
   U3210 : AOI22_X1 port map( A1 => io_out2_2_47_port, A2 => n2947, B1 => 
                           io_out2_3_47_port, B2 => n2941, ZN => n2740);
   U3211 : AOI22_X1 port map( A1 => loc_out2_0_47_port, A2 => n2959, B1 => 
                           io_out2_0_47_port, B2 => n2953, ZN => n2741);
   U3212 : AOI22_X1 port map( A1 => loc_out2_1_47_port, A2 => n2971, B1 => 
                           loc_out2_3_47_port, B2 => n2965, ZN => n2742);
   U3213 : NAND4_X1 port map( A1 => n2736, A2 => n2737, A3 => n2738, A4 => 
                           n2739, ZN => N1180);
   U3214 : AOI22_X1 port map( A1 => io_out2_2_48_port, A2 => n2948, B1 => 
                           io_out2_3_48_port, B2 => n2942, ZN => n2736);
   U3215 : AOI22_X1 port map( A1 => loc_out2_0_48_port, A2 => n2960, B1 => 
                           io_out2_0_48_port, B2 => n2954, ZN => n2737);
   U3216 : AOI22_X1 port map( A1 => loc_out2_1_48_port, A2 => n2972, B1 => 
                           loc_out2_3_48_port, B2 => n2966, ZN => n2738);
   U3217 : NAND4_X1 port map( A1 => n2732, A2 => n2733, A3 => n2734, A4 => 
                           n2735, ZN => N1181);
   U3218 : AOI22_X1 port map( A1 => io_out2_2_49_port, A2 => n2948, B1 => 
                           io_out2_3_49_port, B2 => n2942, ZN => n2732);
   U3219 : AOI22_X1 port map( A1 => loc_out2_0_49_port, A2 => n2960, B1 => 
                           io_out2_0_49_port, B2 => n2954, ZN => n2733);
   U3220 : AOI22_X1 port map( A1 => loc_out2_1_49_port, A2 => n2972, B1 => 
                           loc_out2_3_49_port, B2 => n2966, ZN => n2734);
   U3221 : NAND4_X1 port map( A1 => n2728, A2 => n2729, A3 => n2730, A4 => 
                           n2731, ZN => N1182);
   U3222 : AOI22_X1 port map( A1 => io_out2_2_50_port, A2 => n2948, B1 => 
                           io_out2_3_50_port, B2 => n2942, ZN => n2728);
   U3223 : AOI22_X1 port map( A1 => loc_out2_0_50_port, A2 => n2960, B1 => 
                           io_out2_0_50_port, B2 => n2954, ZN => n2729);
   U3224 : AOI22_X1 port map( A1 => loc_out2_1_50_port, A2 => n2972, B1 => 
                           loc_out2_3_50_port, B2 => n2966, ZN => n2730);
   U3225 : NAND4_X1 port map( A1 => n2724, A2 => n2725, A3 => n2726, A4 => 
                           n2727, ZN => N1183);
   U3226 : AOI22_X1 port map( A1 => io_out2_2_51_port, A2 => n2948, B1 => 
                           io_out2_3_51_port, B2 => n2942, ZN => n2724);
   U3227 : AOI22_X1 port map( A1 => loc_out2_0_51_port, A2 => n2960, B1 => 
                           io_out2_0_51_port, B2 => n2954, ZN => n2725);
   U3228 : AOI22_X1 port map( A1 => loc_out2_1_51_port, A2 => n2972, B1 => 
                           loc_out2_3_51_port, B2 => n2966, ZN => n2726);
   U3229 : NAND4_X1 port map( A1 => n2720, A2 => n2721, A3 => n2722, A4 => 
                           n2723, ZN => N1184);
   U3230 : AOI22_X1 port map( A1 => io_out2_2_52_port, A2 => n2948, B1 => 
                           io_out2_3_52_port, B2 => n2942, ZN => n2720);
   U3231 : AOI22_X1 port map( A1 => loc_out2_0_52_port, A2 => n2960, B1 => 
                           io_out2_0_52_port, B2 => n2954, ZN => n2721);
   U3232 : AOI22_X1 port map( A1 => loc_out2_1_52_port, A2 => n2972, B1 => 
                           loc_out2_3_52_port, B2 => n2966, ZN => n2722);
   U3233 : NAND4_X1 port map( A1 => n2716, A2 => n2717, A3 => n2718, A4 => 
                           n2719, ZN => N1185);
   U3234 : AOI22_X1 port map( A1 => io_out2_2_53_port, A2 => n2948, B1 => 
                           io_out2_3_53_port, B2 => n2942, ZN => n2716);
   U3235 : AOI22_X1 port map( A1 => loc_out2_0_53_port, A2 => n2960, B1 => 
                           io_out2_0_53_port, B2 => n2954, ZN => n2717);
   U3236 : AOI22_X1 port map( A1 => loc_out2_1_53_port, A2 => n2972, B1 => 
                           loc_out2_3_53_port, B2 => n2966, ZN => n2718);
   U3237 : NAND4_X1 port map( A1 => n2712, A2 => n2713, A3 => n2714, A4 => 
                           n2715, ZN => N1186);
   U3238 : AOI22_X1 port map( A1 => io_out2_2_54_port, A2 => n2948, B1 => 
                           io_out2_3_54_port, B2 => n2942, ZN => n2712);
   U3239 : AOI22_X1 port map( A1 => loc_out2_0_54_port, A2 => n2960, B1 => 
                           io_out2_0_54_port, B2 => n2954, ZN => n2713);
   U3240 : AOI22_X1 port map( A1 => loc_out2_1_54_port, A2 => n2972, B1 => 
                           loc_out2_3_54_port, B2 => n2966, ZN => n2714);
   U3241 : NAND4_X1 port map( A1 => n2708, A2 => n2709, A3 => n2710, A4 => 
                           n2711, ZN => N1187);
   U3242 : AOI22_X1 port map( A1 => io_out2_2_55_port, A2 => n2948, B1 => 
                           io_out2_3_55_port, B2 => n2942, ZN => n2708);
   U3243 : AOI22_X1 port map( A1 => loc_out2_0_55_port, A2 => n2960, B1 => 
                           io_out2_0_55_port, B2 => n2954, ZN => n2709);
   U3244 : AOI22_X1 port map( A1 => loc_out2_1_55_port, A2 => n2972, B1 => 
                           loc_out2_3_55_port, B2 => n2966, ZN => n2710);
   U3245 : NAND4_X1 port map( A1 => n2704, A2 => n2705, A3 => n2706, A4 => 
                           n2707, ZN => N1188);
   U3246 : AOI22_X1 port map( A1 => io_out2_2_56_port, A2 => n2948, B1 => 
                           io_out2_3_56_port, B2 => n2942, ZN => n2704);
   U3247 : AOI22_X1 port map( A1 => loc_out2_0_56_port, A2 => n2960, B1 => 
                           io_out2_0_56_port, B2 => n2954, ZN => n2705);
   U3248 : AOI22_X1 port map( A1 => loc_out2_1_56_port, A2 => n2972, B1 => 
                           loc_out2_3_56_port, B2 => n2966, ZN => n2706);
   U3249 : NAND4_X1 port map( A1 => n2700, A2 => n2701, A3 => n2702, A4 => 
                           n2703, ZN => N1189);
   U3250 : AOI22_X1 port map( A1 => io_out2_2_57_port, A2 => n2948, B1 => 
                           io_out2_3_57_port, B2 => n2942, ZN => n2700);
   U3251 : AOI22_X1 port map( A1 => loc_out2_0_57_port, A2 => n2960, B1 => 
                           io_out2_0_57_port, B2 => n2954, ZN => n2701);
   U3252 : AOI22_X1 port map( A1 => loc_out2_1_57_port, A2 => n2972, B1 => 
                           loc_out2_3_57_port, B2 => n2966, ZN => n2702);
   U3253 : NAND4_X1 port map( A1 => n2696, A2 => n2697, A3 => n2698, A4 => 
                           n2699, ZN => N1190);
   U3254 : AOI22_X1 port map( A1 => io_out2_2_58_port, A2 => n2948, B1 => 
                           io_out2_3_58_port, B2 => n2942, ZN => n2696);
   U3255 : AOI22_X1 port map( A1 => loc_out2_0_58_port, A2 => n2960, B1 => 
                           io_out2_0_58_port, B2 => n2954, ZN => n2697);
   U3256 : AOI22_X1 port map( A1 => loc_out2_1_58_port, A2 => n2972, B1 => 
                           loc_out2_3_58_port, B2 => n2966, ZN => n2698);
   U3257 : NAND4_X1 port map( A1 => n2692, A2 => n2693, A3 => n2694, A4 => 
                           n2695, ZN => N1191);
   U3258 : AOI22_X1 port map( A1 => io_out2_2_59_port, A2 => n2948, B1 => 
                           io_out2_3_59_port, B2 => n2942, ZN => n2692);
   U3259 : AOI22_X1 port map( A1 => loc_out2_0_59_port, A2 => n2960, B1 => 
                           io_out2_0_59_port, B2 => n2954, ZN => n2693);
   U3260 : AOI22_X1 port map( A1 => loc_out2_1_59_port, A2 => n2972, B1 => 
                           loc_out2_3_59_port, B2 => n2966, ZN => n2694);
   U3261 : CLKBUF_X1 port map( A => n2679, Z => n2943);
   U3262 : CLKBUF_X1 port map( A => n2678, Z => n2949);
   U3263 : CLKBUF_X1 port map( A => n2677, Z => n2955);
   U3264 : CLKBUF_X1 port map( A => n2676, Z => n2961);
   U3265 : CLKBUF_X1 port map( A => n2675, Z => n2967);
   U3266 : CLKBUF_X1 port map( A => n2674, Z => n2973);
   U3267 : CLKBUF_X1 port map( A => n2673, Z => n2979);
   U3268 : CLKBUF_X1 port map( A => n2672, Z => n2985);
   U3269 : CLKBUF_X1 port map( A => n2160, Z => n2991);
   U3270 : CLKBUF_X1 port map( A => n2159, Z => n2997);
   U3271 : CLKBUF_X1 port map( A => n2158, Z => n3003);
   U3272 : CLKBUF_X1 port map( A => n2157, Z => n3009);
   U3273 : CLKBUF_X1 port map( A => n2156, Z => n3015);
   U3274 : CLKBUF_X1 port map( A => n2155, Z => n3021);
   U3275 : CLKBUF_X1 port map( A => n2154, Z => n3027);
   U3276 : CLKBUF_X1 port map( A => n2153, Z => n3033);
   U3277 : CLKBUF_X1 port map( A => n2152, Z => n3039);
   U3278 : CLKBUF_X1 port map( A => n2147, Z => n3045);
   U3279 : CLKBUF_X1 port map( A => n2145, Z => n3051);
   U3280 : CLKBUF_X1 port map( A => n2144, Z => n3057);
   U3281 : CLKBUF_X1 port map( A => n2143, Z => n3063);

end SYN_BEHAVIORAL;
